
package interleaver_svc_pkg;

   import avm_pkg::*;
   import interleaver_tr_pkg::*;

   `include "interleaver_monitor.svh"
   `include "interleaver_nb_driver.svh"
   `include "interleaver_stimulus.svh"
   `include "interleaver_score.svh"
   `include "interleaver_cover.svh"
   `include "test_status.sv"

endpackage // interleaver_svc_pkg

