module 2b_multiply(m,a,b);
input [1:0]a,[1:0]b;
output wire [1:0]m;
assign m=a*b;
endmodule
