
module count_WIDTH8_DW01_inc_0 ( A, SUM );
  input [7:0] A;
  output [7:0] SUM;

  wire   [7:2] carry;

  HALF_ADD U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  HALF_ADD U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  HALF_ADD U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  HALF_ADD U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  HALF_ADD U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  HALF_ADD U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  INV U1 ( .I(A[0]), .ZN(SUM[0]) );
  XOR2 U2 ( .A1(carry[7]), .A2(A[7]), .Z(SUM[7]) );
endmodule


module fifo_shift_ram_DW01_inc_21 ( A, SUM );
  input [10:0] A;
  output [10:0] SUM;

  wire   [10:2] carry;

  HALF_ADD U1_1_9 ( .A(A[9]), .B(carry[9]), .CO(carry[10]), .S(SUM[9]) );
  HALF_ADD U1_1_8 ( .A(A[8]), .B(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  HALF_ADD U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  HALF_ADD U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  HALF_ADD U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  HALF_ADD U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  HALF_ADD U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  HALF_ADD U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  HALF_ADD U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  INV U1 ( .I(A[0]), .ZN(SUM[0]) );
  XOR2 U2 ( .A1(carry[10]), .A2(A[10]), .Z(SUM[10]) );
endmodule


module fifo_shift_ram_DW01_inc_20 ( A, SUM );
  input [10:0] A;
  output [10:0] SUM;

  wire   [10:2] carry;

  HALF_ADD U1_1_9 ( .A(A[9]), .B(carry[9]), .CO(carry[10]), .S(SUM[9]) );
  HALF_ADD U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  HALF_ADD U1_1_8 ( .A(A[8]), .B(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  HALF_ADD U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  HALF_ADD U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  HALF_ADD U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  HALF_ADD U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  HALF_ADD U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  HALF_ADD U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  INV U1 ( .I(A[0]), .ZN(SUM[0]) );
  XOR2 U2 ( .A1(carry[10]), .A2(A[10]), .Z(SUM[10]) );
endmodule


module fifo_shift_ram_DW01_inc_19 ( A, SUM );
  input [10:0] A;
  output [10:0] SUM;

  wire   [10:2] carry;

  HALF_ADD U1_1_9 ( .A(A[9]), .B(carry[9]), .CO(carry[10]), .S(SUM[9]) );
  HALF_ADD U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  HALF_ADD U1_1_8 ( .A(A[8]), .B(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  HALF_ADD U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  HALF_ADD U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  HALF_ADD U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  HALF_ADD U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  HALF_ADD U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  HALF_ADD U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  INV U1 ( .I(A[0]), .ZN(SUM[0]) );
  XOR2 U2 ( .A1(carry[10]), .A2(A[10]), .Z(SUM[10]) );
endmodule


module fifo_shift_ram_DW01_inc_18 ( A, SUM );
  input [10:0] A;
  output [10:0] SUM;

  wire   [10:2] carry;

  HALF_ADD U1_1_9 ( .A(A[9]), .B(carry[9]), .CO(carry[10]), .S(SUM[9]) );
  HALF_ADD U1_1_8 ( .A(A[8]), .B(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  HALF_ADD U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  HALF_ADD U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  HALF_ADD U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  HALF_ADD U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  HALF_ADD U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  HALF_ADD U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  HALF_ADD U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  INV U1 ( .I(A[0]), .ZN(SUM[0]) );
  XOR2 U2 ( .A1(carry[10]), .A2(A[10]), .Z(SUM[10]) );
endmodule


module fifo_shift_ram_DW01_inc_17 ( A, SUM );
  input [10:0] A;
  output [10:0] SUM;

  wire   [10:2] carry;

  HALF_ADD U1_1_9 ( .A(A[9]), .B(carry[9]), .CO(carry[10]), .S(SUM[9]) );
  HALF_ADD U1_1_8 ( .A(A[8]), .B(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  HALF_ADD U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  HALF_ADD U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  HALF_ADD U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  HALF_ADD U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  HALF_ADD U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  HALF_ADD U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  HALF_ADD U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  INV U1 ( .I(A[0]), .ZN(SUM[0]) );
  XOR2 U2 ( .A1(carry[10]), .A2(A[10]), .Z(SUM[10]) );
endmodule


module fifo_shift_ram_DW01_inc_16 ( A, SUM );
  input [10:0] A;
  output [10:0] SUM;

  wire   [10:2] carry;

  HALF_ADD U1_1_9 ( .A(A[9]), .B(carry[9]), .CO(carry[10]), .S(SUM[9]) );
  HALF_ADD U1_1_8 ( .A(A[8]), .B(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  HALF_ADD U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  HALF_ADD U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  HALF_ADD U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  HALF_ADD U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  HALF_ADD U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  HALF_ADD U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  HALF_ADD U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  INV U1 ( .I(A[0]), .ZN(SUM[0]) );
  XOR2 U2 ( .A1(carry[10]), .A2(A[10]), .Z(SUM[10]) );
endmodule


module fifo_shift_ram_DW01_inc_15 ( A, SUM );
  input [10:0] A;
  output [10:0] SUM;

  wire   [10:2] carry;

  HALF_ADD U1_1_9 ( .A(A[9]), .B(carry[9]), .CO(carry[10]), .S(SUM[9]) );
  HALF_ADD U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  HALF_ADD U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  HALF_ADD U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  HALF_ADD U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  HALF_ADD U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  HALF_ADD U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  HALF_ADD U1_1_8 ( .A(A[8]), .B(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  HALF_ADD U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  INV U1 ( .I(A[0]), .ZN(SUM[0]) );
  XOR2 U2 ( .A1(carry[10]), .A2(A[10]), .Z(SUM[10]) );
endmodule


module fifo_shift_ram_DW01_inc_14 ( A, SUM );
  input [10:0] A;
  output [10:0] SUM;

  wire   [10:2] carry;

  HALF_ADD U1_1_9 ( .A(A[9]), .B(carry[9]), .CO(carry[10]), .S(SUM[9]) );
  HALF_ADD U1_1_8 ( .A(A[8]), .B(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  HALF_ADD U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  HALF_ADD U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  HALF_ADD U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  HALF_ADD U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  HALF_ADD U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  HALF_ADD U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  HALF_ADD U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  INV U1 ( .I(A[0]), .ZN(SUM[0]) );
  XOR2 U2 ( .A1(carry[10]), .A2(A[10]), .Z(SUM[10]) );
endmodule


module fifo_shift_ram_DW01_inc_13 ( A, SUM );
  input [10:0] A;
  output [10:0] SUM;

  wire   [10:2] carry;

  HALF_ADD U1_1_9 ( .A(A[9]), .B(carry[9]), .CO(carry[10]), .S(SUM[9]) );
  HALF_ADD U1_1_8 ( .A(A[8]), .B(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  HALF_ADD U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  HALF_ADD U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  HALF_ADD U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  HALF_ADD U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  HALF_ADD U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  HALF_ADD U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  HALF_ADD U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  INV U1 ( .I(A[0]), .ZN(SUM[0]) );
  XOR2 U2 ( .A1(carry[10]), .A2(A[10]), .Z(SUM[10]) );
endmodule


module fifo_shift_ram_DW01_inc_12 ( A, SUM );
  input [10:0] A;
  output [10:0] SUM;

  wire   [10:2] carry;

  HALF_ADD U1_1_9 ( .A(A[9]), .B(carry[9]), .CO(carry[10]), .S(SUM[9]) );
  HALF_ADD U1_1_8 ( .A(A[8]), .B(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  HALF_ADD U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  HALF_ADD U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  HALF_ADD U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  HALF_ADD U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  HALF_ADD U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  HALF_ADD U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  HALF_ADD U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  INV U1 ( .I(A[0]), .ZN(SUM[0]) );
  XOR2 U2 ( .A1(carry[10]), .A2(A[10]), .Z(SUM[10]) );
endmodule


module fifo_shift_ram_DW01_inc_11 ( A, SUM );
  input [10:0] A;
  output [10:0] SUM;

  wire   [10:2] carry;

  HALF_ADD U1_1_9 ( .A(A[9]), .B(carry[9]), .CO(carry[10]), .S(SUM[9]) );
  HALF_ADD U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  HALF_ADD U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  HALF_ADD U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  HALF_ADD U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  HALF_ADD U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  HALF_ADD U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  HALF_ADD U1_1_8 ( .A(A[8]), .B(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  HALF_ADD U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  INV U1 ( .I(A[0]), .ZN(SUM[0]) );
  XOR2 U2 ( .A1(carry[10]), .A2(A[10]), .Z(SUM[10]) );
endmodule


module fifo_shift_ram_DW01_inc_10 ( A, SUM );
  input [10:0] A;
  output [10:0] SUM;

  wire   [10:2] carry;

  HALF_ADD U1_1_9 ( .A(A[9]), .B(carry[9]), .CO(carry[10]), .S(SUM[9]) );
  HALF_ADD U1_1_8 ( .A(A[8]), .B(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  HALF_ADD U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  HALF_ADD U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  HALF_ADD U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  HALF_ADD U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  HALF_ADD U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  HALF_ADD U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  HALF_ADD U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  INV U1 ( .I(A[0]), .ZN(SUM[0]) );
  XOR2 U2 ( .A1(carry[10]), .A2(A[10]), .Z(SUM[10]) );
endmodule


module fifo_shift_ram_DW01_inc_9 ( A, SUM );
  input [10:0] A;
  output [10:0] SUM;

  wire   [10:2] carry;

  HALF_ADD U1_1_9 ( .A(A[9]), .B(carry[9]), .CO(carry[10]), .S(SUM[9]) );
  HALF_ADD U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  HALF_ADD U1_1_8 ( .A(A[8]), .B(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  HALF_ADD U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  HALF_ADD U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  HALF_ADD U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  HALF_ADD U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  HALF_ADD U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  HALF_ADD U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  INV U1 ( .I(A[0]), .ZN(SUM[0]) );
  XOR2 U2 ( .A1(carry[10]), .A2(A[10]), .Z(SUM[10]) );
endmodule


module fifo_shift_ram_DW01_inc_8 ( A, SUM );
  input [10:0] A;
  output [10:0] SUM;

  wire   [10:2] carry;

  HALF_ADD U1_1_9 ( .A(A[9]), .B(carry[9]), .CO(carry[10]), .S(SUM[9]) );
  HALF_ADD U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  HALF_ADD U1_1_8 ( .A(A[8]), .B(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  HALF_ADD U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  HALF_ADD U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  HALF_ADD U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  HALF_ADD U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  HALF_ADD U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  HALF_ADD U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  INV U1 ( .I(A[0]), .ZN(SUM[0]) );
  XOR2 U2 ( .A1(carry[10]), .A2(A[10]), .Z(SUM[10]) );
endmodule


module fifo_shift_ram_DW01_inc_7 ( A, SUM );
  input [10:0] A;
  output [10:0] SUM;

  wire   [10:2] carry;

  HALF_ADD U1_1_9 ( .A(A[9]), .B(carry[9]), .CO(carry[10]), .S(SUM[9]) );
  HALF_ADD U1_1_8 ( .A(A[8]), .B(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  HALF_ADD U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  HALF_ADD U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  HALF_ADD U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  HALF_ADD U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  HALF_ADD U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  HALF_ADD U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  HALF_ADD U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  INV U1 ( .I(A[0]), .ZN(SUM[0]) );
  XOR2 U2 ( .A1(carry[10]), .A2(A[10]), .Z(SUM[10]) );
endmodule


module fifo_shift_ram_DW01_inc_6 ( A, SUM );
  input [10:0] A;
  output [10:0] SUM;

  wire   [10:2] carry;

  HALF_ADD U1_1_9 ( .A(A[9]), .B(carry[9]), .CO(carry[10]), .S(SUM[9]) );
  HALF_ADD U1_1_8 ( .A(A[8]), .B(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  HALF_ADD U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  HALF_ADD U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  HALF_ADD U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  HALF_ADD U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  HALF_ADD U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  HALF_ADD U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  HALF_ADD U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  INV U1 ( .I(A[0]), .ZN(SUM[0]) );
  XOR2 U2 ( .A1(carry[10]), .A2(A[10]), .Z(SUM[10]) );
endmodule


module fifo_shift_ram_DW01_inc_5 ( A, SUM );
  input [10:0] A;
  output [10:0] SUM;

  wire   [10:2] carry;

  HALF_ADD U1_1_9 ( .A(A[9]), .B(carry[9]), .CO(carry[10]), .S(SUM[9]) );
  HALF_ADD U1_1_8 ( .A(A[8]), .B(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  HALF_ADD U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  HALF_ADD U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  HALF_ADD U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  HALF_ADD U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  HALF_ADD U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  HALF_ADD U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  HALF_ADD U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  INV U1 ( .I(A[0]), .ZN(SUM[0]) );
  XOR2 U2 ( .A1(carry[10]), .A2(A[10]), .Z(SUM[10]) );
endmodule


module fifo_shift_ram_DW01_inc_4 ( A, SUM );
  input [10:0] A;
  output [10:0] SUM;

  wire   [10:2] carry;

  HALF_ADD U1_1_9 ( .A(A[9]), .B(carry[9]), .CO(carry[10]), .S(SUM[9]) );
  HALF_ADD U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  HALF_ADD U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  HALF_ADD U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  HALF_ADD U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  HALF_ADD U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  HALF_ADD U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  HALF_ADD U1_1_8 ( .A(A[8]), .B(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  HALF_ADD U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  INV U1 ( .I(A[0]), .ZN(SUM[0]) );
  XOR2 U2 ( .A1(carry[10]), .A2(A[10]), .Z(SUM[10]) );
endmodule


module fifo_shift_ram_DW01_inc_3 ( A, SUM );
  input [10:0] A;
  output [10:0] SUM;

  wire   [10:2] carry;

  HALF_ADD U1_1_9 ( .A(A[9]), .B(carry[9]), .CO(carry[10]), .S(SUM[9]) );
  HALF_ADD U1_1_8 ( .A(A[8]), .B(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  HALF_ADD U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  HALF_ADD U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  HALF_ADD U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  HALF_ADD U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  HALF_ADD U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  HALF_ADD U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  HALF_ADD U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  INV U1 ( .I(A[0]), .ZN(SUM[0]) );
  XOR2 U2 ( .A1(carry[10]), .A2(A[10]), .Z(SUM[10]) );
endmodule


module fifo_shift_ram_DW01_inc_2 ( A, SUM );
  input [10:0] A;
  output [10:0] SUM;

  wire   [10:2] carry;

  HALF_ADD U1_1_9 ( .A(A[9]), .B(carry[9]), .CO(carry[10]), .S(SUM[9]) );
  HALF_ADD U1_1_8 ( .A(A[8]), .B(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  HALF_ADD U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  HALF_ADD U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  HALF_ADD U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  HALF_ADD U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  HALF_ADD U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  HALF_ADD U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  HALF_ADD U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  INV U1 ( .I(A[0]), .ZN(SUM[0]) );
  XOR2 U2 ( .A1(carry[10]), .A2(A[10]), .Z(SUM[10]) );
endmodule


module fifo_shift_ram_DW01_inc_1 ( A, SUM );
  input [10:0] A;
  output [10:0] SUM;

  wire   [10:2] carry;

  HALF_ADD U1_1_9 ( .A(A[9]), .B(carry[9]), .CO(carry[10]), .S(SUM[9]) );
  HALF_ADD U1_1_8 ( .A(A[8]), .B(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  HALF_ADD U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  HALF_ADD U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  HALF_ADD U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  HALF_ADD U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  HALF_ADD U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  HALF_ADD U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  HALF_ADD U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  INV U1 ( .I(A[0]), .ZN(SUM[0]) );
  XOR2 U2 ( .A1(carry[10]), .A2(A[10]), .Z(SUM[10]) );
endmodule


module fifo_shift_ram_DW01_inc_0 ( A, SUM );
  input [10:0] A;
  output [10:0] SUM;

  wire   [10:2] carry;

  HALF_ADD U1_1_9 ( .A(A[9]), .B(carry[9]), .CO(carry[10]), .S(SUM[9]) );
  HALF_ADD U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  HALF_ADD U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  HALF_ADD U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  HALF_ADD U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  HALF_ADD U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  HALF_ADD U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  HALF_ADD U1_1_8 ( .A(A[8]), .B(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  HALF_ADD U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  INV U1 ( .I(A[0]), .ZN(SUM[0]) );
  XOR2 U2 ( .A1(carry[10]), .A2(A[10]), .Z(SUM[10]) );
endmodule


module mem_ctrl_DW01_inc_0 ( A, SUM );
  input [7:0] A;
  output [7:0] SUM;

  wire   [7:2] carry;

  HALF_ADD U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  HALF_ADD U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  HALF_ADD U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  HALF_ADD U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  HALF_ADD U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  HALF_ADD U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  INV U1 ( .I(A[0]), .ZN(SUM[0]) );
  XOR2 U2 ( .A1(carry[7]), .A2(A[7]), .Z(SUM[7]) );
endmodule


module rdyacpt_WIDTH8_1 ( clk, reset_n, upstream_rdy, downstream_acpt, 
        upstream_data, downstream_rdy, upstream_acpt, downstream_data );
  input [7:0] upstream_data;
  output [7:0] downstream_data;
  input clk, reset_n, upstream_rdy, downstream_acpt;
  output downstream_rdy, upstream_acpt;
  wire   v1, ready_reg, N3, N29, n1, n3, n16, n17, n18, n19, n20, n21, n22,
         n23, n24, n25, n26, n27;
  wire   [7:0] d1;

  DFF_RST v0_reg ( .D(n3), .CP(clk), .CDN(reset_n), .Q(downstream_rdy) );
  DFF_EN d1_reg_7_ ( .D(upstream_data[7]), .E(N29), .CP(clk), .Q(d1[7]) );
  DFF_EN d1_reg_5_ ( .D(upstream_data[5]), .E(N29), .CP(clk), .Q(d1[5]) );
  DFF_EN d1_reg_3_ ( .D(upstream_data[3]), .E(N29), .CP(clk), .Q(d1[3]) );
  DFF_EN d1_reg_1_ ( .D(upstream_data[1]), .E(N29), .CP(clk), .Q(d1[1]) );
  DFF_EN d1_reg_0_ ( .D(upstream_data[0]), .E(N29), .CP(clk), .Q(d1[0]) );
  DFF_EN d1_reg_2_ ( .D(upstream_data[2]), .E(N29), .CP(clk), .Q(d1[2]) );
  DFF_EN d1_reg_4_ ( .D(upstream_data[4]), .E(N29), .CP(clk), .Q(d1[4]) );
  DFF_EN d1_reg_6_ ( .D(upstream_data[6]), .E(N29), .CP(clk), .Q(d1[6]) );
  DFF d0_reg_7_ ( .D(n23), .CP(clk), .Q(downstream_data[7]) );
  DFF d0_reg_5_ ( .D(n21), .CP(clk), .Q(downstream_data[5]) );
  DFF d0_reg_3_ ( .D(n19), .CP(clk), .Q(downstream_data[3]) );
  DFF d0_reg_1_ ( .D(n17), .CP(clk), .Q(downstream_data[1]) );
  DFF d0_reg_0_ ( .D(n16), .CP(clk), .Q(downstream_data[0]) );
  DFF d0_reg_2_ ( .D(n18), .CP(clk), .Q(downstream_data[2]) );
  DFF d0_reg_4_ ( .D(n20), .CP(clk), .Q(downstream_data[4]) );
  DFF d0_reg_6_ ( .D(n22), .CP(clk), .Q(downstream_data[6]) );
  DFF_EN ready_reg_reg ( .D(N3), .E(reset_n), .CP(clk), .Q(ready_reg) );
  DFF_EN_RST v1_reg ( .D(upstream_rdy), .E(upstream_acpt), .CP(clk), .CDN(
        reset_n), .Q(v1) );
  INV U2 ( .I(reset_n), .ZN(n1) );
  NOR2 U3 ( .A1(n25), .A2(upstream_acpt), .ZN(n27) );
  NOR2 U4 ( .A1(n25), .A2(n24), .ZN(n26) );
  NOR2 U5 ( .A1(n24), .A2(n1), .ZN(N29) );
  NAND2 U6 ( .A1(N3), .A2(reset_n), .ZN(n25) );
  I_NAND3 U7 ( .A1(upstream_rdy), .B1(upstream_acpt), .B2(N3), .ZN(n3) );
  I_NOR2 U8 ( .A1(v1), .B1(ready_reg), .ZN(n24) );
  I_NAND2 U9 ( .A1(downstream_acpt), .B1(downstream_rdy), .ZN(N3) );
  AO222 U10 ( .A1(d1[6]), .A2(n27), .B1(upstream_data[6]), .B2(n26), .C1(
        downstream_data[6]), .C2(n25), .Z(n22) );
  AO222 U11 ( .A1(d1[4]), .A2(n27), .B1(upstream_data[4]), .B2(n26), .C1(
        downstream_data[4]), .C2(n25), .Z(n20) );
  AO222 U12 ( .A1(d1[2]), .A2(n27), .B1(upstream_data[2]), .B2(n26), .C1(
        downstream_data[2]), .C2(n25), .Z(n18) );
  AO222 U13 ( .A1(d1[0]), .A2(n27), .B1(upstream_data[0]), .B2(n26), .C1(
        downstream_data[0]), .C2(n25), .Z(n16) );
  AO222 U14 ( .A1(d1[1]), .A2(n27), .B1(upstream_data[1]), .B2(n26), .C1(
        downstream_data[1]), .C2(n25), .Z(n17) );
  AO222 U15 ( .A1(d1[3]), .A2(n27), .B1(upstream_data[3]), .B2(n26), .C1(
        downstream_data[3]), .C2(n25), .Z(n19) );
  AO222 U16 ( .A1(d1[5]), .A2(n27), .B1(upstream_data[5]), .B2(n26), .C1(
        downstream_data[5]), .C2(n25), .Z(n21) );
  AO222 U17 ( .A1(d1[7]), .A2(n27), .B1(upstream_data[7]), .B2(n26), .C1(
        downstream_data[7]), .C2(n25), .Z(n23) );
  INV U18 ( .I(n24), .ZN(upstream_acpt) );
endmodule


module ram2p_2kx8 ( wclk, we, re, rclk, din, waddr, raddr, dout );
  input [7:0] din;
  input [10:0] waddr;
  input [10:0] raddr;
  output [7:0] dout;
  input wclk, we, re, rclk;
  wire   N29, N30, N31, N32, N33, N34, N35, N36, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n25, n26, n28, n29, n31, n32, n34, n35, n37,
         n38, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52,
         n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66,
         n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80,
         n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94,
         n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128,
         n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139,
         n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150,
         n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
         n162, n163, n164, n165, n166, n167, n169, n170, n172, n173, n175,
         n176, n178, n179, n181, n182, n184, n185, n187, n188, n190, n191,
         n193, n194, n196, n197, n199, n200, n202, n203, n205, n206, n208,
         n209, n211, n212, n214, n215, n216, n217, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244,
         n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
         n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266,
         n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277,
         n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288,
         n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
         n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
         n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
         n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831,
         n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842,
         n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
         n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
         n865, n866, n867, n869, n870, n871, n872, n873, n874, n875, n876,
         n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
         n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
         n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
         n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
         n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
         n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
         n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964,
         n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
         n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
         n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
         n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
         n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
         n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
         n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038,
         n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048,
         n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058,
         n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068,
         n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078,
         n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
         n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
         n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108,
         n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118,
         n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1129,
         n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
         n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
         n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
         n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
         n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
         n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
         n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
         n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
         n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
         n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
         n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
         n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
         n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1259, n1260,
         n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270,
         n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280,
         n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290,
         n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300,
         n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310,
         n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320,
         n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330,
         n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340,
         n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350,
         n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360,
         n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370,
         n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380,
         n1381, n1382, n1383, n1384, n1385, n1386, n1388, n1389, n1390, n1391,
         n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401,
         n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411,
         n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421,
         n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431,
         n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441,
         n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451,
         n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461,
         n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471,
         n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481,
         n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491,
         n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501,
         n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511,
         n1512, n1513, n1514, n1515, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653,
         n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663,
         n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673,
         n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683,
         n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693,
         n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703,
         n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713,
         n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723,
         n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733,
         n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743,
         n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753,
         n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763,
         n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773,
         n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784,
         n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794,
         n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804,
         n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814,
         n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824,
         n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834,
         n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844,
         n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854,
         n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864,
         n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874,
         n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884,
         n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894,
         n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1904, n1905,
         n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915,
         n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925,
         n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935,
         n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945,
         n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955,
         n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965,
         n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975,
         n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985,
         n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995,
         n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005,
         n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015,
         n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025,
         n2026, n2027, n2028, n2029, n2030, n2031, n2033, n2034, n2035, n2036,
         n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046,
         n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056,
         n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066,
         n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076,
         n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086,
         n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096,
         n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106,
         n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116,
         n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126,
         n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136,
         n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146,
         n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156,
         n2157, n2158, n2159, n2160, n2162, n2163, n2164, n2165, n2166, n2167,
         n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177,
         n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187,
         n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197,
         n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207,
         n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217,
         n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227,
         n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237,
         n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247,
         n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257,
         n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267,
         n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277,
         n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287,
         n2288, n2289, n2290, n2292, n2293, n2294, n2295, n2296, n2297, n2298,
         n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308,
         n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318,
         n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328,
         n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338,
         n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348,
         n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358,
         n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368,
         n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378,
         n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388,
         n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398,
         n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408,
         n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418,
         n2419, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429,
         n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439,
         n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449,
         n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459,
         n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469,
         n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479,
         n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489,
         n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499,
         n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509,
         n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519,
         n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529,
         n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539,
         n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2550,
         n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560,
         n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570,
         n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580,
         n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590,
         n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600,
         n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610,
         n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620,
         n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630,
         n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640,
         n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650,
         n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660,
         n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670,
         n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2679, n2680, n2681,
         n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691,
         n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701,
         n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711,
         n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721,
         n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731,
         n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741,
         n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751,
         n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761,
         n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771,
         n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781,
         n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791,
         n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801,
         n2802, n2803, n2804, n2805, n2806, n2808, n2809, n2810, n2811, n2812,
         n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
         n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
         n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842,
         n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
         n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
         n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882,
         n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892,
         n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902,
         n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912,
         n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922,
         n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932,
         n2933, n2934, n2935, n2937, n2938, n2939, n2940, n2941, n2942, n2943,
         n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953,
         n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963,
         n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973,
         n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983,
         n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993,
         n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003,
         n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013,
         n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023,
         n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033,
         n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043,
         n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053,
         n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063,
         n3064, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074,
         n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084,
         n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094,
         n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104,
         n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114,
         n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124,
         n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134,
         n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144,
         n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154,
         n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164,
         n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174,
         n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184,
         n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3195,
         n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205,
         n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215,
         n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225,
         n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235,
         n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245,
         n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255,
         n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265,
         n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275,
         n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285,
         n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295,
         n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305,
         n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315,
         n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3325, n3326,
         n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336,
         n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346,
         n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356,
         n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366,
         n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376,
         n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386,
         n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396,
         n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406,
         n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416,
         n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426,
         n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436,
         n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446,
         n3447, n3448, n3449, n3450, n3451, n3452, n3454, n3455, n3456, n3457,
         n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467,
         n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477,
         n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487,
         n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497,
         n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507,
         n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517,
         n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527,
         n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537,
         n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547,
         n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557,
         n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567,
         n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577,
         n3578, n3579, n3580, n3581, n3583, n3584, n3585, n3586, n3587, n3588,
         n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598,
         n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608,
         n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618,
         n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628,
         n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638,
         n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648,
         n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658,
         n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668,
         n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678,
         n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688,
         n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698,
         n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708,
         n3709, n3710, n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719,
         n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729,
         n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739,
         n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749,
         n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759,
         n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769,
         n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779,
         n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789,
         n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799,
         n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809,
         n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819,
         n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829,
         n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839,
         n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850,
         n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860,
         n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870,
         n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880,
         n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890,
         n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900,
         n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910,
         n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920,
         n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930,
         n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940,
         n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950,
         n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960,
         n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3970, n3971,
         n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981,
         n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991,
         n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001,
         n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011,
         n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021,
         n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031,
         n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041,
         n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051,
         n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061,
         n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071,
         n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081,
         n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091,
         n4092, n4093, n4094, n4095, n4096, n4097, n4099, n4100, n4101, n4102,
         n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112,
         n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122,
         n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132,
         n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142,
         n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152,
         n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162,
         n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172,
         n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182,
         n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192,
         n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202,
         n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212,
         n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222,
         n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232,
         n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242,
         n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252,
         n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262,
         n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272,
         n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282,
         n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292,
         n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302,
         n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312,
         n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322,
         n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332,
         n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342,
         n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352,
         n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362,
         n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372,
         n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382,
         n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392,
         n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402,
         n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412,
         n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422,
         n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432,
         n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442,
         n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452,
         n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462,
         n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472,
         n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482,
         n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492,
         n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502,
         n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512,
         n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522,
         n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532,
         n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542,
         n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552,
         n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562,
         n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572,
         n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582,
         n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592,
         n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602,
         n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612,
         n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622,
         n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632,
         n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642,
         n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652,
         n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662,
         n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672,
         n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682,
         n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692,
         n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702,
         n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712,
         n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722,
         n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732,
         n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742,
         n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752,
         n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762,
         n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772,
         n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782,
         n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792,
         n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802,
         n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812,
         n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822,
         n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832,
         n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842,
         n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852,
         n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862,
         n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872,
         n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882,
         n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892,
         n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902,
         n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912,
         n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922,
         n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932,
         n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942,
         n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952,
         n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962,
         n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972,
         n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982,
         n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992,
         n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002,
         n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012,
         n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022,
         n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032,
         n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042,
         n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052,
         n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062,
         n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072,
         n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082,
         n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092,
         n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102,
         n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112,
         n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122,
         n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132,
         n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142,
         n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152,
         n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162,
         n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172,
         n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182,
         n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192,
         n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202,
         n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212,
         n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222,
         n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232,
         n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242,
         n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252,
         n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262,
         n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272,
         n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282,
         n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292,
         n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302,
         n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312,
         n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322,
         n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332,
         n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342,
         n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352,
         n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362,
         n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372,
         n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382,
         n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392,
         n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402,
         n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412,
         n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422,
         n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432,
         n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442,
         n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452,
         n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462,
         n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472,
         n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482,
         n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492,
         n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502,
         n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512,
         n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522,
         n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532,
         n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542,
         n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552,
         n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562,
         n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572,
         n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582,
         n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592,
         n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602,
         n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612,
         n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622,
         n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632,
         n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642,
         n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652,
         n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662,
         n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672,
         n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682,
         n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692,
         n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702,
         n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712,
         n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722,
         n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732,
         n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742,
         n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752,
         n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762,
         n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772,
         n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782,
         n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792,
         n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802,
         n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812,
         n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822,
         n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832,
         n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842,
         n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852,
         n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862,
         n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872,
         n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882,
         n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892,
         n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902,
         n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912,
         n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922,
         n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932,
         n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942,
         n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952,
         n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962,
         n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972,
         n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982,
         n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992,
         n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002,
         n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012,
         n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022,
         n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032,
         n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042,
         n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052,
         n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062,
         n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072,
         n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082,
         n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092,
         n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102,
         n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112,
         n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122,
         n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132,
         n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142,
         n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152,
         n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162,
         n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172,
         n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182,
         n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192,
         n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202,
         n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212,
         n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222,
         n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232,
         n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242,
         n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252,
         n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262,
         n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272,
         n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282,
         n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292,
         n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302,
         n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312,
         n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322,
         n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332,
         n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342,
         n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352,
         n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362,
         n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372,
         n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382,
         n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392,
         n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402,
         n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412,
         n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422,
         n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432,
         n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442,
         n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452,
         n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462,
         n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472,
         n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482,
         n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492,
         n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502,
         n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512,
         n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522,
         n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532,
         n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542,
         n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552,
         n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562,
         n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572,
         n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582,
         n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592,
         n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602,
         n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612,
         n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622,
         n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632,
         n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642,
         n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652,
         n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662,
         n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672,
         n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682,
         n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692,
         n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702,
         n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712,
         n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722,
         n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732,
         n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742,
         n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752,
         n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762,
         n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772,
         n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782,
         n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792,
         n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802,
         n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812,
         n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822,
         n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832,
         n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842,
         n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852,
         n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862,
         n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872,
         n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882,
         n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892,
         n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902,
         n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912,
         n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922,
         n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932,
         n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942,
         n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952,
         n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962,
         n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972,
         n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982,
         n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992,
         n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002,
         n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012,
         n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022,
         n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032,
         n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042,
         n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052,
         n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062,
         n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072,
         n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082,
         n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092,
         n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102,
         n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112,
         n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122,
         n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132,
         n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142,
         n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152,
         n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162,
         n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172,
         n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182,
         n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192,
         n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202,
         n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212,
         n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222,
         n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232,
         n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242,
         n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252,
         n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262,
         n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272,
         n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282,
         n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292,
         n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302,
         n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312,
         n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322,
         n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332,
         n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342,
         n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352,
         n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362,
         n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372,
         n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382,
         n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392,
         n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402,
         n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412,
         n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422,
         n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432,
         n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442,
         n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452,
         n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462,
         n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472,
         n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482,
         n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492,
         n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502,
         n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512,
         n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522,
         n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532,
         n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542,
         n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552,
         n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562,
         n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572,
         n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582,
         n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592,
         n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602,
         n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612,
         n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622,
         n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632,
         n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642,
         n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652,
         n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662,
         n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672,
         n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682,
         n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692,
         n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702,
         n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712,
         n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722,
         n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732,
         n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742,
         n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752,
         n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762,
         n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772,
         n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782,
         n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792,
         n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802,
         n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812,
         n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822,
         n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832,
         n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842,
         n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852,
         n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862,
         n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872,
         n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882,
         n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892,
         n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902,
         n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912,
         n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922,
         n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932,
         n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942,
         n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952,
         n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962,
         n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972,
         n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982,
         n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992,
         n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002,
         n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012,
         n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022,
         n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032,
         n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042,
         n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052,
         n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062,
         n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072,
         n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082,
         n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092,
         n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102,
         n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112,
         n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122,
         n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132,
         n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142,
         n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152,
         n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162,
         n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172,
         n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182,
         n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192,
         n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202,
         n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212,
         n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222,
         n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232,
         n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242,
         n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252,
         n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262,
         n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272,
         n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282,
         n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292,
         n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302,
         n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312,
         n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322,
         n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332,
         n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342,
         n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352,
         n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362,
         n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372,
         n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382,
         n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392,
         n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402,
         n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412,
         n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422,
         n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432,
         n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442,
         n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452,
         n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462,
         n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472,
         n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482,
         n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492,
         n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502,
         n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512,
         n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522,
         n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532,
         n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542,
         n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552,
         n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562,
         n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572,
         n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582,
         n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592,
         n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602,
         n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612,
         n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622,
         n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632,
         n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642,
         n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652,
         n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662,
         n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672,
         n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682,
         n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692,
         n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702,
         n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712,
         n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722,
         n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732,
         n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742,
         n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752,
         n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762,
         n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772,
         n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782,
         n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792,
         n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802,
         n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812,
         n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822,
         n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832,
         n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842,
         n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852,
         n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862,
         n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872,
         n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882,
         n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892,
         n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902,
         n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912,
         n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922,
         n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932,
         n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942,
         n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952,
         n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962,
         n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972,
         n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982,
         n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992,
         n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002,
         n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012,
         n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022,
         n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032,
         n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042,
         n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052,
         n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062,
         n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072,
         n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082,
         n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092,
         n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102,
         n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112,
         n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122,
         n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132,
         n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142,
         n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152,
         n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162,
         n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172,
         n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182,
         n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192,
         n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202,
         n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212,
         n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222,
         n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232,
         n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242,
         n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252,
         n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262,
         n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272,
         n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282,
         n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292,
         n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302,
         n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312,
         n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322,
         n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332,
         n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342,
         n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352,
         n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362,
         n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372,
         n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382,
         n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392,
         n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402,
         n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412,
         n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422,
         n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432,
         n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442,
         n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452,
         n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462,
         n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472,
         n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482,
         n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492,
         n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502,
         n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512,
         n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522,
         n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532,
         n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542,
         n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552,
         n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562,
         n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572,
         n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582,
         n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592,
         n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602,
         n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612,
         n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622,
         n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632,
         n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642,
         n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652,
         n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662,
         n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672,
         n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682,
         n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692,
         n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702,
         n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712,
         n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722,
         n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732,
         n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742,
         n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752,
         n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762,
         n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772,
         n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782,
         n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792,
         n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802,
         n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812,
         n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822,
         n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832,
         n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842,
         n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852,
         n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862,
         n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872,
         n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882,
         n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892,
         n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902,
         n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912,
         n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922,
         n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932,
         n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942,
         n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952,
         n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962,
         n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972,
         n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982,
         n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992,
         n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001,
         n10002, n10003, n10004, n10005, n10006, n10007, n10008, n10009,
         n10010, n10011, n10012, n10013, n10014, n10015, n10016, n10017,
         n10018, n10019, n10020, n10021, n10022, n10023, n10024, n10025,
         n10026, n10027, n10028, n10029, n10030, n10031, n10032, n10033,
         n10034, n10035, n10036, n10037, n10038, n10039, n10040, n10041,
         n10042, n10043, n10044, n10045, n10046, n10047, n10048, n10049,
         n10050, n10051, n10052, n10053, n10054, n10055, n10056, n10057,
         n10058, n10059, n10060, n10061, n10062, n10063, n10064, n10065,
         n10066, n10067, n10068, n10069, n10070, n10071, n10072, n10073,
         n10074, n10075, n10076, n10077, n10078, n10079, n10080, n10081,
         n10082, n10083, n10084, n10085, n10086, n10087, n10088, n10089,
         n10090, n10091, n10092, n10093, n10094, n10095, n10096, n10097,
         n10098, n10099, n10100, n10101, n10102, n10103, n10104, n10105,
         n10106, n10107, n10108, n10109, n10110, n10111, n10112, n10113,
         n10114, n10115, n10116, n10117, n10118, n10119, n10120, n10121,
         n10122, n10123, n10124, n10125, n10126, n10127, n10128, n10129,
         n10130, n10131, n10132, n10133, n10134, n10135, n10136, n10137,
         n10138, n10139, n10140, n10141, n10142, n10143, n10144, n10145,
         n10146, n10147, n10148, n10149, n10150, n10151, n10152, n10153,
         n10154, n10155, n10156, n10157, n10158, n10159, n10160, n10161,
         n10162, n10163, n10164, n10165, n10166, n10167, n10168, n10169,
         n10170, n10171, n10172, n10173, n10174, n10175, n10176, n10177,
         n10178, n10179, n10180, n10181, n10182, n10183, n10184, n10185,
         n10186, n10187, n10188, n10189, n10190, n10191, n10192, n10193,
         n10194, n10195, n10196, n10197, n10198, n10199, n10200, n10201,
         n10202, n10203, n10204, n10205, n10206, n10207, n10208, n10209,
         n10210, n10211, n10212, n10213, n10214, n10215, n10216, n10217,
         n10218, n10219, n10220, n10221, n10222, n10223, n10224, n10225,
         n10226, n10227, n10228, n10229, n10230, n10231, n10232, n10233,
         n10234, n10235, n10236, n10237, n10238, n10239, n10240, n10241,
         n10242, n10243, n10244, n10245, n10246, n10247, n10248, n10249,
         n10250, n10251, n10252, n10253, n10254, n10255, n10256, n10257,
         n10258, n10259, n10260, n10261, n10262, n10263, n10264, n10265,
         n10266, n10267, n10268, n10269, n10270, n10271, n10272, n10273,
         n10274, n10275, n10276, n10277, n10278, n10279, n10280, n10281,
         n10282, n10283, n10284, n10285, n10286, n10287, n10288, n10289,
         n10290, n10291, n10292, n10293, n10294, n10295, n10296, n10297,
         n10298, n10299, n10300, n10301, n10302, n10303, n10304, n10305,
         n10306, n10307, n10308, n10309, n10310, n10311, n10312, n10313,
         n10314, n10315, n10316, n10317, n10318, n10319, n10320, n10321,
         n10322, n10323, n10324, n10325, n10326, n10327, n10328, n10329,
         n10330, n10331, n10332, n10333, n10334, n10335, n10336, n10337,
         n10338, n10339, n10340, n10341, n10342, n10343, n10344, n10345,
         n10346, n10347, n10348, n10349, n10350, n10351, n10352, n10353,
         n10354, n10355, n10356, n10357, n10358, n10359, n10360, n10361,
         n10362, n10363, n10364, n10365, n10366, n10367, n10368, n10369,
         n10370, n10371, n10372, n10373, n10374, n10375, n10376, n10377,
         n10378, n10379, n10380, n10381, n10382, n10383, n10384, n10385,
         n10386, n10387, n10388, n10389, n10390, n10391, n10392, n10393,
         n10394, n10395, n10396, n10397, n10398, n10399, n10400, n10401,
         n10402, n10403, n10404, n10405, n10406, n10407, n10408, n10409,
         n10410, n10411, n10412, n10413, n10414, n10415, n10416, n10417,
         n10418, n10419, n10420, n10421, n10422, n10423, n10424, n10425,
         n10426, n10427, n10428, n10429, n10430, n10431, n10432, n10433,
         n10434, n10435, n10436, n10437, n10438, n10439, n10440, n10441,
         n10442, n10443, n10444, n10445, n10446, n10447, n10448, n10449,
         n10450, n10451, n10452, n10453, n10454, n10455, n10456, n10457,
         n10458, n10459, n10460, n10461, n10462, n10463, n10464, n10465,
         n10466, n10467, n10468, n10469, n10470, n10471, n10472, n10473,
         n10474, n10475, n10476, n10477, n10478, n10479, n10480, n10481,
         n10482, n10483, n10484, n10485, n10486, n10487, n10488, n10489,
         n10490, n10491, n10492, n10493, n10494, n10495, n10496, n10497,
         n10498, n10499, n10500, n10501, n10502, n10503, n10504, n10505,
         n10506, n10507, n10508, n10509, n10510, n10511, n10512, n10513,
         n10514, n10515, n10516, n10517, n10518, n10519, n10520, n10521,
         n10522, n10523, n10524, n10525, n10526, n10527, n10528, n10529,
         n10530, n10531, n10532, n10533, n10534, n10535, n10536, n10537,
         n10538, n10539, n10540, n10541, n10542, n10543, n10544, n10545,
         n10546, n10547, n10548, n10549, n10550, n10551, n10552, n10553,
         n10554, n10555, n10556, n10557, n10558, n10559, n10560, n10561,
         n10562, n10563, n10564, n10565, n10566, n10567, n10568, n10569,
         n10570, n10571, n10572, n10573, n10574, n10575, n10576, n10577,
         n10578, n10579, n10580, n10581, n10582, n10583, n10584, n10585,
         n10586, n10587, n10588, n10589, n10590, n10591, n10592, n10593,
         n10594, n10595, n10596, n10597, n10598, n10599, n10600, n10601,
         n10602, n10603, n10604, n10605, n10606, n10607, n10608, n10609,
         n10610, n10611, n10612, n10613, n10614, n10615, n10616, n10617,
         n10618, n10619, n10620, n10621, n10622, n10623, n10624, n10625,
         n10626, n10627, n10628, n10629, n10630, n10631, n10632, n10633,
         n10634, n10635, n10636, n10637, n10638, n10639, n10640, n10641,
         n10642, n10643, n10644, n10645, n10646, n10647, n10648, n10649,
         n10650, n10651, n10652, n10653, n10654, n10655, n10656, n10657,
         n10658, n10659, n10660, n10661, n10662, n10663, n10664, n10665,
         n10666, n10667, n10668, n10669, n10670, n10671, n10672, n10673,
         n10674, n10675, n10676, n10677, n10678, n10679, n10680, n10681,
         n10682, n10683, n10684, n10685, n10686, n10687, n10688, n10689,
         n10690, n10691, n10692, n10693, n10694, n10695, n10696, n10697,
         n10698, n10699, n10700, n10701, n10702, n10703, n10704, n10705,
         n10706, n10707, n10708, n10709, n10710, n10711, n10712, n10713,
         n10714, n10715, n10716, n10717, n10718, n10719, n10720, n10721,
         n10722, n10723, n10724, n10725, n10726, n10727, n10728, n10729,
         n10730, n10731, n10732, n10733, n10734, n10735, n10736, n10737,
         n10738, n10739, n10740, n10741, n10742, n10743, n10744, n10745,
         n10746, n10747, n10748, n10749, n10750, n10751, n10752, n10753,
         n10754, n10755, n10756, n10757, n10758, n10759, n10760, n10761,
         n10762, n10763, n10764, n10765, n10766, n10767, n10768, n10769,
         n10770, n10771, n10772, n10773, n10774, n10775, n10776, n10777,
         n10778, n10779, n10780, n10781, n10782, n10783, n10784, n10785,
         n10786, n10787, n10788, n10789, n10790, n10791, n10792, n10793,
         n10794, n10795, n10796, n10797, n10798, n10799, n10800, n10801,
         n10802, n10803, n10804, n10805, n10806, n10807, n10808, n10809,
         n10810, n10811, n10812, n10813, n10814, n10815, n10816, n10817,
         n10818, n10819, n10820, n10821, n10822, n10823, n10824, n10825,
         n10826, n10827, n10828, n10829, n10830, n10831, n10832, n10833,
         n10834, n10835, n10836, n10837, n10838, n10839, n10840, n10841,
         n10842, n10843, n10844, n10845, n10846, n10847, n10848, n10849,
         n10850, n10851, n10852, n10853, n10854, n10855, n10856, n10857,
         n10858, n10859, n10860, n10861, n10862, n10863, n10864, n10865,
         n10866, n10867, n10868, n10869, n10870, n10871, n10872, n10873,
         n10874, n10875, n10876, n10877, n10878, n10879, n10880, n10881,
         n10882, n10883, n10884, n10885, n10886, n10887, n10888, n10889,
         n10890, n10891, n10892, n10893, n10894, n10895, n10896, n10897,
         n10898, n10899, n10900, n10901, n10902, n10903, n10904, n10905,
         n10906, n10907, n10908, n10909, n10910, n10911, n10912, n10913,
         n10914, n10915, n10916, n10917, n10918, n10919, n10920, n10921,
         n10922, n10923, n10924, n10925, n10926, n10927, n10928, n10929,
         n10930, n10931, n10932, n10933, n10934, n10935, n10936, n10937,
         n10938, n10939, n10940, n10941, n10942, n10943, n10944, n10945,
         n10946, n10947, n10948, n10949, n10950, n10951, n10952, n10953,
         n10954, n10955, n10956, n10957, n10958, n10959, n10960, n10961,
         n10962, n10963, n10964, n10965, n10966, n10967, n10968, n10969,
         n10970, n10971, n10972, n10973, n10974, n10975, n10976, n10977,
         n10978, n10979, n10980, n10981, n10982, n10983, n10984, n10985,
         n10986, n10987, n10988, n10989, n10990, n10991, n10992, n10993,
         n10994, n10995, n10996, n10997, n10998, n10999, n11000, n11001,
         n11002, n11003, n11004, n11005, n11006, n11007, n11008, n11009,
         n11010, n11011, n11012, n11013, n11014, n11015, n11016, n11017,
         n11018, n11019, n11020, n11021, n11022, n11023, n11024, n11025,
         n11026, n11027, n11028, n11029, n11030, n11031, n11032, n11033,
         n11034, n11035, n11036, n11037, n11038, n11039, n11040, n11041,
         n11042, n11043, n11044, n11045, n11046, n11047, n11048, n11049,
         n11050, n11051, n11052, n11053, n11054, n11055, n11056, n11057,
         n11058, n11059, n11060, n11061, n11062, n11063, n11064, n11065,
         n11066, n11067, n11068, n11069, n11070, n11071, n11072, n11073,
         n11074, n11075, n11076, n11077, n11078, n11079, n11080, n11081,
         n11082, n11083, n11084, n11085, n11086, n11087, n11088, n11089,
         n11090, n11091, n11092, n11093, n11094, n11095, n11096, n11097,
         n11098, n11099, n11100, n11101, n11102, n11103, n11104, n11105,
         n11106, n11107, n11108, n11109, n11110, n11111, n11112, n11113,
         n11114, n11115, n11116, n11117, n11118, n11119, n11120, n11121,
         n11122, n11123, n11124, n11125, n11126, n11127, n11128, n11129,
         n11130, n11131, n11132, n11133, n11134, n11135, n11136, n11137,
         n11138, n11139, n11140, n11141, n11142, n11143, n11144, n11145,
         n11146, n11147, n11148, n11149, n11150, n11151, n11152, n11153,
         n11154, n11155, n11156, n11157, n11158, n11159, n11160, n11161,
         n11162, n11163, n11164, n11165, n11166, n11167, n11168, n11169,
         n11170, n11171, n11172, n11173, n11174, n11175, n11176, n11177,
         n11178, n11179, n11180, n11181, n11182, n11183, n11184, n11185,
         n11186, n11187, n11188, n11189, n11190, n11191, n11192, n11193,
         n11194, n11195, n11196, n11197, n11198, n11199, n11200, n11201,
         n11202, n11203, n11204, n11205, n11206, n11207, n11208, n11209,
         n11210, n11211, n11212, n11213, n11214, n11215, n11216, n11217,
         n11218, n11219, n11220, n11221, n11222, n11223, n11224, n11225,
         n11226, n11227, n11228, n11229, n11230, n11231, n11232, n11233,
         n11234, n11235, n11236, n11237, n11238, n11239, n11240, n11241,
         n11242, n11243, n11244, n11245, n11246, n11247, n11248, n11249,
         n11250, n11251, n11252, n11253, n11254, n11255, n11256, n11257,
         n11258, n11259, n11260, n11261, n11262, n11263, n11264, n11265,
         n11266, n11267, n11268, n11269, n11270, n11271, n11272, n11273,
         n11274, n11275, n11276, n11277, n11278, n11279, n11280, n11281,
         n11282, n11283, n11284, n11285, n11286, n11287, n11288, n11289,
         n11290, n11291, n11292, n11293, n11294, n11295, n11296, n11297,
         n11298, n11299, n11300, n11301, n11302, n11303, n11304, n11305,
         n11306, n11307, n11308, n11309, n11310, n11311, n11312, n11313,
         n11314, n11315, n11316, n11317, n11318, n11319, n11320, n11321,
         n11322, n11323, n11324, n11325, n11326, n11327, n11328, n11329,
         n11330, n11331, n11332, n11333, n11334, n11335, n11336, n11337,
         n11338, n11339, n11340, n11341, n11342, n11343, n11344, n11345,
         n11346, n11347, n11348, n11349, n11350, n11351, n11352, n11353,
         n11354, n11355, n11356, n11357, n11358, n11359, n11360, n11361,
         n11362, n11363, n11364, n11365, n11366, n11367, n11368, n11369,
         n11370, n11371, n11372, n11373, n11374, n11375, n11376, n11377,
         n11378, n11379, n11380, n11381, n11382, n11383, n11384, n11385,
         n11386, n11387, n11388, n11389, n11390, n11391, n11392, n11393,
         n11394, n11395, n11396, n11397, n11398, n11399, n11400, n11401,
         n11402, n11403, n11404, n11405, n11406, n11407, n11408, n11409,
         n11410, n11411, n11412, n11413, n11414, n11415, n11416, n11417,
         n11418, n11419, n11420, n11421, n11422, n11423, n11424, n11425,
         n11426, n11427, n11428, n11429, n11430, n11431, n11432, n11433,
         n11434, n11435, n11436, n11437, n11438, n11439, n11440, n11441,
         n11442, n11443, n11444, n11445, n11446, n11447, n11448, n11449,
         n11450, n11451, n11452, n11453, n11454, n11455, n11456, n11457,
         n11458, n11459, n11460, n11461, n11462, n11463, n11464, n11465,
         n11466, n11467, n11468, n11469, n11470, n11471, n11472, n11473,
         n11474, n11475, n11476, n11477, n11478, n11479, n11480, n11481,
         n11482, n11483, n11484, n11485, n11486, n11487, n11488, n11489,
         n11490, n11491, n11492, n11493, n11494, n11495, n11496, n11497,
         n11498, n11499, n11500, n11501, n11502, n11503, n11504, n11505,
         n11506, n11507, n11508, n11509, n11510, n11511, n11512, n11513,
         n11514, n11515, n11516, n11517, n11518, n11519, n11520, n11521,
         n11522, n11523, n11524, n11525, n11526, n11527, n11528, n11529,
         n11530, n11531, n11532, n11533, n11534, n11535, n11536, n11537,
         n11538, n11539, n11540, n11541, n11542, n11543, n11544, n11545,
         n11546, n11547, n11548, n11549, n11550, n11551, n11552, n11553,
         n11554, n11555, n11556, n11557, n11558, n11559, n11560, n11561,
         n11562, n11563, n11564, n11565, n11566, n11567, n11568, n11569,
         n11570, n11571, n11572, n11573, n11574, n11575, n11576, n11577,
         n11578, n11579, n11580, n11581, n11582, n11583, n11584, n11585,
         n11586, n11587, n11588, n11589, n11590, n11591, n11592, n11593,
         n11594, n11595, n11596, n11597, n11598, n11599, n11600, n11601,
         n11602, n11603, n11604, n11605, n11606, n11607, n11608, n11609,
         n11610, n11611, n11612, n11613, n11614, n11615, n11616, n11617,
         n11618, n11619, n11620, n11621, n11622, n11623, n11624, n11625,
         n11626, n11627, n11628, n11629, n11630, n11631, n11632, n11633,
         n11634, n11635, n11636, n11637, n11638, n11639, n11640, n11641,
         n11642, n11643, n11644, n11645, n11646, n11647, n11648, n11649,
         n11650, n11651, n11652, n11653, n11654, n11655, n11656, n11657,
         n11658, n11659, n11660, n11661, n11662, n11663, n11664, n11665,
         n11666, n11667, n11668, n11669, n11670, n11671, n11672, n11673,
         n11674, n11675, n11676, n11677, n11678, n11679, n11680, n11681,
         n11682, n11683, n11684, n11685, n11686, n11687, n11688, n11689,
         n11690, n11691, n11692, n11693, n11694, n11695, n11696, n11697,
         n11698, n11699, n11700, n11701, n11702, n11703, n11704, n11705,
         n11706, n11707, n11708, n11709, n11710, n11711, n11712, n11713,
         n11714, n11715, n11716, n11717, n11718, n11719, n11720, n11721,
         n11722, n11723, n11724, n11725, n11726, n11727, n11728, n11729,
         n11730, n11731, n11732, n11733, n11734, n11735, n11736, n11737,
         n11738, n11739, n11740, n11741, n11742, n11743, n11744, n11745,
         n11746, n11747, n11748, n11749, n11750, n11751, n11752, n11753,
         n11754, n11755, n11756, n11757, n11758, n11759, n11760, n11761,
         n11762, n11763, n11764, n11765, n11766, n11767, n11768, n11769,
         n11770, n11771, n11772, n11773, n11774, n11775, n11776, n11777,
         n11778, n11779, n11780, n11781, n11782, n11783, n11784, n11785,
         n11786, n11787, n11788, n11789, n11790, n11791, n11792, n11793,
         n11794, n11795, n11796, n11797, n11798, n11799, n11800, n11801,
         n11802, n11803, n11804, n11805, n11806, n11807, n11808, n11809,
         n11810, n11811, n11812, n11813, n11814, n11815, n11816, n11817,
         n11818, n11819, n11820, n11821, n11822, n11823, n11824, n11825,
         n11826, n11827, n11828, n11829, n11830, n11831, n11832, n11833,
         n11834, n11835, n11836, n11837, n11838, n11839, n11840, n11841,
         n11842, n11843, n11844, n11845, n11846, n11847, n11848, n11849,
         n11850, n11851, n11852, n11853, n11854, n11855, n11856, n11857,
         n11858, n11859, n11860, n11861, n11862, n11863, n11864, n11865,
         n11866, n11867, n11868, n11869, n11870, n11871, n11872, n11873,
         n11874, n11875, n11876, n11877, n11878, n11879, n11880, n11881,
         n11882, n11883, n11884, n11885, n11886, n11887, n11888, n11889,
         n11890, n11891, n11892, n11893, n11894, n11895, n11896, n11897,
         n11898, n11899, n11900, n11901, n11902, n11903, n11904, n11905,
         n11906, n11907, n11908, n11909, n11910, n11911, n11912, n11913,
         n11914, n11915, n11916, n11917, n11918, n11919, n11920, n11921,
         n11922, n11923, n11924, n11925, n11926, n11927, n11928, n11929,
         n11930, n11931, n11932, n11933, n11934, n11935, n11936, n11937,
         n11938, n11939, n11940, n11941, n11942, n11943, n11944, n11945,
         n11946, n11947, n11948, n11949, n11950, n11951, n11952, n11953,
         n11954, n11955, n11956, n11957, n11958, n11959, n11960, n11961,
         n11962, n11963, n11964, n11965, n11966, n11967, n11968, n11969,
         n11970, n11971, n11972, n11973, n11974, n11975, n11976, n11977,
         n11978, n11979, n11980, n11981, n11982, n11983, n11984, n11985,
         n11986, n11987, n11988, n11989, n11990, n11991, n11992, n11993,
         n11994, n11995, n11996, n11997, n11998, n11999, n12000, n12001,
         n12002, n12003, n12004, n12005, n12006, n12007, n12008, n12009,
         n12010, n12011, n12012, n12013, n12014, n12015, n12016, n12017,
         n12018, n12019, n12020, n12021, n12022, n12023, n12024, n12025,
         n12026, n12027, n12028, n12029, n12030, n12031, n12032, n12033,
         n12034, n12035, n12036, n12037, n12038, n12039, n12040, n12041,
         n12042, n12043, n12044, n12045, n12046, n12047, n12048, n12049,
         n12050, n12051, n12052, n12053, n12054, n12055, n12056, n12057,
         n12058, n12059, n12060, n12061, n12062, n12063, n12064, n12065,
         n12066, n12067, n12068, n12069, n12070, n12071, n12072, n12073,
         n12074, n12075, n12076, n12077, n12078, n12079, n12080, n12081,
         n12082, n12083, n12084, n12085, n12086, n12087, n12088, n12089,
         n12090, n12091, n12092, n12093, n12094, n12095, n12096, n12097,
         n12098, n12099, n12100, n12101, n12102, n12103, n12104, n12105,
         n12106, n12107, n12108, n12109, n12110, n12111, n12112, n12113,
         n12114, n12115, n12116, n12117, n12118, n12119, n12120, n12121,
         n12122, n12123, n12124, n12125, n12126, n12127, n12128, n12129,
         n12130, n12131, n12132, n12133, n12134, n12135, n12136, n12137,
         n12138, n12139, n12140, n12141, n12142, n12143, n12144, n12145,
         n12146, n12147, n12148, n12149, n12150, n12151, n12152, n12153,
         n12154, n12155, n12156, n12157, n12158, n12159, n12160, n12161,
         n12162, n12163, n12164, n12165, n12166, n12167, n12168, n12169,
         n12170, n12171, n12172, n12173, n12174, n12175, n12176, n12177,
         n12178, n12179, n12180, n12181, n12182, n12183, n12184, n12185,
         n12186, n12187, n12188, n12189, n12190, n12191, n12192, n12193,
         n12194, n12195, n12196, n12197, n12198, n12199, n12200, n12201,
         n12202, n12203, n12204, n12205, n12206, n12207, n12208, n12209,
         n12210, n12211, n12212, n12213, n12214, n12215, n12216, n12217,
         n12218, n12219, n12220, n12221, n12222, n12223, n12224, n12225,
         n12226, n12227, n12228, n12229, n12230, n12231, n12232, n12233,
         n12234, n12235, n12236, n12237, n12238, n12239, n12240, n12241,
         n12242, n12243, n12244, n12245, n12246, n12247, n12248, n12249,
         n12250, n12251, n12252, n12253, n12254, n12255, n12256, n12257,
         n12258, n12259, n12260, n12261, n12262, n12263, n12264, n12265,
         n12266, n12267, n12268, n12269, n12270, n12271, n12272, n12273,
         n12274, n12275, n12276, n12277, n12278, n12279, n12280, n12281,
         n12282, n12283, n12284, n12285, n12286, n12287, n12288, n12289,
         n12290, n12291, n12292, n12293, n12294, n12295, n12296, n12297,
         n12298, n12299, n12300, n12301, n12302, n12303, n12304, n12305,
         n12306, n12307, n12308, n12309, n12310, n12311, n12312, n12313,
         n12314, n12315, n12316, n12317, n12318, n12319, n12320, n12321,
         n12322, n12323, n12324, n12325, n12326, n12327, n12328, n12329,
         n12330, n12331, n12332, n12333, n12334, n12335, n12336, n12337,
         n12338, n12339, n12340, n12341, n12342, n12343, n12344, n12345,
         n12346, n12347, n12348, n12349, n12350, n12351, n12352, n12353,
         n12354, n12355, n12356, n12357, n12358, n12359, n12360, n12361,
         n12362, n12363, n12364, n12365, n12366, n12367, n12368, n12369,
         n12370, n12371, n12372, n12373, n12374, n12375, n12376, n12377,
         n12378, n12379, n12380, n12381, n12382, n12383, n12384, n12385,
         n12386, n12387, n12388, n12389, n12390, n12391, n12392, n12393,
         n12394, n12395, n12396, n12397, n12398, n12399, n12400, n12401,
         n12402, n12403, n12404, n12405, n12406, n12407, n12408, n12409,
         n12410, n12411, n12412, n12413, n12414, n12415, n12416, n12417,
         n12418, n12419, n12420, n12421, n12422, n12423, n12424, n12425,
         n12426, n12427, n12428, n12429, n12430, n12431, n12432, n12433,
         n12434, n12435, n12436, n12437, n12438, n12439, n12440, n12441,
         n12442, n12443, n12444, n12445, n12446, n12447, n12448, n12449,
         n12450, n12451, n12452, n12453, n12454, n12455, n12456, n12457,
         n12458, n12459, n12460, n12461, n12462, n12463, n12464, n12465,
         n12466, n12467, n12468, n12469, n12470, n12471, n12472, n12473,
         n12474, n12475, n12476, n12477, n12478, n12479, n12480, n12481,
         n12482, n12483, n12484, n12485, n12486, n12487, n12488, n12489,
         n12490, n12491, n12492, n12493, n12494, n12495, n12496, n12497,
         n12498, n12499, n12500, n12501, n12502, n12503, n12504, n12505,
         n12506, n12507, n12508, n12509, n12510, n12511, n12512, n12513,
         n12514, n12515, n12516, n12517, n12518, n12519, n12520, n12521,
         n12522, n12523, n12524, n12525, n12526, n12527, n12528, n12529,
         n12530, n12531, n12532, n12533, n12534, n12535, n12536, n12537,
         n12538, n12539, n12540, n12541, n12542, n12543, n12544, n12545,
         n12546, n12547, n12548, n12549, n12550, n12551, n12552, n12553,
         n12554, n12555, n12556, n12557, n12558, n12559, n12560, n12561,
         n12562, n12563, n12564, n12565, n12566, n12567, n12568, n12569,
         n12570, n12571, n12572, n12573, n12574, n12575, n12576, n12577,
         n12578, n12579, n12580, n12581, n12582, n12583, n12584, n12585,
         n12586, n12587, n12588, n12589, n12590, n12591, n12592, n12593,
         n12594, n12595, n12596, n12597, n12598, n12599, n12600, n12601,
         n12602, n12603, n12604, n12605, n12606, n12607, n12608, n12609,
         n12610, n12611, n12612, n12613, n12614, n12615, n12616, n12617,
         n12618, n12619, n12620, n12621, n12622, n12623, n12624, n12625,
         n12626, n12627, n12628, n12629, n12630, n12631, n12632, n12633,
         n12634, n12635, n12636, n12637, n12638, n12639, n12640, n12641,
         n12642, n12643, n12644, n12645, n12646, n12647, n12648, n12649,
         n12650, n12651, n12652, n12653, n12654, n12655, n12656, n12657,
         n12658, n12659, n12660, n12661, n12662, n12663, n12664, n12665,
         n12666, n12667, n12668, n12669, n12670, n12671, n12672, n12673,
         n12674, n12675, n12676, n12677, n12678, n12679, n12680, n12681,
         n12682, n12683, n12684, n12685, n12686, n12687, n12688, n12689,
         n12690, n12691, n12692, n12693, n12694, n12695, n12696, n12697,
         n12698, n12699, n12700, n12701, n12702, n12703, n12704, n12705,
         n12706, n12707, n12708, n12709, n12710, n12711, n12712, n12713,
         n12714, n12715, n12716, n12717, n12718, n12719, n12720, n12721,
         n12722, n12723, n12724, n12725, n12726, n12727, n12728, n12729,
         n12730, n12731, n12732, n12733, n12734, n12735, n12736, n12737,
         n12738, n12739, n12740, n12741, n12742, n12743, n12744, n12745,
         n12746, n12747, n12748, n12749, n12750, n12751, n12752, n12753,
         n12754, n12755, n12756, n12757, n12758, n12759, n12760, n12761,
         n12762, n12763, n12764, n12765, n12766, n12767, n12768, n12769,
         n12770, n12771, n12772, n12773, n12774, n12775, n12776, n12777,
         n12778, n12779, n12780, n12781, n12782, n12783, n12784, n12785,
         n12786, n12787, n12788, n12789, n12790, n12791, n12792, n12793,
         n12794, n12795, n12796, n12797, n12798, n12799, n12800, n12801,
         n12802, n12803, n12804, n12805, n12806, n12807, n12808, n12809,
         n12810, n12811, n12812, n12813, n12814, n12815, n12816, n12817,
         n12818, n12819, n12820, n12821, n12822, n12823, n12824, n12825,
         n12826, n12827, n12828, n12829, n12830, n12831, n12832, n12833,
         n12834, n12835, n12836, n12837, n12838, n12839, n12840, n12841,
         n12842, n12843, n12844, n12845, n12846, n12847, n12848, n12849,
         n12850, n12851, n12852, n12853, n12854, n12855, n12856, n12857,
         n12858, n12859, n12860, n12861, n12862, n12863, n12864, n12865,
         n12866, n12867, n12868, n12869, n12870, n12871, n12872, n12873,
         n12874, n12875, n12876, n12877, n12878, n12879, n12880, n12881,
         n12882, n12883, n12884, n12885, n12886, n12887, n12888, n12889,
         n12890, n12891, n12892, n12893, n12894, n12895, n12896, n12897,
         n12898, n12899, n12900, n12901, n12902, n12903, n12904, n12905,
         n12906, n12907, n12908, n12909, n12910, n12911, n12912, n12913,
         n12914, n12915, n12916, n12917, n12918, n12919, n12920, n12921,
         n12922, n12923, n12924, n12925, n12926, n12927, n12928, n12929,
         n12930, n12931, n12932, n12933, n12934, n12935, n12936, n12937,
         n12938, n12939, n12940, n12941, n12942, n12943, n12944, n12945,
         n12946, n12947, n12948, n12949, n12950, n12951, n12952, n12953,
         n12954, n12955, n12956, n12957, n12958, n12959, n12960, n12961,
         n12962, n12963, n12964, n12965, n12966, n12967, n12968, n12969,
         n12970, n12971, n12972, n12973, n12974, n12975, n12976, n12977,
         n12978, n12979, n12980, n12981, n12982, n12983, n12984, n12985,
         n12986, n12987, n12988, n12989, n12990, n12991, n12992, n12993,
         n12994, n12995, n12996, n12997, n12998, n12999, n13000, n13001,
         n13002, n13003, n13004, n13005, n13006, n13007, n13008, n13009,
         n13010, n13011, n13012, n13013, n13014, n13015, n13016, n13017,
         n13018, n13019, n13020, n13021, n13022, n13023, n13024, n13025,
         n13026, n13027, n13028, n13029, n13030, n13031, n13032, n13033,
         n13034, n13035, n13036, n13037, n13038, n13039, n13040, n13041,
         n13042, n13043, n13044, n13045, n13046, n13047, n13048, n13049,
         n13050, n13051, n13052, n13053, n13054, n13055, n13056, n13057,
         n13058, n13059, n13060, n13061, n13062, n13063, n13064, n13065,
         n13066, n13067, n13068, n13069, n13070, n13071, n13072, n13073,
         n13074, n13075, n13076, n13077, n13078, n13079, n13080, n13081,
         n13082, n13083, n13084, n13085, n13086, n13087, n13088, n13089,
         n13090, n13091, n13092, n13093, n13094, n13095, n13096, n13097,
         n13098, n13099, n13100, n13101, n13102, n13103, n13104, n13105,
         n13106, n13107, n13108, n13109, n13110, n13111, n13112, n13113,
         n13114, n13115, n13116, n13117, n13118, n13119, n13120, n13121,
         n13122, n13123, n13124, n13125, n13126, n13127, n13128, n13129,
         n13130, n13131, n13132, n13133, n13134, n13135, n13136, n13137,
         n13138, n13139, n13140, n13141, n13142, n13143, n13144, n13145,
         n13146, n13147, n13148, n13149, n13150, n13151, n13152, n13153,
         n13154, n13155, n13156, n13157, n13158, n13159, n13160, n13161,
         n13162, n13163, n13164, n13165, n13166, n13167, n13168, n13169,
         n13170, n13171, n13172, n13173, n13174, n13175, n13176, n13177,
         n13178, n13179, n13180, n13181, n13182, n13183, n13184, n13185,
         n13186, n13187, n13188, n13189, n13190, n13191, n13192, n13193,
         n13194, n13195, n13196, n13197, n13198, n13199, n13200, n13201,
         n13202, n13203, n13204, n13205, n13206, n13207, n13208, n13209,
         n13210, n13211, n13212, n13213, n13214, n13215, n13216, n13217,
         n13218, n13219, n13220, n13221, n13222, n13223, n13224, n13225,
         n13226, n13227, n13228, n13229, n13230, n13231, n13232, n13233,
         n13234, n13235, n13236, n13237, n13238, n13239, n13240, n13241,
         n13242, n13243, n13244, n13245, n13246, n13247, n13248, n13249,
         n13250, n13251, n13252, n13253, n13254, n13255, n13256, n13257,
         n13258, n13259, n13260, n13261, n13262, n13263, n13264, n13265,
         n13266, n13267, n13268, n13269, n13270, n13271, n13272, n13273,
         n13274, n13275, n13276, n13277, n13278, n13279, n13280, n13281,
         n13282, n13283, n13284, n13285, n13286, n13287, n13288, n13289,
         n13290, n13291, n13292, n13293, n13294, n13295, n13296, n13297,
         n13298, n13299, n13300, n13301, n13302, n13303, n13304, n13305,
         n13306, n13307, n13308, n13309, n13310, n13311, n13312, n13313,
         n13314, n13315, n13316, n13317, n13318, n13319, n13320, n13321,
         n13322, n13323, n13324, n13325, n13326, n13327, n13328, n13329,
         n13330, n13331, n13332, n13333, n13334, n13335, n13336, n13337,
         n13338, n13339, n13340, n13341, n13342, n13343, n13344, n13345,
         n13346, n13347, n13348, n13349, n13350, n13351, n13352, n13353,
         n13354, n13355, n13356, n13357, n13358, n13359, n13360, n13361,
         n13362, n13363, n13364, n13365, n13366, n13367, n13368, n13369,
         n13370, n13371, n13372, n13373, n13374, n13375, n13376, n13377,
         n13378, n13379, n13380, n13381, n13382, n13383, n13384, n13385,
         n13386, n13387, n13388, n13389, n13390, n13391, n13392, n13393,
         n13394, n13395, n13396, n13397, n13398, n13399, n13400, n13401,
         n13402, n13403, n13404, n13405, n13406, n13407, n13408, n13409,
         n13410, n13411, n13412, n13413, n13414, n13415, n13416, n13417,
         n13418, n13419, n13420, n13421, n13422, n13423, n13424, n13425,
         n13426, n13427, n13428, n13429, n13430, n13431, n13432, n13433,
         n13434, n13435, n13436, n13437, n13438, n13439, n13440, n13441,
         n13442, n13443, n13444, n13445, n13446, n13447, n13448, n13449,
         n13450, n13451, n13452, n13453, n13454, n13455, n13456, n13457,
         n13458, n13459, n13460, n13461, n13462, n13463, n13464, n13465,
         n13466, n13467, n13468, n13469, n13470, n13471, n13472, n13473,
         n13474, n13475, n13476, n13477, n13478, n13479, n13480, n13481,
         n13482, n13483, n13484, n13485, n13486, n13487, n13488, n13489,
         n13490, n13491, n13492, n13493, n13494, n13495, n13496, n13497,
         n13498, n13499, n13500, n13501, n13502, n13503, n13504, n13505,
         n13506, n13507, n13508, n13509, n13510, n13511, n13512, n13513,
         n13514, n13515, n13516, n13517, n13518, n13519, n13520, n13521,
         n13522, n13523, n13524, n13525, n13526, n13527, n13528, n13529,
         n13530, n13531, n13532, n13533, n13534, n13535, n13536, n13537,
         n13538, n13539, n13540, n13541, n13542, n13543, n13544, n13545,
         n13546, n13547, n13548, n13549, n13550, n13551, n13552, n13553,
         n13554, n13555, n13556, n13557, n13558, n13559, n13560, n13561,
         n13562, n13563, n13564, n13565, n13566, n13567, n13568, n13569,
         n13570, n13571, n13572, n13573, n13574, n13575, n13576, n13577,
         n13578, n13579, n13580, n13581, n13582, n13583, n13584, n13585,
         n13586, n13587, n13588, n13589, n13590, n13591, n13592, n13593,
         n13594, n13595, n13596, n13597, n13598, n13599, n13600, n13601,
         n13602, n13603, n13604, n13605, n13606, n13607, n13608, n13609,
         n13610, n13611, n13612, n13613, n13614, n13615, n13616, n13617,
         n13618, n13619, n13620, n13621, n13622, n13623, n13624, n13625,
         n13626, n13627, n13628, n13629, n13630, n13631, n13632, n13633,
         n13634, n13635, n13636, n13637, n13638, n13639, n13640, n13641,
         n13642, n13643, n13644, n13645, n13646, n13647, n13648, n13649,
         n13650, n13651, n13652, n13653, n13654, n13655, n13656, n13657,
         n13658, n13659, n13660, n13661, n13662, n13663, n13664, n13665,
         n13666, n13667, n13668, n13669, n13670, n13671, n13672, n13673,
         n13674, n13675, n13676, n13677, n13678, n13679, n13680, n13681,
         n13682, n13683, n13684, n13685, n13686, n13687, n13688, n13689,
         n13690, n13691, n13692, n13693, n13694, n13695, n13696, n13697,
         n13698, n13699, n13700, n13701, n13702, n13703, n13704, n13705,
         n13706, n13707, n13708, n13709, n13710, n13711, n13712, n13713,
         n13714, n13715, n13716, n13717, n13718, n13719, n13720, n13721,
         n13722, n13723, n13724, n13725, n13726, n13727, n13728, n13729,
         n13730, n13731, n13732, n13733, n13734, n13735, n13736, n13737,
         n13738, n13739, n13740, n13741, n13742, n13743, n13744, n13745,
         n13746, n13747, n13748, n13749, n13750, n13751, n13752, n13753,
         n13754, n13755, n13756, n13757, n13758, n13759, n13760, n13761,
         n13762, n13763, n13764, n13765, n13766, n13767, n13768, n13769,
         n13770, n13771, n13772, n13773, n13774, n13775, n13776, n13777,
         n13778, n13779, n13780, n13781, n13782, n13783, n13784, n13785,
         n13786, n13787, n13788, n13789, n13790, n13791, n13792, n13793,
         n13794, n13795, n13796, n13797, n13798, n13799, n13800, n13801,
         n13802, n13803, n13804, n13805, n13806, n13807, n13808, n13809,
         n13810, n13811, n13812, n13813, n13814, n13815, n13816, n13817,
         n13818, n13819, n13820, n13821, n13822, n13823, n13824, n13825,
         n13826, n13827, n13828, n13829, n13830, n13831, n13832, n13833,
         n13834, n13835, n13836, n13837, n13838, n13839, n13840, n13841,
         n13842, n13843, n13844, n13845, n13846, n13847, n13848, n13849,
         n13850, n13851, n13852, n13853, n13854, n13855, n13856, n13857,
         n13858, n13859, n13860, n13861, n13862, n13863, n13864, n13865,
         n13866, n13867, n13868, n13869, n13870, n13871, n13872, n13873,
         n13874, n13875, n13876, n13877, n13878, n13879, n13880, n13881,
         n13882, n13883, n13884, n13885, n13886, n13887, n13888, n13889,
         n13890, n13891, n13892, n13893, n13894, n13895, n13896, n13897,
         n13898, n13899, n13900, n13901, n13902, n13903, n13904, n13905,
         n13906, n13907, n13908, n13909, n13910, n13911, n13912, n13913,
         n13914, n13915, n13916, n13917, n13918, n13919, n13920, n13921,
         n13922, n13923, n13924, n13925, n13926, n13927, n13928, n13929,
         n13930, n13931, n13932, n13933, n13934, n13935, n13936, n13937,
         n13938, n13939, n13940, n13941, n13942, n13943, n13944, n13945,
         n13946, n13947, n13948, n13949, n13950, n13951, n13952, n13953,
         n13954, n13955, n13956, n13957, n13958, n13959, n13960, n13961,
         n13962, n13963, n13964, n13965, n13966, n13967, n13968, n13969,
         n13970, n13971, n13972, n13973, n13974, n13975, n13976, n13977,
         n13978, n13979, n13980, n13981, n13982, n13983, n13984, n13985,
         n13986, n13987, n13988, n13989, n13990, n13991, n13992, n13993,
         n13994, n13995, n13996, n13997, n13998, n13999, n14000, n14001,
         n14002, n14003, n14004, n14005, n14006, n14007, n14008, n14009,
         n14010, n14011, n14012, n14013, n14014, n14015, n14016, n14017,
         n14018, n14019, n14020, n14021, n14022, n14023, n14024, n14025,
         n14026, n14027, n14028, n14029, n14030, n14031, n14032, n14033,
         n14034, n14035, n14036, n14037, n14038, n14039, n14040, n14041,
         n14042, n14043, n14044, n14045, n14046, n14047, n14048, n14049,
         n14050, n14051, n14052, n14053, n14054, n14055, n14056, n14057,
         n14058, n14059, n14060, n14061, n14062, n14063, n14064, n14065,
         n14066, n14067, n14068, n14069, n14070, n14071, n14072, n14073,
         n14074, n14075, n14076, n14077, n14078, n14079, n14080, n14081,
         n14082, n14083, n14084, n14085, n14086, n14087, n14088, n14089,
         n14090, n14091, n14092, n14093, n14094, n14095, n14096, n14097,
         n14098, n14099, n14100, n14101, n14102, n14103, n14104, n14105,
         n14106, n14107, n14108, n14109, n14110, n14111, n14112, n14113,
         n14114, n14115, n14116, n14117, n14118, n14119, n14120, n14121,
         n14122, n14123, n14124, n14125, n14126, n14127, n14128, n14129,
         n14130, n14131, n14132, n14133, n14134, n14135, n14136, n14137,
         n14138, n14139, n14140, n14141, n14142, n14143, n14144, n14145,
         n14146, n14147, n14148, n14149, n14150, n14151, n14152, n14153,
         n14154, n14155, n14156, n14157, n14158, n14159, n14160, n14161,
         n14162, n14163, n14164, n14165, n14166, n14167, n14168, n14169,
         n14170, n14171, n14172, n14173, n14174, n14175, n14176, n14177,
         n14178, n14179, n14180, n14181, n14182, n14183, n14184, n14185,
         n14186, n14187, n14188, n14189, n14190, n14191, n14192, n14193,
         n14194, n14195, n14196, n14197, n14198, n14199, n14200, n14201,
         n14202, n14203, n14204, n14205, n14206, n14207, n14208, n14209,
         n14210, n14211, n14212, n14213, n14214, n14215, n14216, n14217,
         n14218, n14219, n14220, n14221, n14222, n14223, n14224, n14225,
         n14226, n14227, n14228, n14229, n14230, n14231, n14232, n14233,
         n14234, n14235, n14236, n14237, n14238, n14239, n14240, n14241,
         n14242, n14243, n14244, n14245, n14246, n14247, n14248, n14249,
         n14250, n14251, n14252, n14253, n14254, n14255, n14256, n14257,
         n14258, n14259, n14260, n14261, n14262, n14263, n14264, n14265,
         n14266, n14267, n14268, n14269, n14270, n14271, n14272, n14273,
         n14274, n14275, n14276, n14277, n14278, n14279, n14280, n14281,
         n14282, n14283, n14284, n14285, n14286, n14287, n14288, n14289,
         n14290, n14291, n14292, n14293, n14294, n14295, n14296, n14297,
         n14298, n14299, n14300, n14301, n14302, n14303, n14304, n14305,
         n14306, n14307, n14308, n14309, n14310, n14311, n14312, n14313,
         n14314, n14315, n14316, n14317, n14318, n14319, n14320, n14321,
         n14322, n14323, n14324, n14325, n14326, n14327, n14328, n14329,
         n14330, n14331, n14332, n14333, n14334, n14335, n14336, n14337,
         n14338, n14339, n14340, n14341, n14342, n14343, n14344, n14345,
         n14346, n14347, n14348, n14349, n14350, n14351, n14352, n14353,
         n14354, n14355, n14356, n14357, n14358, n14359, n14360, n14361,
         n14362, n14363, n14364, n14365, n14366, n14367, n14368, n14369,
         n14370, n14371, n14372, n14373, n14374, n14375, n14376, n14377,
         n14378, n14379, n14380, n14381, n14382, n14383, n14384, n14385,
         n14386, n14387, n14388, n14389, n14390, n14391, n14392, n14393,
         n14394, n14395, n14396, n14397, n14398, n14399, n14400, n14401,
         n14402, n14403, n14404, n14405, n14406, n14407, n14408, n14409,
         n14410, n14411, n14412, n14413, n14414, n14415, n14416, n14417,
         n14418, n14419, n14420, n14421, n14422, n14423, n14424, n14425,
         n14426, n14427, n14428, n14429, n14430, n14431, n14432, n14433,
         n14434, n14435, n14436, n14437, n14438, n14439, n14440, n14441,
         n14442, n14443, n14444, n14445, n14446, n14447, n14448, n14449,
         n14450, n14451, n14452, n14453, n14454, n14455, n14456, n14457,
         n14458, n14459, n14460, n14461, n14462, n14463, n14464, n14465,
         n14466, n14467, n14468, n14469, n14470, n14471, n14472, n14473,
         n14474, n14475, n14476, n14477, n14478, n14479, n14480, n14481,
         n14482, n14483, n14484, n14485, n14486, n14487, n14488, n14489,
         n14490, n14491, n14492, n14493, n14494, n14495, n14496, n14497,
         n14498, n14499, n14500, n14501, n14502, n14503, n14504, n14505,
         n14506, n14507, n14508, n14509, n14510, n14511, n14512, n14513,
         n14514, n14515, n14516, n14517, n14518, n14519, n14520, n14521,
         n14522, n14523, n14524, n14525, n14526, n14527, n14528, n14529,
         n14530, n14531, n14532, n14533, n14534, n14535, n14536, n14537,
         n14538, n14539, n14540, n14541, n14542, n14543, n14544, n14545,
         n14546, n14547, n14548, n14549, n14550, n14551, n14552, n14553,
         n14554, n14555, n14556, n14557, n14558, n14559, n14560, n14561,
         n14562, n14563, n14564, n14565, n14566, n14567, n14568, n14569,
         n14570, n14571, n14572, n14573, n14574, n14575, n14576, n14577,
         n14578, n14579, n14580, n14581, n14582, n14583, n14584, n14585,
         n14586, n14587, n14588, n14589, n14590, n14591, n14592, n14593,
         n14594, n14595, n14596, n14597, n14598, n14599, n14600, n14601,
         n14602, n14603, n14604, n14605, n14606, n14607, n14608, n14609,
         n14610, n14611, n14612, n14613, n14614, n14615, n14616, n14617,
         n14618, n14619, n14620, n14621, n14622, n14623, n14624, n14625,
         n14626, n14627, n14628, n14629, n14630, n14631, n14632, n14633,
         n14634, n14635, n14636, n14637, n14638, n14639, n14640, n14641,
         n14642, n14643, n14644, n14645, n14646, n14647, n14648, n14649,
         n14650, n14651, n14652, n14653, n14654, n14655, n14656, n14657,
         n14658, n14659, n14660, n14661, n14662, n14663, n14664, n14665,
         n14666, n14667, n14668, n14669, n14670, n14671, n14672, n14673,
         n14674, n14675, n14676, n14677, n14678, n14679, n14680, n14681,
         n14682, n14683, n14684, n14685, n14686, n14687, n14688, n14689,
         n14690, n14691, n14692, n14693, n14694, n14695, n14696, n14697,
         n14698, n14699, n14700, n14701, n14702, n14703, n14704, n14705,
         n14706, n14707, n14708, n14709, n14710, n14711, n14712, n14713,
         n14714, n14715, n14716, n14717, n14718, n14719, n14720, n14721,
         n14722, n14723, n14724, n14725, n14726, n14727, n14728, n14729,
         n14730, n14731, n14732, n14733, n14734, n14735, n14736, n14737,
         n14738, n14739, n14740, n14741, n14742, n14743, n14744, n14745,
         n14746, n14747, n14748, n14749, n14750, n14751, n14752, n14753,
         n14754, n14755, n14756, n14757, n14758, n14759, n14760, n14761,
         n14762, n14763, n14764, n14765, n14766, n14767, n14768, n14769,
         n14770, n14771, n14772, n14773, n14774, n14775, n14776, n14777,
         n14778, n14779, n14780, n14781, n14782, n14783, n14784, n14785,
         n14786, n14787, n14788, n14789, n14790, n14791, n14792, n14793,
         n14794, n14795, n14796, n14797, n14798, n14799, n14800, n14801,
         n14802, n14803, n14804, n14805, n14806, n14807, n14808, n14809,
         n14810, n14811, n14812, n14813, n14814, n14815, n14816, n14817,
         n14818, n14819, n14820, n14821, n14822, n14823, n14824, n14825,
         n14826, n14827, n14828, n14829, n14830, n14831, n14832, n14833,
         n14834, n14835, n14836, n14837, n14838, n14839, n14840, n14841,
         n14842, n14843, n14844, n14845, n14846, n14847, n14848, n14849,
         n14850, n14851, n14852, n14853, n14854, n14855, n14856, n14857,
         n14858, n14859, n14860, n14861, n14862, n14863, n14864, n14865,
         n14866, n14867, n14868, n14869, n14870, n14871, n14872, n14873,
         n14874, n14875, n14876, n14877, n14878, n14879, n14880, n14881,
         n14882, n14883, n14884, n14885, n14886, n14887, n14888, n14889,
         n14890, n14891, n14892, n14893, n14894, n14895, n14896, n14897,
         n14898, n14899, n14900, n14901, n14902, n14903, n14904, n14905,
         n14906, n14907, n14908, n14909, n14910, n14911, n14912, n14913,
         n14914, n14915, n14916, n14917, n14918, n14919, n14920, n14921,
         n14922, n14923, n14924, n14925, n14926, n14927, n14928, n14929,
         n14930, n14931, n14932, n14933, n14934, n14935, n14936, n14937,
         n14938, n14939, n14940, n14941, n14942, n14943, n14944, n14945,
         n14946, n14947, n14948, n14949, n14950, n14951, n14952, n14953,
         n14954, n14955, n14956, n14957, n14958, n14959, n14960, n14961,
         n14962, n14963, n14964, n14965, n14966, n14967, n14968, n14969,
         n14970, n14971, n14972, n14973, n14974, n14975, n14976, n14977,
         n14978, n14979, n14980, n14981, n14982, n14983, n14984, n14985,
         n14986, n14987, n14988, n14989, n14990, n14991, n14992, n14993,
         n14994, n14995, n14996, n14997, n14998, n14999, n15000, n15001,
         n15002, n15003, n15004, n15005, n15006, n15007, n15008, n15009,
         n15010, n15011, n15012, n15013, n15014, n15015, n15016, n15017,
         n15018, n15019, n15020, n15021, n15022, n15023, n15024, n15025,
         n15026, n15027, n15028, n15029, n15030, n15031, n15032, n15033,
         n15034, n15035, n15036, n15037, n15038, n15039, n15040, n15041,
         n15042, n15043, n15044, n15045, n15046, n15047, n15048, n15049,
         n15050, n15051, n15052, n15053, n15054, n15055, n15056, n15057,
         n15058, n15059, n15060, n15061, n15062, n15063, n15064, n15065,
         n15066, n15067, n15068, n15069, n15070, n15071, n15072, n15073,
         n15074, n15075, n15076, n15077, n15078, n15079, n15080, n15081,
         n15082, n15083, n15084, n15085, n15086, n15087, n15088, n15089,
         n15090, n15091, n15092, n15093, n15094, n15095, n15096, n15097,
         n15098, n15099, n15100, n15101, n15102, n15103, n15104, n15105,
         n15106, n15107, n15108, n15109, n15110, n15111, n15112, n15113,
         n15114, n15115, n15116, n15117, n15118, n15119, n15120, n15121,
         n15122, n15123, n15124, n15125, n15126, n15127, n15128, n15129,
         n15130, n15131, n15132, n15133, n15134, n15135, n15136, n15137,
         n15138, n15139, n15140, n15141, n15142, n15143, n15144, n15145,
         n15146, n15147, n15148, n15149, n15150, n15151, n15152, n15153,
         n15154, n15155, n15156, n15157, n15158, n15159, n15160, n15161,
         n15162, n15163, n15164, n15165, n15166, n15167, n15168, n15169,
         n15170, n15171, n15172, n15173, n15174, n15175, n15176, n15177,
         n15178, n15179, n15180, n15181, n15182, n15183, n15184, n15185,
         n15186, n15187, n15188, n15189, n15190, n15191, n15192, n15193,
         n15194, n15195, n15196, n15197, n15198, n15199, n15200, n15201,
         n15202, n15203, n15204, n15205, n15206, n15207, n15208, n15209,
         n15210, n15211, n15212, n15213, n15214, n15215, n15216, n15217,
         n15218, n15219, n15220, n15221, n15222, n15223, n15224, n15225,
         n15226, n15227, n15228, n15229, n15230, n15231, n15232, n15233,
         n15234, n15235, n15236, n15237, n15238, n15239, n15240, n15241,
         n15242, n15243, n15244, n15245, n15246, n15247, n15248, n15249,
         n15250, n15251, n15252, n15253, n15254, n15255, n15256, n15257,
         n15258, n15259, n15260, n15261, n15262, n15263, n15264, n15265,
         n15266, n15267, n15268, n15269, n15270, n15271, n15272, n15273,
         n15274, n15275, n15276, n15277, n15278, n15279, n15280, n15281,
         n15282, n15283, n15284, n15285, n15286, n15287, n15288, n15289,
         n15290, n15291, n15292, n15293, n15294, n15295, n15296, n15297,
         n15298, n15299, n15300, n15301, n15302, n15303, n15304, n15305,
         n15306, n15307, n15308, n15309, n15310, n15311, n15312, n15313,
         n15314, n15315, n15316, n15317, n15318, n15319, n15320, n15321,
         n15322, n15323, n15324, n15325, n15326, n15327, n15328, n15329,
         n15330, n15331, n15332, n15333, n15334, n15335, n15336, n15337,
         n15338, n15339, n15340, n15341, n15342, n15343, n15344, n15345,
         n15346, n15347, n15348, n15349, n15350, n15351, n15352, n15353,
         n15354, n15355, n15356, n15357, n15358, n15359, n15360, n15361,
         n15362, n15363, n15364, n15365, n15366, n15367, n15368, n15369,
         n15370, n15371, n15372, n15373, n15374, n15375, n15376, n15377,
         n15378, n15379, n15380, n15381, n15382, n15383, n15384, n15385,
         n15386, n15387, n15388, n15389, n15390, n15391, n15392, n15393,
         n15394, n15395, n15396, n15397, n15398, n15399, n15400, n15401,
         n15402, n15403, n15404, n15405, n15406, n15407, n15408, n15409,
         n15410, n15411, n15412, n15413, n15414, n15415, n15416, n15417,
         n15418, n15419, n15420, n15421, n15422, n15423, n15424, n15425,
         n15426, n15427, n15428, n15429, n15430, n15431, n15432, n15433,
         n15434, n15435, n15436, n15437, n15438, n15439, n15440, n15441,
         n15442, n15443, n15444, n15445, n15446, n15447, n15448, n15449,
         n15450, n15451, n15452, n15453, n15454, n15455, n15456, n15457,
         n15458, n15459, n15460, n15461, n15462, n15463, n15464, n15465,
         n15466, n15467, n15468, n15469, n15470, n15471, n15472, n15473,
         n15474, n15475, n15476, n15477, n15478, n15479, n15480, n15481,
         n15482, n15483, n15484, n15485, n15486, n15487, n15488, n15489,
         n15490, n15491, n15492, n15493, n15494, n15495, n15496, n15497,
         n15498, n15499, n15500, n15501, n15502, n15503, n15504, n15505,
         n15506, n15507, n15508, n15509, n15510, n15511, n15512, n15513,
         n15514, n15515, n15516, n15517, n15518, n15519, n15520, n15521,
         n15522, n15523, n15524, n15525, n15526, n15527, n15528, n15529,
         n15530, n15531, n15532, n15533, n15534, n15535, n15536, n15537,
         n15538, n15539, n15540, n15541, n15542, n15543, n15544, n15545,
         n15546, n15547, n15548, n15549, n15550, n15551, n15552, n15553,
         n15554, n15555, n15556, n15557, n15558, n15559, n15560, n15561,
         n15562, n15563, n15564, n15565, n15566, n15567, n15568, n15569,
         n15570, n15571, n15572, n15573, n15574, n15575, n15576, n15577,
         n15578, n15579, n15580, n15581, n15582, n15583, n15584, n15585,
         n15586, n15587, n15588, n15589, n15590, n15591, n15592, n15593,
         n15594, n15595, n15596, n15597, n15598, n15599, n15600, n15601,
         n15602, n15603, n15604, n15605, n15606, n15607, n15608, n15609,
         n15610, n15611, n15612, n15613, n15614, n15615, n15616, n15617,
         n15618, n15619, n15620, n15621, n15622, n15623, n15624, n15625,
         n15626, n15627, n15628, n15629, n15630, n15631, n15632, n15633,
         n15634, n15635, n15636, n15637, n15638, n15639, n15640, n15641,
         n15642, n15643, n15644, n15645, n15646, n15647, n15648, n15649,
         n15650, n15651, n15652, n15653, n15654, n15655, n15656, n15657,
         n15658, n15659, n15660, n15661, n15662, n15663, n15664, n15665,
         n15666, n15667, n15668, n15669, n15670, n15671, n15672, n15673,
         n15674, n15675, n15676, n15677, n15678, n15679, n15680, n15681,
         n15682, n15683, n15684, n15685, n15686, n15687, n15688, n15689,
         n15690, n15691, n15692, n15693, n15694, n15695, n15696, n15697,
         n15698, n15699, n15700, n15701, n15702, n15703, n15704, n15705,
         n15706, n15707, n15708, n15709, n15710, n15711, n15712, n15713,
         n15714, n15715, n15716, n15717, n15718, n15719, n15720, n15721,
         n15722, n15723, n15724, n15725, n15726, n15727, n15728, n15729,
         n15730, n15731, n15732, n15733, n15734, n15735, n15736, n15737,
         n15738, n15739, n15740, n15741, n15742, n15743, n15744, n15745,
         n15746, n15747, n15748, n15749, n15750, n15751, n15752, n15753,
         n15754, n15755, n15756, n15757, n15758, n15759, n15760, n15761,
         n15762, n15763, n15764, n15765, n15766, n15767, n15768, n15769,
         n15770, n15771, n15772, n15773, n15774, n15775, n15776, n15777,
         n15778, n15779, n15780, n15781, n15782, n15783, n15784, n15785,
         n15786, n15787, n15788, n15789, n15790, n15791, n15792, n15793,
         n15794, n15795, n15796, n15797, n15798, n15799, n15800, n15801,
         n15802, n15803, n15804, n15805, n15806, n15807, n15808, n15809,
         n15810, n15811, n15812, n15813, n15814, n15815, n15816, n15817,
         n15818, n15819, n15820, n15821, n15822, n15823, n15824, n15825,
         n15826, n15827, n15828, n15829, n15830, n15831, n15832, n15833,
         n15834, n15835, n15836, n15837, n15838, n15839, n15840, n15841,
         n15842, n15843, n15844, n15845, n15846, n15847, n15848, n15849,
         n15850, n15851, n15852, n15853, n15854, n15855, n15856, n15857,
         n15858, n15859, n15860, n15861, n15862, n15863, n15864, n15865,
         n15866, n15867, n15868, n15869, n15870, n15871, n15872, n15873,
         n15874, n15875, n15876, n15877, n15878, n15879, n15880, n15881,
         n15882, n15883, n15884, n15885, n15886, n15887, n15888, n15889,
         n15890, n15891, n15892, n15893, n15894, n15895, n15896, n15897,
         n15898, n15899, n15900, n15901, n15902, n15903, n15904, n15905,
         n15906, n15907, n15908, n15909, n15910, n15911, n15912, n15913,
         n15914, n15915, n15916, n15917, n15918, n15919, n15920, n15921,
         n15922, n15923, n15924, n15925, n15926, n15927, n15928, n15929,
         n15930, n15931, n15932, n15933, n15934, n15935, n15936, n15937,
         n15938, n15939, n15940, n15941, n15942, n15943, n15944, n15945,
         n15946, n15947, n15948, n15949, n15950, n15951, n15952, n15953,
         n15954, n15955, n15956, n15957, n15958, n15959, n15960, n15961,
         n15962, n15963, n15964, n15965, n15966, n15967, n15968, n15969,
         n15970, n15971, n15972, n15973, n15974, n15975, n15976, n15977,
         n15978, n15979, n15980, n15981, n15982, n15983, n15984, n15985,
         n15986, n15987, n15988, n15989, n15990, n15991, n15992, n15993,
         n15994, n15995, n15996, n15997, n15998, n15999, n16000, n16001,
         n16002, n16003, n16004, n16005, n16006, n16007, n16008, n16009,
         n16010, n16011, n16012, n16013, n16014, n16015, n16016, n16017,
         n16018, n16019, n16020, n16021, n16022, n16023, n16024, n16025,
         n16026, n16027, n16028, n16029, n16030, n16031, n16032, n16033,
         n16034, n16035, n16036, n16037, n16038, n16039, n16040, n16041,
         n16042, n16043, n16044, n16045, n16046, n16047, n16048, n16049,
         n16050, n16051, n16052, n16053, n16054, n16055, n16056, n16057,
         n16058, n16059, n16060, n16061, n16062, n16063, n16064, n16065,
         n16066, n16067, n16068, n16069, n16070, n16071, n16072, n16073,
         n16074, n16075, n16076, n16077, n16078, n16079, n16080, n16081,
         n16082, n16083, n16084, n16085, n16086, n16087, n16088, n16089,
         n16090, n16091, n16092, n16093, n16094, n16095, n16096, n16097,
         n16098, n16099, n16100, n16101, n16102, n16103, n16104, n16105,
         n16106, n16107, n16108, n16109, n16110, n16111, n16112, n16113,
         n16114, n16115, n16116, n16117, n16118, n16119, n16120, n16121,
         n16122, n16123, n16124, n16125, n16126, n16127, n16128, n16129,
         n16130, n16131, n16132, n16133, n16134, n16135, n16136, n16137,
         n16138, n16139, n16140, n16141, n16142, n16143, n16144, n16145,
         n16146, n16147, n16148, n16149, n16150, n16151, n16152, n16153,
         n16154, n16155, n16156, n16157, n16158, n16159, n16160, n16161,
         n16162, n16163, n16164, n16165, n16166, n16167, n16168, n16169,
         n16170, n16171, n16172, n16173, n16174, n16175, n16176, n16177,
         n16178, n16179, n16180, n16181, n16182, n16183, n16184, n16185,
         n16186, n16187, n16188, n16189, n16190, n16191, n16192, n16193,
         n16194, n16195, n16196, n16197, n16198, n16199, n16200, n16201,
         n16202, n16203, n16204, n16205, n16206, n16207, n16208, n16209,
         n16210, n16211, n16212, n16213, n16214, n16215, n16216, n16217,
         n16218, n16219, n16220, n16221, n16222, n16223, n16224, n16225,
         n16226, n16227, n16228, n16229, n16230, n16231, n16232, n16233,
         n16234, n16235, n16236, n16237, n16238, n16239, n16240, n16241,
         n16242, n16243, n16244, n16245, n16246, n16247, n16248, n16249,
         n16250, n16251, n16252, n16253, n16254, n16255, n16256, n16257,
         n16258, n16259, n16260, n16261, n16262, n16263, n16264, n16265,
         n16266, n16267, n16268, n16269, n16270, n16271, n16272, n16273,
         n16274, n16275, n16276, n16277, n16278, n16279, n16280, n16281,
         n16282, n16283, n16284, n16285, n16286, n16287, n16288, n16289,
         n16290, n16291, n16292, n16293, n16294, n16295, n16296, n16297,
         n16298, n16299, n16300, n16301, n16302, n16303, n16304, n16305,
         n16306, n16307, n16308, n16309, n16310, n16311, n16312, n16313,
         n16314, n16315, n16316, n16317, n16318, n16319, n16320, n16321,
         n16322, n16323, n16324, n16325, n16326, n16327, n16328, n16329,
         n16330, n16331, n16332, n16333, n16334, n16335, n16336, n16337,
         n16338, n16339, n16340, n16341, n16342, n16343, n16344, n16345,
         n16346, n16347, n16348, n16349, n16350, n16351, n16352, n16353,
         n16354, n16355, n16356, n16357, n16358, n16359, n16360, n16361,
         n16362, n16363, n16364, n16365, n16366, n16367, n16368, n16369,
         n16370, n16371, n16372, n16373, n16374, n16375, n16376, n16377,
         n16378, n16379, n16380, n16381, n16382, n16383, n16384, n16385,
         n16386, n16387, n16388, n16389, n16390, n16391, n16392, n16393,
         n16394, n16395, n16396, n16397, n16398, n16399, n16400, n16401,
         n16402, n16403, n16404, n16405, n16406, n16407, n16408, n16409,
         n16410, n16411, n16412, n16413, n16414, n16415, n16416, n16417,
         n16418, n16419, n16420, n16421, n16422, n16423, n16424, n16425,
         n16426, n16427, n16428, n16429, n16430, n16431, n16432, n16433,
         n16434, n16435, n16436, n16437, n16438, n16439, n16440, n16441,
         n16442, n16443, n16444, n16445, n16446, n16447, n16448, n16449,
         n16450, n16451, n16452, n16453, n16454, n16455, n16456, n16457,
         n16458, n16459, n16460, n16461, n16462, n16463, n16464, n16465,
         n16466, n16467, n16468, n16469, n16470, n16471, n16472, n16473,
         n16474, n16475, n16476, n16477, n16478, n16479, n16480, n16481,
         n16482, n16483, n16484, n16485, n16486, n16487, n16488, n16489,
         n16490, n16491, n16492, n16493, n16494, n16495, n16496, n16497,
         n16498, n16499, n16500, n16501, n16502, n16503, n16504, n16505,
         n16506, n16507, n16508, n16509, n16510, n16511, n16512, n16513,
         n16514, n16515, n16516, n16517, n16518, n16519, n16520, n16521,
         n16522, n16523, n16524, n16525, n16526, n16527, n16528, n16529,
         n16530, n16531, n16532, n16533, n16534, n16535, n16536, n16537,
         n16538, n16539, n16540, n16541, n16542, n16543, n16544, n16545,
         n16546, n16547, n16548, n16549, n16550, n16551, n16552, n16553,
         n16554, n16555, n16556, n16557, n16558, n16559, n16560, n16561,
         n16562, n16563, n16564, n16565, n16566, n16567, n16568, n16569,
         n16570, n16571, n16572, n16573, n16574, n16575, n16576, n16577,
         n16578, n16579, n16580, n16581, n16582, n16583, n16584, n16585,
         n16586, n16587, n16588, n16589, n16590, n16591, n16592, n16593,
         n16594, n16595, n16596, n16597, n16598, n16599, n16600, n16601,
         n16602, n16603, n16604, n16605, n16606, n16607, n16608, n16609,
         n16610, n16611, n16612, n16613, n16614, n16615, n16616, n16617,
         n16618, n16619, n16620, n16621, n16622, n16623, n16624, n16625,
         n16626, n16627, n16628, n16629, n16630, n16631, n16632, n16633,
         n16634, n16635, n16636, n16637, n16638, n16639, n16640, n16641,
         n16642, n16643, n16644, n16645, n16646, n16647, n16648, n16649,
         n16650, n16651, n16652, n16653, n16654, n16655, n16656, n16657,
         n16658, n16659, n16660, n16661, n16662, n16663, n16664, n16665,
         n16666, n16667, n16668, n16669, n16670, n16671, n16672, n16673,
         n16674, n16675, n16676, n16677, n16678, n16679, n16680, n16681,
         n16682, n16683, n16684, n16685, n16686, n16687, n16688, n16689,
         n16690, n16691, n16692, n16693, n16694, n16695, n16696, n16697,
         n16698, n16699, n16700, n16701, n16702, n16703, n16704, n16705,
         n16706, n16707, n16708, n16709, n16710, n16711, n16712, n16713,
         n16714, n16715, n16716, n16717, n16718, n16719, n16720, n16721,
         n16722, n16723, n16724, n16725, n16726, n16727, n16728, n16729,
         n16730, n16731, n16732, n16733, n16734, n16735, n16736, n16737,
         n16738, n16739, n16740, n16741, n16742, n16743, n16744, n16745,
         n16746, n16747, n16748, n16749, n16750, n16751, n16752, n16753,
         n16754, n16755, n16756, n16757, n16758, n16759, n16760, n16761,
         n16762, n16763, n16764, n16765, n16766, n16767, n16768, n16769,
         n16770, n16771, n16772, n16773, n16774, n16775, n16776, n16777,
         n16778, n16779, n16780, n16781, n16782, n16783, n16784, n16785,
         n16786, n16787, n16788, n16789, n16790, n16791, n16792, n16793,
         n16794, n16795, n16796, n16797, n16798, n16799, n16800, n16801,
         n16802, n16803, n16804, n16805, n16806, n16807, n16808, n16809,
         n16810, n16811, n16812, n16813, n16814, n16815, n16816, n16817,
         n16818, n16819, n16820, n16821, n16822, n16823, n16824, n16825,
         n16826, n16827, n16828, n16829, n16830, n16831, n16832, n16833,
         n16834, n16835, n16836, n16837, n16838, n16839, n16840, n16841,
         n16842, n16843, n16844, n16845, n16846, n16847, n16848, n16849,
         n16850, n16851, n16852, n16853, n16854, n16855, n16856, n16857,
         n16858, n16859, n16860, n16861, n16862, n16863, n16864, n16865,
         n16866, n16867, n16868, n16869, n16870, n16871, n16872, n16873,
         n16874, n16875, n16876, n16877, n16878, n16879, n16880, n16881,
         n16882, n16883, n16884, n16885, n16886, n16887, n16888, n16889,
         n16890, n16891, n16892, n16893, n16894, n16895, n16896, n16897,
         n16898, n16899, n16900, n16901, n16902, n16903, n16904, n16905,
         n16906, n16907, n16908, n16909, n16910, n16911, n16912, n16913,
         n16914, n16915, n16916, n16917, n16918, n16919, n16920, n16921,
         n16922, n16923, n16924, n16925, n16926, n16927, n16928, n16929,
         n16930, n16931, n16932, n16933, n16934, n16935, n16936, n16937,
         n16938, n16939, n16940, n16941, n16942, n16943, n16944, n16945,
         n16946, n16947, n16948, n16949, n16950, n16951, n16952, n16953,
         n16954, n16955, n16956, n16957, n16958, n16959, n16960, n16961,
         n16962, n16963, n16964, n16965, n16966, n16967, n16968, n16969,
         n16970, n16971, n16972, n16973, n16974, n16975, n16976, n16977,
         n16978, n16979, n16980, n16981, n16982, n16983, n16984, n16985,
         n16986, n16987, n16988, n16989, n16990, n16991, n16992, n16993,
         n16994, n16995, n16996, n16997, n16998, n16999, n17000, n17001,
         n17002, n17003, n17004, n17005, n17006, n17007, n17008, n17009,
         n17010, n17011, n17012, n17013, n17014, n17015, n17016, n17017,
         n17018, n17019, n17020, n17021, n17022, n17023, n17024, n17025,
         n17026, n17027, n17028, n17029, n17030, n17031, n17032, n17033,
         n17034, n17035, n17036, n17037, n17038, n17039, n17040, n17041,
         n17042, n17043, n17044, n17045, n17046, n17047, n17048, n17049,
         n17050, n17051, n17052, n17053, n17054, n17055, n17056, n17057,
         n17058, n17059, n17060, n17061, n17062, n17063, n17064, n17065,
         n17066, n17067, n17068, n17069, n17070, n17071, n17072, n17073,
         n17074, n17075, n17076, n17077, n17078, n17079, n17080, n17081,
         n17082, n17083, n17084, n17085, n17086, n17087, n17088, n17089,
         n17090, n17091, n17092, n17093, n17094, n17095, n17096, n17097,
         n17098, n17099, n17100, n17101, n17102, n17103, n17104, n17105,
         n17106, n17107, n17108, n17109, n17110, n17111, n17112, n17113,
         n17114, n17115, n17116, n17117, n17118, n17119, n17120, n17121,
         n17122, n17123, n17124, n17125, n17126, n17127, n17128, n17129,
         n17130, n17131, n17132, n17133, n17134, n17135, n17136, n17137,
         n17138, n17139, n17140, n17141, n17142, n17143, n17144, n17145,
         n17146, n17147, n17148, n17149, n17150, n17151, n17152, n17153,
         n17154, n17155, n17156, n17157, n17158, n17159, n17160, n17161,
         n17162, n17163, n17164, n17165, n17166, n17167, n17168, n17169,
         n17170, n17171, n17172, n17173, n17174, n17175, n17176, n17177,
         n17178, n17179, n17180, n17181, n17182, n17183, n17184, n17185,
         n17186, n17187, n17188, n17189, n17190, n17191, n17192, n17193,
         n17194, n17195, n17196, n17197, n17198, n17199, n17200, n17201,
         n17202, n17203, n17204, n17205, n17206, n17207, n17208, n17209,
         n17210, n17211, n17212, n17213, n17214, n17215, n17216, n17217,
         n17218, n17219, n17220, n17221, n17222, n17223, n17224, n17225,
         n17226, n17227, n17228, n17229, n17230, n17231, n17232, n17233,
         n17234, n17235, n17236, n17237, n17238, n17239, n17240, n17241,
         n17242, n17243, n17244, n17245, n17246, n17247, n17248, n17249,
         n17250, n17251, n17252, n17253, n17254, n17255, n17256, n17257,
         n17258, n17259, n17260, n17261, n17262, n17263, n17264, n17265,
         n17266, n17267, n17268, n17269, n17270, n17271, n17272, n17273,
         n17274, n17275, n17276, n17277, n17278, n17279, n17280, n17281,
         n17282, n17283, n17284, n17285, n17286, n17287, n17288, n17289,
         n17290, n17291, n17292, n17293, n17294, n17295, n17296, n17297,
         n17298, n17299, n17300, n17301, n17302, n17303, n17304, n17305,
         n17306, n17307, n17308, n17309, n17310, n17311, n17312, n17313,
         n17314, n17315, n17316, n17317, n17318, n17319, n17320, n17321,
         n17322, n17323, n17324, n17325, n17326, n17327, n17328, n17329,
         n17330, n17331, n17332, n17333, n17334, n17335, n17336, n17337,
         n17338, n17339, n17340, n17341, n17342, n17343, n17344, n17345,
         n17346, n17347, n17348, n17349, n17350, n17351, n17352, n17353,
         n17354, n17355, n17356, n17357, n17358, n17359, n17360, n17361,
         n17362, n17363, n17364, n17365, n17366, n17367, n17368, n17369,
         n17370, n17371, n17372, n17373, n17374, n17375, n17376, n17377,
         n17378, n17379, n17380, n17381, n17382, n17383, n17384, n17385,
         n17386, n17387, n17388, n17389, n17390, n17391, n17392, n17393,
         n17394, n17395, n17396, n17397, n17398, n17399, n17400, n17401,
         n17402, n17403, n17404, n17405, n17406, n17407, n17408, n17409,
         n17410, n17411, n17412, n17413, n17414, n17415, n17416, n17417,
         n17418, n17419, n17420, n17421, n17422, n17423, n17424, n17425,
         n17426, n17427, n17428, n17429, n17430, n17431, n17432, n17433,
         n17434, n17435, n17436, n17437, n17438, n17439, n17440, n17441,
         n17442, n17443, n17444, n17445, n17446, n17447, n17448, n17449,
         n17450, n17451, n17452, n17453, n17454, n17455, n17456, n17457,
         n17458, n17459, n17460, n17461, n17462, n17463, n17464, n17465,
         n17466, n17467, n17468, n17469, n17470, n17471, n17472, n17473,
         n17474, n17475, n17476, n17477, n17478, n17479, n17480, n17481,
         n17482, n17483, n17484, n17485, n17486, n17487, n17488, n17489,
         n17490, n17491, n17492, n17493, n17494, n17495, n17496, n17497,
         n17498, n17499, n17500, n17501, n17502, n17503, n17504, n17505,
         n17506, n17507, n17508, n17509, n17510, n17511, n17512, n17513,
         n17514, n17515, n17516, n17517, n17518, n17519, n17520, n17521,
         n17522, n17523, n17524, n17525, n17526, n17527, n17528, n17529,
         n17530, n17531, n17532, n17533, n17534, n17535, n17536, n17537,
         n17538, n17539, n17540, n17541, n17542, n17543, n17544, n17545,
         n17546, n17547, n17548, n17549, n17550, n17551, n17552, n17553,
         n17554, n17555, n17556, n17557, n17558, n17559, n17560, n17561,
         n17562, n17563, n17564, n17565, n17566, n17567, n17568, n17569,
         n17570, n17571, n17572, n17573, n17574, n17575, n17576, n17577,
         n17578, n17579, n17580, n17581, n17582, n17583, n17584, n17585,
         n17586, n17587, n17588, n17589, n17590, n17591, n17592, n17593,
         n17594, n17595, n17596, n17597, n17598, n17599, n17600, n17601,
         n17602, n17603, n17604, n17605, n17606, n17607, n17608, n17609,
         n17610, n17611, n17612, n17613, n17614, n17615, n17616, n17617,
         n17618, n17619, n17620, n17621, n17622, n17623, n17624, n17625,
         n17626, n17627, n17628, n17629, n17630, n17631, n17632, n17633,
         n17634, n17635, n17636, n17637, n17638, n17639, n17640, n17641,
         n17642, n17643, n17644, n17645, n17646, n17647, n17648, n17649,
         n17650, n17651, n17652, n17653, n17654, n17655, n17656, n17657,
         n17658, n17659, n17660, n17661, n17662, n17663, n17664, n17665,
         n17666, n17667, n17668, n17669, n17670, n17671, n17672, n17673,
         n17674, n17675, n17676, n17677, n17678, n17679, n17680, n17681,
         n17682, n17683, n17684, n17685, n17686, n17687, n17688, n17689,
         n17690, n17691, n17692, n17693, n17694, n17695, n17696, n17697,
         n17698, n17699, n17700, n17701, n17702, n17703, n17704, n17705,
         n17706, n17707, n17708, n17709, n17710, n17711, n17712, n17713,
         n17714, n17715, n17716, n17717, n17718, n17719, n17720, n17721,
         n17722, n17723, n17724, n17725, n17726, n17727, n17728, n17729,
         n17730, n17731, n17732, n17733, n17734, n17735, n17736, n17737,
         n17738, n17739, n17740, n17741, n17742, n17743, n17744, n17745,
         n17746, n17747, n17748, n17749, n17750, n17751, n17752, n17753,
         n17754, n17755, n17756, n17757, n17758, n17759, n17760, n17761,
         n17762, n17763, n17764, n17765, n17766, n17767, n17768, n17769,
         n17770, n17771, n17772, n17773, n17774, n17775, n17776, n17777,
         n17778, n17779, n17780, n17781, n17782, n17783, n17784, n17785,
         n17786, n17787, n17788, n17789, n17790, n17791, n17792, n17793,
         n17794, n17795, n17796, n17797, n17798, n17799, n17800, n17801,
         n17802, n17803, n17804, n17805, n17806, n17807, n17808, n17809,
         n17810, n17811, n17812, n17813, n17814, n17815, n17816, n17817,
         n17818, n17819, n17820, n17821, n17822, n17823, n17824, n17825,
         n17826, n17827, n17828, n17829, n17830, n17831, n17832, n17833,
         n17834, n17835, n17836, n17837, n17838, n17839, n17840, n17841,
         n17842, n17843, n17844, n17845, n17846, n17847, n17848, n17849,
         n17850, n17851, n17852, n17853, n17854, n17855, n17856, n17857,
         n17858, n17859, n17860, n17861, n17862, n17863, n17864, n17865,
         n17866, n17867, n17868, n17869, n17870, n17871, n17872, n17873,
         n17874, n17875, n17876, n17877, n17878, n17879, n17880, n17881,
         n17882, n17883, n17884, n17885, n17886, n17887, n17888, n17889,
         n17890, n17891, n17892, n17893, n17894, n17895, n17896, n17897,
         n17898, n17899, n17900, n17901, n17902, n17903, n17904, n17905,
         n17906, n17907, n17908, n17909, n17910, n17911, n17912, n17913,
         n17914, n17915, n17916, n17917, n17918, n17919, n17920, n17921,
         n17922, n17923, n17924, n17925, n17926, n17927, n17928, n17929,
         n17930, n17931, n17932, n17933, n17934, n17935, n17936, n17937,
         n17938, n17939, n17940, n17941, n17942, n17943, n17944, n17945,
         n17946, n17947, n17948, n17949, n17950, n17951, n17952, n17953,
         n17954, n17955, n17956, n17957, n17958, n17959, n17960, n17961,
         n17962, n17963, n17964, n17965, n17966, n17967, n17968, n17969,
         n17970, n17971, n17972, n17973, n17974, n17975, n17976, n17977,
         n17978, n17979, n17980, n17981, n17982, n17983, n17984, n17985,
         n17986, n17987, n17988, n17989, n17990, n17991, n17992, n17993,
         n17994, n17995, n17996, n17997, n17998, n17999, n18000, n18001,
         n18002, n18003, n18004, n18005, n18006, n18007, n18008, n18009,
         n18010, n18011, n18012, n18013, n18014, n18015, n18016, n18017,
         n18018, n18019, n18020, n18021, n18022, n18023, n18024, n18025,
         n18026, n18027, n18028, n18029, n18030, n18031, n18032, n18033,
         n18034, n18035, n18036, n18037, n18038, n18039, n18040, n18041,
         n18042, n18043, n18044, n18045, n18046, n18047, n18048, n18049,
         n18050, n18051, n18052, n18053, n18054, n18055, n18056, n18057,
         n18058, n18059, n18060, n18061, n18062, n18063, n18064, n18065,
         n18066, n18067, n18068, n18069, n18070, n18071, n18072, n18073,
         n18074, n18075, n18076, n18077, n18078, n18079, n18080, n18081,
         n18082, n18083, n18084, n18085, n18086, n18087, n18088, n18089,
         n18090, n18091, n18092, n18093, n18094, n18095, n18096, n18097,
         n18098, n18099, n18100, n18101, n18102, n18103, n18104, n18105,
         n18106, n18107, n18108, n18109, n18110, n18111, n18112, n18113,
         n18114, n18115, n18116, n18117, n18118, n18119, n18120, n18121,
         n18122, n18123, n18124, n18125, n18126, n18127, n18128, n18129,
         n18130, n18131, n18132, n18133, n18134, n18135, n18136, n18137,
         n18138, n18139, n18140, n18141, n18142, n18143, n18144, n18145,
         n18146, n18147, n18148, n18149, n18150, n18151, n18152, n18153,
         n18154, n18155, n18156, n18157, n18158, n18159, n18160, n18161,
         n18162, n18163, n18164, n18165, n18166, n18167, n18168, n18169,
         n18170, n18171, n18172, n18173, n18174, n18175, n18176, n18177,
         n18178, n18179, n18180, n18181, n18182, n18183, n18184, n18185,
         n18186, n18187, n18188, n18189, n18190, n18191, n18192, n18193,
         n18194, n18195, n18196, n18197, n18198, n18199, n18200, n18201,
         n18202, n18203, n18204, n18205, n18206, n18207, n18208, n18209,
         n18210, n18211, n18212, n18213, n18214, n18215, n18216, n18217,
         n18218, n18219, n18220, n18221, n18222, n18223, n18224, n18225,
         n18226, n18227, n18228, n18229, n18230, n18231, n18232, n18233,
         n18234, n18235, n18236, n18237, n18238, n18239, n18240, n18241,
         n18242, n18243, n18244, n18245, n18246, n18247, n18248, n18249,
         n18250, n18251, n18252, n18253, n18254, n18255, n18256, n18257,
         n18258, n18259, n18260, n18261, n18262, n18263, n18264, n18265,
         n18266, n18267, n18268, n18269, n18270, n18271, n18272, n18273,
         n18274, n18275, n18276, n18277, n18278, n18279, n18280, n18281,
         n18282, n18283, n18284, n18285, n18286, n18287, n18288, n18289,
         n18290, n18291, n18292, n18293, n18294, n18295, n18296, n18297,
         n18298, n18299, n18300, n18301, n18302, n18303, n18304, n18305,
         n18306, n18307, n18308, n18309, n18310, n18311, n18312, n18313,
         n18314, n18315, n18316, n18317, n18318, n18319, n18320, n18321,
         n18322, n18323, n18324, n18325, n18326, n18327, n18328, n18329,
         n18330, n18331, n18332, n18333, n18334, n18335, n18336, n18337,
         n18338, n18339, n18340, n18341, n18342, n18343, n18344, n18345,
         n18346, n18347, n18348, n18349, n18350, n18351, n18352, n18353,
         n18354, n18355, n18356, n18357, n18358, n18359, n18360, n18361,
         n18362, n18363, n18364, n18365, n18366, n18367, n18368, n18369,
         n18370, n18371, n18372, n18373, n18374, n18375, n18376, n18377,
         n18378, n18379, n18380, n18381, n18382, n18383, n18384, n18385,
         n18386, n18387, n18388, n18389, n18390, n18391, n18392, n18393,
         n18394, n18395, n18396, n18397, n18398, n18399, n18400, n18401,
         n18402, n18403, n18404, n18405, n18406, n18407, n18408, n18409,
         n18410, n18411, n18412, n18413, n18414, n18415, n18416, n18417,
         n18418, n18419, n18420, n18421, n18422, n18423, n18424, n18425,
         n18426, n18427, n18428, n18429, n18430, n18431, n18432, n18433,
         n18434, n18435, n18436, n18437, n18438, n18439, n18440, n18441,
         n18442, n18443, n18444, n18445, n18446, n18447, n18448, n18449,
         n18450, n18451, n18452, n18453, n18454, n18455, n18456, n18457,
         n18458, n18459, n18460, n18461, n18462, n18463, n18464, n18465,
         n18466, n18467, n18468, n18469, n18470, n18471, n18472, n18473,
         n18474, n18475, n18476, n18477, n18478, n18479, n18480, n18481,
         n18482, n18483, n18484, n18485, n18486, n18487, n18488, n18489,
         n18490, n18491, n18492, n18493, n18494, n18495, n18496, n18497,
         n18498, n18499, n18500, n18501, n18502, n18503, n18504, n18505,
         n18506, n18507, n18508, n18509, n18510, n18511, n18512, n18513,
         n18514, n18515, n18516, n18517, n18518, n18519, n18520, n18521,
         n18522, n18523, n18524, n18525, n18526, n18527, n18528, n18529,
         n18530, n18531, n18532, n18533, n18534, n18535, n18536, n18537,
         n18538, n18539, n18540, n18541, n18542, n18543, n18544, n18545,
         n18546, n18547, n18548, n18549, n18550, n18551, n18552, n18553,
         n18554, n18555, n18556, n18557, n18558, n18559, n18560, n18561,
         n18562, n18563, n18564, n18565, n18566, n18567, n18568, n18569,
         n18570, n18571, n18572, n18573, n18574, n18575, n18576, n18577,
         n18578, n18579, n18580, n18581, n18582, n18583, n18584, n18585,
         n18586, n18587, n18588, n18589, n18590, n18591, n18592, n18593,
         n18594, n18595, n18596, n18597, n18598, n18599, n18600, n18601,
         n18602, n18603, n18604, n18605, n18606, n18607, n18608, n18609,
         n18610, n18611, n18612, n18613, n18614, n18615, n18616, n18617,
         n18618, n18619, n18620, n18621, n18622, n18623, n18624, n18625,
         n18626, n18627, n18628, n18629, n18630, n18631, n18632, n18633,
         n18634, n18635, n18636, n18637, n18638, n18639, n18640, n18641,
         n18642, n18643, n18644, n18645, n18646, n18647, n18648, n18649,
         n18650, n18651, n18652, n18653, n18654, n18655, n18656, n18657,
         n18658, n18659, n18660, n18661, n18662, n18663, n18664, n18665,
         n18666, n18667, n18668, n18669, n18670, n18671, n18672, n18673,
         n18674, n18675, n18676, n18677, n18678, n18679, n18680, n18681,
         n18682, n18683, n18684, n18685, n18686, n18687, n18688, n18689,
         n18690, n18691, n18692, n18693, n18694, n18695, n18696, n18697,
         n18698, n18699, n18700, n18701, n18702, n18703, n18704, n18705,
         n18706, n18707, n18708, n18709, n18710, n18711, n18712, n18713,
         n18714, n18715, n18716, n18717, n18718, n18719, n18720, n18721,
         n18722, n18723, n18724, n18725, n18726, n18727, n18728, n18729,
         n18730, n18731, n18732, n18733, n18734, n18735, n18736, n18737,
         n18738, n18739, n18740, n18741, n18742, n18743, n18744, n18745,
         n18746, n18747, n18748, n18749, n18750, n18751, n18752, n18753,
         n18754, n18755, n18756, n18757, n18758, n18759, n18760, n18761,
         n18762, n18763, n18764, n18765, n18766, n18767, n18768, n18769,
         n18770, n18771, n18772, n18773, n18774, n18775, n18776, n18777,
         n18778, n18779, n18780, n18781, n18782, n18783, n18784, n18785,
         n18786, n18787, n18788, n18789, n18790, n18791, n18792, n18793,
         n18794, n18795, n18796, n18797, n18798, n18799, n18800, n18801,
         n18802, n18803, n18804, n18805, n18806, n18807, n18808, n18809,
         n18810, n18811, n18812, n18813, n18814, n18815, n18816, n18817,
         n18818, n18819, n18820, n18821, n18822, n18823, n18824, n18825,
         n18826, n18827, n18828, n18829, n18830, n18831, n18832, n18833,
         n18834, n18835, n18836, n18837, n18838, n18839, n18840, n18841,
         n18842, n18843, n18844, n18845, n18846, n18847, n18848, n18849,
         n18850, n18851, n18852, n18853, n18854, n18855, n18856, n18857,
         n18858, n18859, n18860, n18861, n18862, n18863, n18864, n18865,
         n18866, n18867, n18868, n18869, n18870, n18871, n18872, n18873,
         n18874, n18875, n18876, n18877, n18878, n18879, n18880, n18881,
         n18882, n18883, n18884, n18885, n18886, n18887, n18888, n18889,
         n18890, n18891, n18892, n18893, n18894, n18895, n18896, n18897,
         n18898, n18899, n18900, n18901, n18902, n18903, n18904, n18905,
         n18906, n18907, n18908, n18909, n18910, n18911, n18912, n18913,
         n18914, n18915, n18916, n18917, n18918, n18919, n18920, n18921,
         n18922, n18923, n18924, n18925, n18926, n18927, n18928, n18929,
         n18930, n18931, n18932, n18933, n18934, n18935, n18936, n18937,
         n18938, n18939, n18940, n18941, n18942, n18943, n18944, n18945,
         n18946, n18947, n18948, n18949, n18950, n18951, n18952, n18953,
         n18954, n18955, n18956, n18957, n18958, n18959, n18960, n18961,
         n18962, n18963, n18964, n18965, n18966, n18967, n18968, n18969,
         n18970, n18971, n18972, n18973, n18974, n18975, n18976, n18977,
         n18978, n18979, n18980, n18981, n18982, n18983, n18984, n18985,
         n18986, n18987, n18988, n18989, n18990, n18991, n18992, n18993,
         n18994, n18995, n18996, n18997, n18998, n18999, n19000, n19001,
         n19002, n19003, n19004, n19005, n19006, n19007, n19008, n19009,
         n19010, n19011, n19012, n19013, n19014, n19015, n19016, n19017,
         n19018, n19019, n19020, n19021, n19022, n19023, n19024, n19025,
         n19026, n19027, n19028, n19029, n19030, n19031, n19032, n19033,
         n19034, n19035, n19036, n19037, n19038, n19039, n19040, n19041,
         n19042, n19043, n19044, n19045, n19046, n19047, n19048, n19049,
         n19050, n19051, n19052, n19053, n19054, n19055, n19056, n19057,
         n19058, n19059, n19060, n19061, n19062, n19063, n19064, n19065,
         n19066, n19067, n19068, n19069, n19070, n19071, n19072, n19073,
         n19074, n19075, n19076, n19077, n19078, n19079, n19080, n19081,
         n19082, n19083, n19084, n19085, n19086, n19087, n19088, n19089,
         n19090, n19091, n19092, n19093, n19094, n19095, n19096, n19097,
         n19098, n19099, n19100, n19101, n19102, n19103, n19104, n19105,
         n19106, n19107, n19108, n19109, n19110, n19111, n19112, n19113,
         n19114, n19115, n19116, n19117, n19118, n19119, n19120, n19121,
         n19122, n19123, n19124, n19125, n19126, n19127, n19128, n19129,
         n19130, n19131, n19132, n19133, n19134, n19135, n19136, n19137,
         n19138, n19139, n19140, n19141, n19142, n19143, n19144, n19145,
         n19146, n19147, n19148, n19149, n19150, n19151, n19152, n19153,
         n19154, n19155, n19156, n19157, n19158, n19159, n19160, n19161,
         n19162, n19163, n19164, n19165, n19166, n19167, n19168, n19169,
         n19170, n19171, n19172, n19173, n19174, n19175, n19176, n19177,
         n19178, n19179, n19180, n19181, n19182, n19183, n19184, n19185,
         n19186, n19187, n19188, n19189, n19190, n19191, n19192, n19193,
         n19194, n19195, n19196, n19197, n19198, n19199, n19200, n19201,
         n19202, n19203, n19204, n19205, n19206, n19207, n19208, n19209,
         n19210, n19211, n19212, n19213, n19214, n19215, n19216, n19217,
         n19218, n19219, n19220, n19221, n19222, n19223, n19224, n19225,
         n19226, n19227, n19228, n19229, n19230, n19231, n19232, n19233,
         n19234, n19235, n19236, n19237, n19238, n19239, n19240, n19241,
         n19242, n19243, n19244, n19245, n19246, n19247, n19248, n19249,
         n19250, n19251, n19252, n19253, n19254, n19255, n19256, n19257,
         n19258, n19259, n19260, n19261, n19262, n19263, n19264, n19265,
         n19266, n19267, n19268, n19269, n19270, n19271, n19272, n19273,
         n19274, n19275, n19276, n19277, n19278, n19279, n19280, n19281,
         n19282, n19283, n19284, n19285, n19286, n19287, n19288, n19289,
         n19290, n19291, n19292, n19293, n19294, n19295, n19296, n19297,
         n19298, n19299, n19300, n19301, n19302, n19303, n19304, n19305,
         n19306, n19307, n19308, n19309, n19310, n19311, n19312, n19313,
         n19314, n19315, n19316, n19317, n19318, n19319, n19320, n19321,
         n19322, n19323, n19324, n19325, n19326, n19327, n19328, n19329,
         n19330, n19331, n19332, n19333, n19334, n19335, n19336, n19337,
         n19338, n19339, n19340, n19341, n19342, n19343, n19344, n19345,
         n19346, n19347, n19348, n19349, n19350, n19351, n19352, n19353,
         n19354, n19355, n19356, n19357, n19358, n19359, n19360, n19361,
         n19362, n19363, n19364, n19365, n19366, n19367, n19368, n19369,
         n19370, n19371, n19372, n19373, n19374, n19375, n19376, n19377,
         n19378, n19379, n19380, n19381, n19382, n19383, n19384, n19385,
         n19386, n19387, n19388, n19389, n19390, n19391, n19392, n19393,
         n19394, n19395, n19396, n19397, n19398, n19399, n19400, n19401,
         n19402, n19403, n19404, n19405, n19406, n19407, n19408, n19409,
         n19410, n19411, n19412, n19413, n19414, n19415, n19416, n19417,
         n19418, n19419, n19420, n19421, n19422, n19423, n19424, n19425,
         n19426, n19427, n19428, n19429, n19430, n19431, n19432, n19433,
         n19434, n19435, n19436, n19437, n19438, n19439, n19440, n19441,
         n19442, n19443, n19444, n19445, n19446, n19447, n19448, n19449,
         n19450, n19451, n19452, n19453, n19454, n19455, n19456, n19457,
         n19458, n19459, n19460, n19461, n19462, n19463, n19464, n19465,
         n19466, n19467, n19468, n19469, n19470, n19471, n19472, n19473,
         n19474, n19475, n19476, n19477, n19478, n19479, n19480, n19481,
         n19482, n19483, n19484, n19485, n19486, n19487, n19488, n19489,
         n19490, n19491, n19492, n19493, n19494, n19495, n19496, n19497,
         n19498, n19499, n19500, n19501, n19502, n19503, n19504, n19505,
         n19506, n19507, n19508, n19509, n19510, n19511, n19512, n19513,
         n19514, n19515, n19516, n19517, n19518, n19519, n19520, n19521,
         n19522, n19523, n19524, n19525, n19526, n19527, n19528, n19529,
         n19530, n19531, n19532, n19533, n19534, n19535, n19536, n19537,
         n19538, n19539, n19540, n19541, n19542, n19543, n19544, n19545,
         n19546, n19547, n19548, n19549, n19550, n19551, n19552, n19553,
         n19554, n19555, n19556, n19557, n19558, n19559, n19560, n19561,
         n19562, n19563, n19564, n19565, n19566, n19567, n19568, n19569,
         n19570, n19571, n19572, n19573, n19574, n19575, n19576, n19577,
         n19578, n19579, n19580, n19581, n19582, n19583, n19584, n19585,
         n19586, n19587, n19588, n19589, n19590, n19591, n19592, n19593,
         n19594, n19595, n19596, n19597, n19598, n19599, n19600, n19601,
         n19602, n19603, n19604, n19605, n19606, n19607, n19608, n19609,
         n19610, n19611, n19612, n19613, n19614, n19615, n19616, n19617,
         n19618, n19619, n19620, n19621, n19622, n19623, n19624, n19625,
         n19626, n19627, n19628, n19629, n19630, n19631, n19632, n19633,
         n19634, n19635, n19636, n19637, n19638, n19639, n19640, n19641,
         n19642, n19643, n19644, n19645, n19646, n19647, n19648, n19649,
         n19650, n19651, n19652, n19653, n19654, n19655, n19656, n19657,
         n19658, n19659, n19660, n19661, n19662, n19663, n19664, n19665,
         n19666, n19667, n19668, n19669, n19670, n19671, n19672, n19673,
         n19674, n19675, n19676, n19677, n19678, n19679, n19680, n19681,
         n19682, n19683, n19684, n19685, n19686, n19687, n19688, n19689,
         n19690, n19691, n19692, n19693, n19694, n19695, n19696, n19697,
         n19698, n19699, n19700, n19701, n19702, n19703, n19704, n19705,
         n19706, n19707, n19708, n19709, n19710, n19711, n19712, n19713,
         n19714, n19715, n19716, n19717, n19718, n19719, n19720, n19721,
         n19722, n19723, n19724, n19725, n19726, n19727, n19728, n19729,
         n19730, n19731, n19732, n19733, n19734, n19735, n19736, n19737,
         n19738, n19739, n19740, n19741, n19742, n19743, n19744, n19745,
         n19746, n19747, n19748, n19749, n19750, n19751, n19752, n19753,
         n19754, n19755, n19756, n19757, n19758, n19759, n19760, n19761,
         n19762, n19763, n19764, n19765, n19766, n19767, n19768, n19769,
         n19770, n19771, n19772, n19773, n19774, n19775, n19776, n19777,
         n19778, n19779, n19780, n19781, n19782, n19783, n19784, n19785,
         n19786, n19787, n19788, n19789, n19790, n19791, n19792, n19793,
         n19794, n19795, n19796, n19797, n19798, n19799, n19800, n19801,
         n19802, n19803, n19804, n19805, n19806, n19807, n19808, n19809,
         n19810, n19811, n19812, n19813, n19814, n19815, n19816, n19817,
         n19818, n19819, n19820, n19821, n19822, n19823, n19824, n19825,
         n19826, n19827, n19828, n19829, n19830, n19831, n19832, n19833,
         n19834, n19835, n19836, n19837, n19838, n19839, n19840, n19841,
         n19842, n19843, n19844, n19845, n19846, n19847, n19848, n19849,
         n19850, n19851, n19852, n19853, n19854, n19855, n19856, n19857,
         n19858, n19859, n19860, n19861, n19862, n19863, n19864, n19865,
         n19866, n19867, n19868, n19869, n19870, n19871, n19872, n19873,
         n19874, n19875, n19876, n19877, n19878, n19879, n19880, n19881,
         n19882, n19883, n19884, n19885, n19886, n19887, n19888, n19889,
         n19890, n19891, n19892, n19893, n19894, n19895, n19896, n19897,
         n19898, n19899, n19900, n19901, n19902, n19903, n19904, n19905,
         n19906, n19907, n19908, n19909, n19910, n19911, n19912, n19913,
         n19914, n19915, n19916, n19917, n19918, n19919, n19920, n19921,
         n19922, n19923, n19924, n19925, n19926, n19927, n19928, n19929,
         n19930, n19931, n19932, n19933, n19934, n19935, n19936, n19937,
         n19938, n19939, n19940, n19941, n19942, n19943, n19944, n19945,
         n19946, n19947, n19948, n19949, n19950, n19951, n19952, n19953,
         n19954, n19955, n19956, n19957, n19958, n19959, n19960, n19961,
         n19962, n19963, n19964, n19965, n19966, n19967, n19968, n19969,
         n19970, n19971, n19972, n19973, n19974, n19975, n19976, n19977,
         n19978, n19979, n19980, n19981, n19982, n19983, n19984, n19985,
         n19986, n19987, n19988, n19989, n19990, n19991, n19992, n19993,
         n19994, n19995, n19996, n19997, n19998, n19999, n20000, n20001,
         n20002, n20003, n20004, n20005, n20006, n20007, n20008, n20009,
         n20010, n20011, n20012, n20013, n20014, n20015, n20016, n20017,
         n20018, n20019, n20020, n20021, n20022, n20023, n20024, n20025,
         n20026, n20027, n20028, n20029, n20030, n20031, n20032, n20033,
         n20034, n20035, n20036, n20037, n20038, n20039, n20040, n20041,
         n20042, n20043, n20044, n20045, n20046, n20047, n20048, n20049,
         n20050, n20051, n20052, n20053, n20054, n20055, n20056, n20057,
         n20058, n20059, n20060, n20061, n20062, n20063, n20064, n20065,
         n20066, n20067, n20068, n20069, n20070, n20071, n20072, n20073,
         n20074, n20075, n20076, n20077, n20078, n20079, n20080, n20081,
         n20082, n20083, n20084, n20085, n20086, n20087, n20088, n20089,
         n20090, n20091, n20092, n20093, n20094, n20095, n20096, n20097,
         n20098, n20099, n20100, n20101, n20102, n20103, n20104, n20105,
         n20106, n20107, n20108, n20109, n20110, n20111, n20112, n20113,
         n20114, n20115, n20116, n20117, n20118, n20119, n20120, n20121,
         n20122, n20123, n20124, n20125, n20126, n20127, n20128, n20129,
         n20130, n20131, n20132, n20133, n20134, n20135, n20136, n20137,
         n20138, n20139, n20140, n20141, n20142, n20143, n20144, n20145,
         n20146, n20147, n20148, n20149, n20150, n20151, n20152, n20153,
         n20154, n20155, n20156, n20157, n20158, n20159, n20160, n20161,
         n20162, n20163, n20164, n20165, n20166, n20167, n20168, n20169,
         n20170, n20171, n20172, n20173, n20174, n20175, n20176, n20177,
         n20178, n20179, n20180, n20181, n20182, n20183, n20184, n20185,
         n20186, n20187, n20188, n20189, n20190, n20191, n20192, n20193,
         n20194, n20195, n20196, n20197, n20198, n20199, n20200, n20201,
         n20202, n20203, n20204, n20205, n20206, n20207, n20208, n20209,
         n20210, n20211, n20212, n20213, n20214, n20215, n20216, n20217,
         n20218, n20219, n20220, n20221, n20222, n20223, n20224, n20225,
         n20226, n20227, n20228, n20229, n20230, n20231, n20232, n20233,
         n20234, n20235, n20236, n20237, n20238, n20239, n20240, n20241,
         n20242, n20243, n20244, n20245, n20246, n20247, n20248, n20249,
         n20250, n20251, n20252, n20253, n20254, n20255, n20256, n20257,
         n20258, n20259, n20260, n20261, n20262, n20263, n20264, n20265,
         n20266, n20267, n20268, n20269, n20270, n20271, n20272, n20273,
         n20274, n20275, n20276, n20277, n20278, n20279, n20280, n20281,
         n20282, n20283, n20284, n20285, n20286, n20287, n20288, n20289,
         n20290, n20291, n20292, n20293, n20294, n20295, n20296, n20297,
         n20298, n20299, n20300, n20301, n20302, n20303, n20304, n20305,
         n20306, n20307, n20308, n20309, n20310, n20311, n20312, n20313,
         n20314, n20315, n20316, n20317, n20318, n20319, n20320, n20321,
         n20322, n20323, n20324, n20325, n20326, n20327, n20328, n20329,
         n20330, n20331, n20332, n20333, n20334, n20335, n20336, n20337,
         n20338, n20339, n20340, n20341, n20342, n20343, n20344, n20345,
         n20346, n20347, n20348, n20349, n20350, n20351, n20352, n20353,
         n20354, n20355, n20356, n20357, n20358, n20359, n20360, n20361,
         n20362, n20363, n20364, n20365, n20366, n20367, n20368, n20369,
         n20370, n20371, n20372, n20373, n20374, n20375, n20376, n20377,
         n20378, n20379, n20380, n20381, n20382, n20383, n20384, n20385,
         n20386, n20387, n20388, n20389, n20390, n20391, n20392, n20393,
         n20394, n20395, n20396, n20397, n20398, n20399, n20400, n20401,
         n20402, n20403, n20404, n20405, n20406, n20407, n20408, n20409,
         n20410, n20411, n20412, n20413, n20414, n20415, n20416, n20417,
         n20418, n20419, n20420, n20421, n20422, n20423, n20424, n20425,
         n20426, n20427, n20428, n20429, n20430, n20431, n20432, n20433,
         n20434, n20435, n20436, n20437, n20438, n20439, n20440, n20441,
         n20442, n20443, n20444, n20445, n20446, n20447, n20448, n20449,
         n20450, n20451, n20452, n20453, n20454, n20455, n20456, n20457,
         n20458, n20459, n20460, n20461, n20462, n20463, n20464, n20465,
         n20466, n20467, n20468, n20469, n20470, n20471, n20472, n20473,
         n20474, n20475, n20476, n20477, n20478, n20479, n20480, n20481,
         n20482, n20483, n20484, n20485, n20486, n20487, n20488, n20489,
         n20490, n20491, n20492, n20493, n20494, n20495, n20496, n20497,
         n20498, n20499, n20500, n20501, n20502, n20503, n20504, n20505,
         n20506, n20507, n20508, n20509, n20510, n20511, n20512, n20513,
         n20514, n20515, n20516, n20517, n20518, n20519, n20520, n20521,
         n20522, n20523, n20524, n20525, n20526, n20527, n20528, n20529,
         n20530, n20531, n20532, n20533, n20534, n20535, n20536, n20537,
         n20538, n20539, n20540, n20541, n20542, n20543, n20544, n20545,
         n20546, n20547, n20548, n20549, n20550, n20551, n20552, n20553,
         n20554, n20555, n20556, n20557, n20558, n20559, n20560, n20561,
         n20562, n20563, n20564, n20565, n20566, n20567, n20568, n20569,
         n20570, n20571, n20572, n20573, n20574, n20575, n20576, n20577,
         n20578, n20579, n20580, n20581, n20582, n20583, n20584, n20585,
         n20586, n20587, n20588, n20589, n20590, n20591, n20592, n20593,
         n20594, n20595, n20596, n20597, n20598, n20599, n20600, n20601,
         n20602, n20603, n20604, n20605, n20606, n20607, n20608, n20609,
         n20610, n20611, n20612, n20613, n20614, n20615, n20616, n20617,
         n20618, n20619, n20620, n20621, n20622, n20623, n20624, n1, n2, n3,
         n4, n5, n6, n7, n8, n9, n10, n11, n12, n24, n27, n30, n33, n36, n39,
         n168, n171, n174, n177, n180, n183, n186, n189, n192, n195, n198,
         n201, n204, n207, n210, n213, n218, n348, n478, n608, n738, n868,
         n998, n1128, n1258, n1387, n1516, n1645, n1774, n1903, n2032, n2161,
         n2291, n2420, n2549, n2678, n2807, n2936, n3065, n3194, n3324, n3453,
         n3582, n3711, n3840, n3969, n4098, n20625, n20626, n20627, n20628,
         n20629, n20630, n20631, n20632, n20633, n20634, n20635, n20636,
         n20637, n20638, n20639, n20640, n20641, n20642, n20643, n20644,
         n20645, n20646, n20647, n20648, n20649, n20650, n20651, n20652,
         n20653, n20654, n20655, n20656, n20657, n20658, n20659, n20660,
         n20661, n20662, n20663, n20664, n20665, n20666, n20667, n20668,
         n20669, n20670, n20671, n20672, n20673, n20674, n20675, n20676,
         n20677, n20678, n20679, n20680, n20681, n20682, n20683, n20684,
         n20685, n20686, n20687, n20688, n20689, n20690, n20691, n20692,
         n20693, n20694, n20695, n20696, n20697, n20698, n20699, n20700,
         n20701, n20702, n20703, n20704, n20705, n20706, n20707, n20708,
         n20709, n20710, n20711, n20712, n20713, n20714, n20715, n20716,
         n20717, n20718, n20719, n20720, n20721, n20722, n20723, n20724,
         n20725, n20726, n20727, n20728, n20729, n20730, n20731, n20732,
         n20733, n20734, n20735, n20736, n20737, n20738, n20739, n20740,
         n20741, n20742, n20743, n20744, n20745, n20746, n20747, n20748,
         n20749, n20750, n20751, n20752, n20753, n20754, n20755, n20756,
         n20757, n20758, n20759, n20760, n20761, n20762, n20763, n20764,
         n20765, n20766, n20767, n20768, n20769, n20770, n20771, n20772,
         n20773, n20774, n20775, n20776, n20777, n20778, n20779, n20780,
         n20781, n20782, n20783, n20784, n20785, n20786, n20787, n20788,
         n20789, n20790, n20791, n20792, n20793, n20794, n20795, n20796,
         n20797, n20798, n20799, n20800, n20801, n20802, n20803, n20804,
         n20805, n20806, n20807, n20808, n20809, n20810, n20811, n20812,
         n20813, n20814, n20815, n20816, n20817, n20818, n20819, n20820,
         n20821, n20822, n20823, n20824, n20825, n20826, n20827, n20828,
         n20829, n20830, n20831, n20832, n20833, n20834, n20835, n20836,
         n20837, n20838, n20839, n20840, n20841, n20842, n20843, n20844,
         n20845, n20846, n20847, n20848, n20849, n20850, n20851, n20852,
         n20853, n20854, n20855, n20856, n20857, n20858, n20859, n20860,
         n20861, n20862, n20863, n20864, n20865, n20866, n20867, n20868,
         n20869, n20870, n20871, n20872, n20873, n20874, n20875, n20876,
         n20877, n20878, n20879, n20880, n20881, n20882, n20883, n20884,
         n20885, n20886, n20887, n20888, n20889, n20890, n20891, n20892,
         n20893, n20894, n20895, n20896, n20897, n20898, n20899, n20900,
         n20901, n20902, n20903, n20904, n20905, n20906, n20907, n20908,
         n20909, n20910, n20911, n20912, n20913, n20914, n20915, n20916,
         n20917, n20918, n20919, n20920, n20921, n20922, n20923, n20924,
         n20925, n20926, n20927, n20928, n20929, n20930, n20931, n20932,
         n20933, n20934, n20935, n20936, n20937, n20938, n20939, n20940,
         n20941, n20942, n20943, n20944, n20945, n20946, n20947, n20948,
         n20949, n20950, n20951, n20952, n20953, n20954, n20955, n20956,
         n20957, n20958, n20959, n20960, n20961, n20962, n20963, n20964,
         n20965, n20966, n20967, n20968, n20969, n20970, n20971, n20972,
         n20973, n20974, n20975, n20976, n20977, n20978, n20979, n20980,
         n20981, n20982, n20983, n20984, n20985, n20986, n20987, n20988,
         n20989, n20990, n20991, n20992, n20993, n20994, n20995, n20996,
         n20997, n20998, n20999, n21000, n21001, n21002, n21003, n21004,
         n21005, n21006, n21007, n21008, n21009, n21010, n21011, n21012,
         n21013, n21014, n21015, n21016, n21017, n21018, n21019, n21020,
         n21021, n21022, n21023, n21024, n21025, n21026, n21027, n21028,
         n21029, n21030, n21031, n21032, n21033, n21034, n21035, n21036,
         n21037, n21038, n21039, n21040, n21041, n21042, n21043, n21044,
         n21045, n21046, n21047, n21048, n21049, n21050, n21051, n21052,
         n21053, n21054, n21055, n21056, n21057, n21058, n21059, n21060,
         n21061, n21062, n21063, n21064, n21065, n21066, n21067, n21068,
         n21069, n21070, n21071, n21072, n21073, n21074, n21075, n21076,
         n21077, n21078, n21079, n21080, n21081, n21082, n21083, n21084,
         n21085, n21086, n21087, n21088, n21089, n21090, n21091, n21092,
         n21093, n21094, n21095, n21096, n21097, n21098, n21099, n21100,
         n21101, n21102, n21103, n21104, n21105, n21106, n21107, n21108,
         n21109, n21110, n21111, n21112, n21113, n21114, n21115, n21116,
         n21117, n21118, n21119, n21120, n21121, n21122, n21123, n21124,
         n21125, n21126, n21127, n21128, n21129, n21130, n21131, n21132,
         n21133, n21134, n21135, n21136, n21137, n21138, n21139, n21140,
         n21141, n21142, n21143, n21144, n21145, n21146, n21147, n21148,
         n21149, n21150, n21151, n21152, n21153, n21154, n21155, n21156,
         n21157, n21158, n21159, n21160, n21161, n21162, n21163, n21164,
         n21165, n21166, n21167, n21168, n21169, n21170, n21171, n21172,
         n21173, n21174, n21175, n21176, n21177, n21178, n21179, n21180,
         n21181, n21182, n21183, n21184, n21185, n21186, n21187, n21188,
         n21189, n21190, n21191, n21192, n21193, n21194, n21195, n21196,
         n21197, n21198, n21199, n21200, n21201, n21202, n21203, n21204,
         n21205, n21206, n21207, n21208, n21209, n21210, n21211, n21212,
         n21213, n21214, n21215, n21216, n21217, n21218, n21219, n21220,
         n21221, n21222, n21223, n21224, n21225, n21226, n21227, n21228,
         n21229, n21230, n21231, n21232, n21233, n21234, n21235, n21236,
         n21237, n21238, n21239, n21240, n21241, n21242, n21243, n21244,
         n21245, n21246, n21247, n21248, n21249, n21250, n21251, n21252,
         n21253, n21254, n21255, n21256, n21257, n21258, n21259, n21260,
         n21261, n21262, n21263, n21264, n21265, n21266, n21267, n21268,
         n21269, n21270, n21271, n21272, n21273, n21274, n21275, n21276,
         n21277, n21278, n21279, n21280, n21281, n21282, n21283, n21284,
         n21285, n21286, n21287, n21288, n21289, n21290, n21291, n21292,
         n21293, n21294, n21295, n21296, n21297, n21298, n21299, n21300,
         n21301, n21302, n21303, n21304, n21305, n21306, n21307, n21308,
         n21309, n21310, n21311, n21312, n21313, n21314, n21315, n21316,
         n21317, n21318, n21319, n21320, n21321, n21322, n21323, n21324,
         n21325, n21326, n21327, n21328, n21329, n21330, n21331, n21332,
         n21333, n21334, n21335, n21336, n21337, n21338, n21339, n21340,
         n21341, n21342, n21343, n21344, n21345, n21346, n21347, n21348,
         n21349, n21350, n21351, n21352, n21353, n21354, n21355, n21356,
         n21357, n21358, n21359, n21360, n21361, n21362, n21363, n21364,
         n21365, n21366, n21367, n21368, n21369, n21370, n21371, n21372,
         n21373, n21374, n21375, n21376, n21377, n21378, n21379, n21380,
         n21381, n21382, n21383, n21384, n21385, n21386, n21387, n21388,
         n21389, n21390, n21391, n21392, n21393, n21394, n21395, n21396,
         n21397, n21398, n21399, n21400, n21401, n21402, n21403, n21404,
         n21405, n21406, n21407, n21408, n21409, n21410, n21411, n21412,
         n21413, n21414, n21415, n21416, n21417, n21418, n21419, n21420,
         n21421, n21422, n21423, n21424, n21425, n21426, n21427, n21428,
         n21429, n21430, n21431, n21432, n21433, n21434, n21435, n21436,
         n21437, n21438, n21439, n21440, n21441, n21442, n21443, n21444,
         n21445, n21446, n21447, n21448, n21449, n21450, n21451, n21452,
         n21453, n21454, n21455, n21456, n21457, n21458, n21459, n21460,
         n21461, n21462, n21463, n21464, n21465, n21466, n21467, n21468,
         n21469, n21470, n21471, n21472, n21473, n21474, n21475, n21476,
         n21477, n21478, n21479, n21480, n21481, n21482, n21483, n21484,
         n21485, n21486, n21487, n21488, n21489, n21490, n21491, n21492,
         n21493, n21494, n21495, n21496, n21497, n21498, n21499, n21500,
         n21501, n21502, n21503, n21504, n21505, n21506, n21507, n21508,
         n21509, n21510, n21511, n21512, n21513, n21514, n21515, n21516,
         n21517, n21518, n21519, n21520, n21521, n21522, n21523, n21524,
         n21525, n21526, n21527, n21528, n21529, n21530, n21531, n21532,
         n21533, n21534, n21535, n21536, n21537, n21538, n21539, n21540,
         n21541, n21542, n21543, n21544, n21545, n21546, n21547, n21548,
         n21549, n21550, n21551, n21552, n21553, n21554, n21555, n21556,
         n21557, n21558, n21559, n21560, n21561, n21562, n21563, n21564,
         n21565, n21566, n21567, n21568, n21569, n21570, n21571, n21572,
         n21573, n21574, n21575, n21576, n21577, n21578, n21579, n21580,
         n21581, n21582, n21583, n21584, n21585, n21586, n21587, n21588,
         n21589, n21590, n21591, n21592, n21593, n21594, n21595, n21596,
         n21597, n21598, n21599, n21600, n21601, n21602, n21603, n21604,
         n21605, n21606, n21607, n21608, n21609, n21610, n21611, n21612,
         n21613, n21614, n21615, n21616, n21617, n21618, n21619, n21620,
         n21621, n21622, n21623, n21624, n21625, n21626, n21627, n21628,
         n21629, n21630, n21631, n21632, n21633, n21634, n21635, n21636,
         n21637, n21638, n21639, n21640, n21641, n21642, n21643, n21644,
         n21645, n21646, n21647, n21648, n21649, n21650, n21651, n21652,
         n21653, n21654, n21655, n21656, n21657, n21658, n21659, n21660,
         n21661, n21662, n21663, n21664, n21665, n21666, n21667, n21668,
         n21669, n21670, n21671, n21672, n21673, n21674, n21675, n21676,
         n21677, n21678, n21679, n21680, n21681, n21682, n21683, n21684,
         n21685, n21686, n21687, n21688, n21689, n21690, n21691, n21692,
         n21693, n21694, n21695, n21696, n21697, n21698, n21699, n21700,
         n21701, n21702, n21703, n21704, n21705, n21706, n21707, n21708,
         n21709, n21710, n21711, n21712, n21713, n21714, n21715, n21716,
         n21717, n21718, n21719, n21720, n21721, n21722, n21723, n21724,
         n21725, n21726, n21727, n21728, n21729, n21730, n21731, n21732,
         n21733, n21734, n21735, n21736, n21737, n21738, n21739, n21740,
         n21741, n21742, n21743, n21744, n21745, n21746, n21747, n21748,
         n21749, n21750, n21751, n21752, n21753, n21754, n21755, n21756,
         n21757, n21758, n21759, n21760, n21761, n21762, n21763, n21764,
         n21765, n21766, n21767, n21768, n21769, n21770, n21771, n21772,
         n21773, n21774, n21775, n21776, n21777, n21778, n21779, n21780,
         n21781, n21782, n21783, n21784, n21785, n21786, n21787, n21788,
         n21789, n21790, n21791, n21792, n21793, n21794, n21795, n21796,
         n21797, n21798, n21799, n21800, n21801, n21802, n21803, n21804,
         n21805, n21806, n21807, n21808, n21809, n21810, n21811, n21812,
         n21813, n21814, n21815, n21816, n21817, n21818, n21819, n21820,
         n21821, n21822, n21823, n21824, n21825, n21826, n21827, n21828,
         n21829, n21830, n21831, n21832, n21833, n21834, n21835, n21836,
         n21837, n21838, n21839, n21840, n21841, n21842, n21843, n21844,
         n21845, n21846, n21847, n21848, n21849, n21850, n21851, n21852,
         n21853, n21854, n21855, n21856, n21857, n21858, n21859, n21860,
         n21861, n21862, n21863, n21864, n21865, n21866, n21867, n21868,
         n21869, n21870, n21871, n21872, n21873, n21874, n21875, n21876,
         n21877, n21878, n21879, n21880, n21881, n21882, n21883, n21884,
         n21885, n21886, n21887, n21888, n21889, n21890, n21891, n21892,
         n21893, n21894, n21895, n21896, n21897, n21898, n21899, n21900,
         n21901, n21902, n21903, n21904, n21905, n21906, n21907, n21908,
         n21909, n21910, n21911, n21912, n21913, n21914, n21915, n21916,
         n21917, n21918, n21919, n21920, n21921, n21922, n21923, n21924,
         n21925, n21926, n21927, n21928, n21929, n21930, n21931, n21932,
         n21933, n21934, n21935, n21936, n21937, n21938, n21939, n21940,
         n21941, n21942, n21943, n21944, n21945, n21946, n21947, n21948,
         n21949, n21950, n21951, n21952, n21953, n21954, n21955, n21956,
         n21957, n21958, n21959, n21960, n21961, n21962, n21963, n21964,
         n21965, n21966, n21967, n21968, n21969, n21970, n21971, n21972,
         n21973, n21974, n21975, n21976, n21977, n21978, n21979, n21980,
         n21981, n21982, n21983, n21984, n21985, n21986, n21987, n21988,
         n21989, n21990, n21991, n21992, n21993, n21994, n21995, n21996,
         n21997, n21998, n21999, n22000, n22001, n22002, n22003, n22004,
         n22005, n22006, n22007, n22008, n22009, n22010, n22011, n22012,
         n22013, n22014, n22015, n22016, n22017, n22018, n22019, n22020,
         n22021, n22022, n22023, n22024, n22025, n22026, n22027, n22028,
         n22029, n22030, n22031, n22032, n22033, n22034, n22035, n22036,
         n22037, n22038, n22039, n22040, n22041, n22042, n22043, n22044,
         n22045, n22046, n22047, n22048, n22049, n22050, n22051, n22052,
         n22053, n22054, n22055, n22056, n22057, n22058, n22059, n22060,
         n22061, n22062, n22063, n22064, n22065, n22066, n22067, n22068,
         n22069, n22070, n22071, n22072, n22073, n22074, n22075, n22076,
         n22077, n22078, n22079, n22080, n22081, n22082, n22083, n22084,
         n22085, n22086, n22087, n22088, n22089, n22090, n22091, n22092,
         n22093, n22094, n22095, n22096, n22097, n22098, n22099, n22100,
         n22101, n22102, n22103, n22104, n22105, n22106, n22107, n22108,
         n22109, n22110, n22111, n22112, n22113, n22114, n22115, n22116,
         n22117, n22118, n22119, n22120, n22121, n22122, n22123, n22124,
         n22125, n22126, n22127, n22128, n22129, n22130, n22131, n22132,
         n22133, n22134, n22135, n22136, n22137, n22138, n22139, n22140,
         n22141, n22142, n22143, n22144, n22145, n22146, n22147, n22148,
         n22149, n22150, n22151, n22152, n22153, n22154, n22155, n22156,
         n22157, n22158, n22159, n22160, n22161, n22162, n22163, n22164,
         n22165, n22166, n22167, n22168, n22169, n22170, n22171, n22172,
         n22173, n22174, n22175, n22176, n22177, n22178, n22179, n22180,
         n22181, n22182, n22183, n22184, n22185, n22186, n22187, n22188,
         n22189, n22190, n22191, n22192, n22193, n22194, n22195, n22196,
         n22197, n22198, n22199, n22200, n22201, n22202, n22203, n22204,
         n22205, n22206, n22207, n22208, n22209, n22210, n22211, n22212,
         n22213, n22214, n22215, n22216, n22217, n22218, n22219, n22220,
         n22221, n22222, n22223, n22224, n22225, n22226, n22227, n22228,
         n22229, n22230, n22231, n22232, n22233, n22234, n22235, n22236,
         n22237, n22238, n22239, n22240, n22241, n22242, n22243, n22244,
         n22245, n22246, n22247, n22248, n22249, n22250, n22251, n22252,
         n22253, n22254, n22255, n22256, n22257, n22258, n22259, n22260,
         n22261, n22262, n22263, n22264, n22265, n22266, n22267, n22268,
         n22269, n22270, n22271, n22272, n22273, n22274, n22275, n22276,
         n22277, n22278, n22279, n22280, n22281, n22282, n22283, n22284,
         n22285, n22286, n22287, n22288, n22289, n22290, n22291, n22292,
         n22293, n22294, n22295, n22296, n22297, n22298, n22299, n22300,
         n22301, n22302, n22303, n22304, n22305, n22306, n22307, n22308,
         n22309, n22310, n22311, n22312, n22313, n22314, n22315, n22316,
         n22317, n22318, n22319, n22320, n22321, n22322, n22323, n22324,
         n22325, n22326, n22327, n22328, n22329, n22330, n22331, n22332,
         n22333, n22334, n22335, n22336, n22337, n22338, n22339, n22340,
         n22341, n22342, n22343, n22344, n22345, n22346, n22347, n22348,
         n22349, n22350, n22351, n22352, n22353, n22354, n22355, n22356,
         n22357, n22358, n22359, n22360, n22361, n22362, n22363, n22364,
         n22365, n22366, n22367, n22368, n22369, n22370, n22371, n22372,
         n22373, n22374, n22375, n22376, n22377, n22378, n22379, n22380,
         n22381, n22382, n22383, n22384, n22385, n22386, n22387, n22388,
         n22389, n22390, n22391, n22392, n22393, n22394, n22395, n22396,
         n22397, n22398, n22399, n22400, n22401, n22402, n22403, n22404,
         n22405, n22406, n22407, n22408, n22409, n22410, n22411, n22412,
         n22413, n22414, n22415, n22416, n22417, n22418, n22419, n22420,
         n22421, n22422, n22423, n22424, n22425, n22426, n22427, n22428,
         n22429, n22430, n22431, n22432, n22433, n22434, n22435, n22436,
         n22437, n22438, n22439, n22440, n22441, n22442, n22443, n22444,
         n22445, n22446, n22447, n22448, n22449, n22450, n22451, n22452,
         n22453, n22454, n22455, n22456, n22457, n22458, n22459, n22460,
         n22461, n22462, n22463, n22464, n22465, n22466, n22467, n22468,
         n22469, n22470, n22471, n22472, n22473, n22474, n22475, n22476,
         n22477, n22478, n22479, n22480, n22481, n22482, n22483, n22484,
         n22485, n22486, n22487, n22488, n22489, n22490, n22491, n22492,
         n22493, n22494, n22495, n22496, n22497, n22498, n22499, n22500,
         n22501, n22502, n22503, n22504, n22505, n22506, n22507, n22508,
         n22509, n22510, n22511, n22512, n22513, n22514, n22515, n22516,
         n22517, n22518, n22519, n22520, n22521, n22522, n22523, n22524,
         n22525, n22526, n22527, n22528, n22529, n22530, n22531, n22532,
         n22533, n22534, n22535, n22536, n22537, n22538, n22539, n22540,
         n22541, n22542, n22543, n22544, n22545, n22546, n22547, n22548,
         n22549, n22550, n22551, n22552, n22553, n22554, n22555, n22556,
         n22557, n22558, n22559, n22560, n22561, n22562, n22563, n22564,
         n22565, n22566, n22567, n22568, n22569, n22570, n22571, n22572,
         n22573, n22574, n22575, n22576, n22577, n22578, n22579, n22580,
         n22581, n22582, n22583, n22584, n22585, n22586, n22587, n22588,
         n22589, n22590, n22591, n22592, n22593, n22594, n22595, n22596,
         n22597, n22598, n22599, n22600, n22601, n22602, n22603, n22604,
         n22605, n22606, n22607, n22608, n22609, n22610, n22611, n22612,
         n22613, n22614, n22615, n22616, n22617, n22618, n22619, n22620,
         n22621, n22622, n22623, n22624, n22625, n22626, n22627, n22628,
         n22629, n22630, n22631, n22632, n22633, n22634, n22635, n22636,
         n22637, n22638, n22639, n22640, n22641, n22642, n22643, n22644,
         n22645, n22646, n22647, n22648, n22649, n22650, n22651, n22652,
         n22653, n22654, n22655, n22656, n22657, n22658, n22659, n22660,
         n22661, n22662, n22663, n22664, n22665, n22666, n22667, n22668,
         n22669, n22670, n22671, n22672, n22673, n22674, n22675, n22676,
         n22677, n22678, n22679, n22680, n22681, n22682, n22683, n22684,
         n22685, n22686, n22687, n22688, n22689, n22690, n22691, n22692,
         n22693, n22694, n22695, n22696, n22697, n22698, n22699, n22700,
         n22701, n22702, n22703, n22704, n22705, n22706, n22707, n22708,
         n22709, n22710, n22711, n22712, n22713, n22714, n22715, n22716,
         n22717, n22718, n22719, n22720, n22721, n22722, n22723, n22724,
         n22725, n22726, n22727, n22728, n22729, n22730, n22731, n22732,
         n22733, n22734, n22735, n22736, n22737, n22738, n22739, n22740,
         n22741, n22742, n22743, n22744, n22745, n22746, n22747, n22748,
         n22749, n22750, n22751, n22752, n22753, n22754, n22755, n22756,
         n22757, n22758, n22759, n22760, n22761, n22762, n22763, n22764,
         n22765, n22766, n22767, n22768, n22769, n22770, n22771, n22772,
         n22773, n22774, n22775, n22776, n22777, n22778, n22779, n22780,
         n22781, n22782, n22783, n22784, n22785, n22786, n22787, n22788,
         n22789, n22790, n22791, n22792, n22793, n22794, n22795, n22796,
         n22797, n22798, n22799, n22800, n22801, n22802, n22803, n22804,
         n22805, n22806, n22807, n22808, n22809, n22810, n22811, n22812,
         n22813, n22814, n22815, n22816, n22817, n22818, n22819, n22820,
         n22821, n22822, n22823, n22824, n22825, n22826, n22827, n22828,
         n22829, n22830, n22831, n22832, n22833, n22834, n22835, n22836,
         n22837, n22838, n22839, n22840, n22841, n22842, n22843, n22844,
         n22845, n22846, n22847, n22848, n22849, n22850, n22851, n22852,
         n22853, n22854, n22855, n22856, n22857, n22858, n22859, n22860,
         n22861, n22862, n22863, n22864, n22865, n22866, n22867, n22868,
         n22869, n22870, n22871, n22872, n22873, n22874, n22875, n22876,
         n22877, n22878, n22879, n22880, n22881, n22882, n22883, n22884,
         n22885, n22886, n22887, n22888, n22889, n22890, n22891, n22892,
         n22893, n22894, n22895, n22896, n22897, n22898, n22899, n22900,
         n22901, n22902, n22903, n22904, n22905, n22906, n22907, n22908,
         n22909, n22910, n22911, n22912, n22913, n22914, n22915, n22916,
         n22917, n22918, n22919, n22920, n22921, n22922, n22923, n22924,
         n22925, n22926, n22927, n22928, n22929, n22930, n22931, n22932,
         n22933, n22934, n22935, n22936, n22937, n22938, n22939, n22940,
         n22941, n22942, n22943, n22944, n22945, n22946, n22947, n22948,
         n22949, n22950, n22951, n22952, n22953, n22954, n22955, n22956,
         n22957, n22958, n22959, n22960, n22961, n22962, n22963, n22964,
         n22965, n22966, n22967, n22968, n22969, n22970, n22971, n22972,
         n22973, n22974, n22975, n22976, n22977, n22978, n22979, n22980,
         n22981, n22982, n22983, n22984, n22985, n22986, n22987, n22988,
         n22989, n22990, n22991, n22992, n22993, n22994, n22995, n22996,
         n22997, n22998, n22999, n23000, n23001, n23002, n23003, n23004,
         n23005, n23006, n23007, n23008, n23009, n23010, n23011, n23012,
         n23013, n23014, n23015, n23016, n23017, n23018, n23019, n23020,
         n23021, n23022, n23023, n23024, n23025, n23026, n23027, n23028,
         n23029, n23030, n23031, n23032, n23033, n23034, n23035, n23036,
         n23037, n23038, n23039, n23040, n23041, n23042, n23043, n23044,
         n23045, n23046, n23047, n23048, n23049, n23050, n23051, n23052,
         n23053, n23054, n23055, n23056, n23057, n23058, n23059, n23060,
         n23061, n23062, n23063, n23064, n23065, n23066, n23067, n23068,
         n23069, n23070, n23071, n23072, n23073, n23074, n23075, n23076,
         n23077, n23078, n23079, n23080, n23081, n23082, n23083, n23084,
         n23085, n23086, n23087, n23088, n23089, n23090, n23091, n23092,
         n23093, n23094, n23095, n23096, n23097, n23098, n23099, n23100,
         n23101, n23102, n23103, n23104, n23105, n23106, n23107, n23108,
         n23109, n23110, n23111, n23112, n23113, n23114, n23115, n23116,
         n23117, n23118, n23119, n23120, n23121, n23122, n23123, n23124,
         n23125, n23126, n23127, n23128, n23129, n23130, n23131, n23132,
         n23133, n23134, n23135, n23136, n23137, n23138, n23139, n23140,
         n23141, n23142, n23143, n23144, n23145, n23146, n23147, n23148,
         n23149, n23150, n23151, n23152, n23153, n23154, n23155, n23156,
         n23157, n23158, n23159, n23160, n23161, n23162, n23163, n23164,
         n23165, n23166, n23167, n23168, n23169, n23170, n23171, n23172,
         n23173, n23174, n23175, n23176, n23177, n23178, n23179, n23180,
         n23181, n23182, n23183, n23184, n23185, n23186, n23187, n23188,
         n23189, n23190, n23191, n23192, n23193, n23194, n23195, n23196,
         n23197, n23198, n23199, n23200, n23201, n23202, n23203, n23204,
         n23205, n23206, n23207, n23208, n23209, n23210, n23211, n23212,
         n23213, n23214, n23215, n23216, n23217, n23218, n23219, n23220,
         n23221, n23222, n23223, n23224, n23225, n23226, n23227, n23228,
         n23229, n23230, n23231, n23232, n23233, n23234, n23235, n23236,
         n23237, n23238, n23239, n23240, n23241, n23242, n23243, n23244,
         n23245, n23246, n23247, n23248, n23249, n23250, n23251, n23252,
         n23253, n23254, n23255, n23256, n23257, n23258, n23259, n23260,
         n23261, n23262, n23263, n23264, n23265, n23266, n23267, n23268,
         n23269, n23270, n23271, n23272, n23273, n23274, n23275, n23276,
         n23277, n23278, n23279, n23280, n23281, n23282, n23283, n23284,
         n23285, n23286, n23287, n23288, n23289, n23290, n23291, n23292,
         n23293, n23294, n23295, n23296, n23297, n23298, n23299, n23300,
         n23301, n23302, n23303, n23304, n23305, n23306, n23307, n23308,
         n23309, n23310, n23311, n23312, n23313, n23314, n23315, n23316,
         n23317, n23318, n23319, n23320, n23321, n23322, n23323, n23324,
         n23325, n23326, n23327, n23328, n23329, n23330, n23331, n23332,
         n23333, n23334, n23335, n23336, n23337, n23338, n23339, n23340,
         n23341, n23342, n23343, n23344, n23345, n23346, n23347, n23348,
         n23349, n23350, n23351, n23352, n23353, n23354, n23355, n23356,
         n23357, n23358, n23359, n23360, n23361, n23362, n23363, n23364,
         n23365, n23366, n23367, n23368, n23369, n23370, n23371, n23372,
         n23373, n23374, n23375, n23376, n23377, n23378, n23379, n23380,
         n23381, n23382, n23383, n23384, n23385, n23386, n23387, n23388,
         n23389, n23390, n23391, n23392, n23393, n23394, n23395, n23396,
         n23397, n23398, n23399, n23400, n23401, n23402, n23403, n23404,
         n23405, n23406, n23407, n23408, n23409, n23410, n23411, n23412,
         n23413, n23414, n23415, n23416, n23417, n23418, n23419, n23420,
         n23421, n23422, n23423, n23424, n23425, n23426, n23427, n23428,
         n23429, n23430, n23431, n23432, n23433, n23434, n23435, n23436,
         n23437, n23438, n23439, n23440, n23441, n23442, n23443, n23444,
         n23445, n23446, n23447, n23448, n23449, n23450, n23451, n23452,
         n23453, n23454, n23455, n23456, n23457, n23458, n23459, n23460,
         n23461, n23462, n23463, n23464, n23465, n23466, n23467, n23468,
         n23469, n23470, n23471, n23472, n23473, n23474, n23475, n23476,
         n23477, n23478, n23479, n23480, n23481, n23482, n23483, n23484,
         n23485, n23486, n23487, n23488, n23489, n23490, n23491, n23492,
         n23493, n23494, n23495, n23496, n23497, n23498, n23499, n23500,
         n23501, n23502, n23503, n23504, n23505, n23506, n23507, n23508,
         n23509, n23510, n23511, n23512, n23513, n23514, n23515, n23516,
         n23517, n23518, n23519, n23520, n23521, n23522, n23523, n23524,
         n23525, n23526, n23527, n23528, n23529, n23530, n23531, n23532,
         n23533, n23534, n23535, n23536, n23537, n23538, n23539, n23540,
         n23541, n23542, n23543, n23544, n23545, n23546, n23547, n23548,
         n23549, n23550, n23551, n23552, n23553, n23554, n23555, n23556,
         n23557, n23558, n23559, n23560, n23561, n23562, n23563, n23564,
         n23565, n23566, n23567, n23568, n23569, n23570, n23571, n23572,
         n23573, n23574, n23575, n23576, n23577, n23578, n23579, n23580,
         n23581, n23582, n23583, n23584, n23585, n23586, n23587, n23588,
         n23589, n23590, n23591, n23592, n23593, n23594, n23595, n23596,
         n23597, n23598, n23599, n23600, n23601, n23602, n23603, n23604,
         n23605, n23606, n23607, n23608, n23609, n23610, n23611, n23612,
         n23613, n23614, n23615, n23616, n23617, n23618, n23619, n23620,
         n23621, n23622, n23623, n23624, n23625, n23626, n23627, n23628,
         n23629, n23630, n23631, n23632, n23633, n23634, n23635, n23636,
         n23637, n23638, n23639, n23640, n23641, n23642, n23643, n23644,
         n23645, n23646, n23647, n23648, n23649, n23650, n23651, n23652,
         n23653, n23654, n23655, n23656, n23657, n23658, n23659, n23660,
         n23661, n23662, n23663, n23664, n23665, n23666, n23667, n23668,
         n23669, n23670, n23671, n23672, n23673, n23674, n23675, n23676,
         n23677, n23678, n23679, n23680, n23681, n23682, n23683, n23684,
         n23685, n23686, n23687, n23688, n23689, n23690, n23691, n23692,
         n23693, n23694, n23695, n23696, n23697, n23698, n23699, n23700,
         n23701, n23702, n23703, n23704, n23705, n23706, n23707, n23708,
         n23709, n23710, n23711, n23712, n23713, n23714, n23715, n23716,
         n23717, n23718, n23719, n23720, n23721, n23722, n23723, n23724,
         n23725, n23726, n23727, n23728, n23729, n23730, n23731, n23732,
         n23733, n23734, n23735, n23736, n23737, n23738, n23739, n23740,
         n23741, n23742, n23743, n23744, n23745, n23746, n23747, n23748,
         n23749, n23750, n23751, n23752, n23753, n23754, n23755, n23756,
         n23757, n23758, n23759, n23760, n23761, n23762, n23763, n23764,
         n23765, n23766, n23767, n23768, n23769, n23770, n23771, n23772,
         n23773, n23774, n23775, n23776, n23777, n23778, n23779, n23780,
         n23781, n23782, n23783, n23784, n23785, n23786, n23787, n23788,
         n23789, n23790, n23791, n23792, n23793, n23794, n23795, n23796,
         n23797, n23798, n23799, n23800, n23801, n23802, n23803, n23804,
         n23805, n23806, n23807, n23808, n23809, n23810, n23811, n23812,
         n23813, n23814, n23815, n23816, n23817, n23818, n23819, n23820,
         n23821, n23822, n23823, n23824, n23825, n23826, n23827, n23828,
         n23829, n23830, n23831, n23832, n23833, n23834, n23835, n23836,
         n23837, n23838, n23839, n23840, n23841, n23842, n23843, n23844,
         n23845, n23846, n23847, n23848, n23849, n23850, n23851, n23852,
         n23853, n23854, n23855, n23856, n23857, n23858, n23859, n23860,
         n23861, n23862, n23863, n23864, n23865, n23866, n23867, n23868,
         n23869, n23870, n23871, n23872, n23873, n23874, n23875, n23876,
         n23877, n23878, n23879, n23880, n23881, n23882, n23883, n23884,
         n23885, n23886, n23887, n23888, n23889, n23890, n23891, n23892,
         n23893, n23894, n23895, n23896, n23897, n23898, n23899, n23900,
         n23901, n23902, n23903, n23904, n23905, n23906, n23907, n23908,
         n23909, n23910, n23911, n23912, n23913, n23914, n23915, n23916,
         n23917, n23918, n23919, n23920, n23921, n23922, n23923, n23924,
         n23925, n23926, n23927, n23928, n23929, n23930, n23931, n23932,
         n23933, n23934, n23935, n23936, n23937, n23938, n23939, n23940,
         n23941, n23942, n23943, n23944, n23945, n23946, n23947, n23948,
         n23949, n23950, n23951, n23952, n23953, n23954, n23955, n23956,
         n23957, n23958, n23959, n23960, n23961, n23962, n23963, n23964,
         n23965, n23966, n23967, n23968, n23969, n23970, n23971, n23972,
         n23973, n23974, n23975, n23976, n23977, n23978, n23979, n23980,
         n23981, n23982, n23983, n23984, n23985, n23986, n23987, n23988,
         n23989, n23990, n23991, n23992, n23993, n23994, n23995, n23996,
         n23997, n23998, n23999, n24000, n24001, n24002, n24003, n24004,
         n24005, n24006, n24007, n24008, n24009, n24010, n24011, n24012,
         n24013, n24014, n24015, n24016, n24017, n24018, n24019, n24020,
         n24021, n24022, n24023, n24024, n24025, n24026, n24027, n24028,
         n24029, n24030, n24031, n24032, n24033, n24034, n24035, n24036,
         n24037, n24038, n24039, n24040, n24041, n24042, n24043, n24044,
         n24045, n24046, n24047, n24048, n24049, n24050, n24051, n24052,
         n24053, n24054, n24055, n24056, n24057, n24058, n24059, n24060,
         n24061, n24062, n24063, n24064, n24065, n24066, n24067, n24068,
         n24069, n24070, n24071, n24072, n24073, n24074, n24075, n24076,
         n24077, n24078, n24079, n24080, n24081, n24082, n24083, n24084,
         n24085, n24086, n24087, n24088, n24089, n24090, n24091, n24092,
         n24093, n24094, n24095, n24096, n24097, n24098, n24099, n24100,
         n24101, n24102, n24103, n24104, n24105, n24106, n24107, n24108,
         n24109, n24110, n24111, n24112, n24113, n24114, n24115, n24116,
         n24117, n24118, n24119, n24120, n24121, n24122, n24123, n24124,
         n24125, n24126, n24127, n24128, n24129, n24130, n24131, n24132,
         n24133, n24134, n24135, n24136, n24137, n24138, n24139, n24140,
         n24141, n24142, n24143, n24144, n24145, n24146, n24147, n24148,
         n24149, n24150, n24151, n24152, n24153, n24154, n24155, n24156,
         n24157, n24158, n24159, n24160, n24161, n24162, n24163, n24164,
         n24165, n24166, n24167, n24168, n24169, n24170, n24171, n24172,
         n24173, n24174, n24175, n24176, n24177, n24178, n24179, n24180,
         n24181, n24182, n24183, n24184, n24185, n24186, n24187, n24188,
         n24189, n24190, n24191, n24192, n24193, n24194, n24195, n24196,
         n24197, n24198, n24199, n24200, n24201, n24202, n24203, n24204,
         n24205, n24206, n24207, n24208, n24209, n24210, n24211, n24212,
         n24213, n24214, n24215, n24216, n24217, n24218, n24219, n24220,
         n24221, n24222, n24223, n24224, n24225, n24226, n24227, n24228,
         n24229, n24230, n24231, n24232, n24233, n24234, n24235, n24236,
         n24237, n24238, n24239, n24240, n24241, n24242, n24243, n24244,
         n24245, n24246, n24247, n24248, n24249, n24250, n24251, n24252,
         n24253, n24254, n24255, n24256, n24257, n24258, n24259, n24260,
         n24261, n24262, n24263, n24264, n24265, n24266, n24267, n24268,
         n24269, n24270, n24271, n24272, n24273, n24274, n24275, n24276,
         n24277, n24278, n24279, n24280, n24281, n24282, n24283, n24284,
         n24285, n24286, n24287, n24288, n24289, n24290, n24291, n24292,
         n24293, n24294, n24295, n24296, n24297, n24298, n24299, n24300,
         n24301, n24302, n24303, n24304, n24305, n24306, n24307, n24308,
         n24309, n24310, n24311, n24312, n24313, n24314, n24315, n24316,
         n24317, n24318, n24319, n24320, n24321, n24322, n24323, n24324,
         n24325, n24326, n24327, n24328, n24329, n24330, n24331, n24332,
         n24333, n24334, n24335, n24336, n24337, n24338, n24339, n24340,
         n24341, n24342, n24343, n24344, n24345, n24346, n24347, n24348,
         n24349, n24350, n24351, n24352, n24353, n24354, n24355, n24356,
         n24357, n24358, n24359, n24360, n24361, n24362, n24363, n24364,
         n24365, n24366, n24367, n24368, n24369, n24370, n24371, n24372,
         n24373, n24374, n24375, n24376, n24377, n24378, n24379, n24380,
         n24381, n24382, n24383, n24384, n24385, n24386, n24387, n24388,
         n24389, n24390, n24391, n24392, n24393, n24394, n24395, n24396,
         n24397, n24398, n24399, n24400, n24401, n24402, n24403, n24404,
         n24405, n24406, n24407, n24408, n24409, n24410, n24411, n24412,
         n24413, n24414, n24415, n24416, n24417, n24418, n24419, n24420,
         n24421, n24422, n24423, n24424, n24425, n24426, n24427, n24428,
         n24429, n24430, n24431, n24432, n24433, n24434, n24435, n24436,
         n24437, n24438, n24439, n24440, n24441, n24442, n24443, n24444,
         n24445, n24446, n24447, n24448, n24449, n24450, n24451, n24452,
         n24453, n24454, n24455, n24456, n24457, n24458, n24459, n24460,
         n24461, n24462, n24463, n24464, n24465, n24466, n24467, n24468,
         n24469, n24470, n24471, n24472, n24473, n24474, n24475, n24476,
         n24477, n24478, n24479, n24480, n24481, n24482, n24483, n24484,
         n24485, n24486, n24487, n24488, n24489, n24490, n24491, n24492,
         n24493, n24494, n24495, n24496, n24497, n24498, n24499, n24500,
         n24501, n24502, n24503, n24504, n24505, n24506, n24507, n24508,
         n24509, n24510, n24511, n24512, n24513, n24514, n24515, n24516,
         n24517, n24518, n24519, n24520, n24521, n24522, n24523, n24524,
         n24525, n24526, n24527, n24528, n24529, n24530, n24531, n24532,
         n24533, n24534, n24535, n24536, n24537, n24538, n24539, n24540,
         n24541, n24542, n24543, n24544, n24545, n24546, n24547, n24548,
         n24549, n24550, n24551, n24552, n24553, n24554, n24555, n24556,
         n24557, n24558, n24559, n24560, n24561, n24562, n24563, n24564,
         n24565, n24566, n24567, n24568, n24569, n24570, n24571, n24572,
         n24573, n24574, n24575, n24576, n24577, n24578, n24579, n24580,
         n24581, n24582, n24583, n24584, n24585, n24586, n24587, n24588,
         n24589, n24590, n24591, n24592, n24593, n24594, n24595, n24596,
         n24597, n24598, n24599, n24600, n24601, n24602, n24603, n24604,
         n24605, n24606, n24607, n24608, n24609, n24610, n24611, n24612,
         n24613, n24614, n24615, n24616, n24617, n24618, n24619, n24620,
         n24621, n24622, n24623, n24624, n24625, n24626, n24627, n24628,
         n24629, n24630, n24631, n24632, n24633, n24634, n24635, n24636,
         n24637, n24638, n24639, n24640, n24641, n24642, n24643, n24644,
         n24645, n24646, n24647, n24648, n24649, n24650, n24651, n24652,
         n24653, n24654, n24655, n24656, n24657, n24658, n24659, n24660,
         n24661, n24662, n24663, n24664, n24665, n24666, n24667, n24668,
         n24669, n24670, n24671, n24672, n24673, n24674, n24675, n24676,
         n24677, n24678, n24679, n24680, n24681, n24682, n24683, n24684,
         n24685, n24686, n24687, n24688, n24689, n24690, n24691, n24692,
         n24693, n24694, n24695, n24696, n24697, n24698, n24699, n24700,
         n24701, n24702, n24703, n24704, n24705, n24706, n24707, n24708,
         n24709, n24710, n24711, n24712, n24713, n24714, n24715, n24716,
         n24717, n24718, n24719, n24720, n24721, n24722, n24723, n24724,
         n24725, n24726, n24727, n24728, n24729, n24730, n24731, n24732,
         n24733, n24734, n24735, n24736, n24737, n24738, n24739, n24740,
         n24741, n24742, n24743, n24744, n24745, n24746, n24747, n24748,
         n24749, n24750, n24751, n24752, n24753, n24754, n24755, n24756,
         n24757, n24758, n24759, n24760, n24761, n24762, n24763, n24764,
         n24765, n24766, n24767, n24768, n24769, n24770, n24771, n24772,
         n24773, n24774, n24775, n24776, n24777, n24778, n24779, n24780,
         n24781, n24782, n24783, n24784, n24785, n24786, n24787, n24788,
         n24789, n24790, n24791, n24792, n24793, n24794, n24795, n24796,
         n24797, n24798, n24799, n24800, n24801, n24802, n24803, n24804,
         n24805, n24806, n24807, n24808, n24809, n24810, n24811, n24812,
         n24813, n24814, n24815, n24816, n24817, n24818, n24819, n24820,
         n24821, n24822, n24823, n24824, n24825, n24826, n24827, n24828,
         n24829, n24830, n24831, n24832, n24833, n24834, n24835, n24836,
         n24837, n24838, n24839, n24840, n24841, n24842, n24843, n24844,
         n24845, n24846, n24847, n24848, n24849, n24850, n24851, n24852,
         n24853, n24854, n24855, n24856, n24857, n24858, n24859, n24860,
         n24861, n24862, n24863, n24864, n24865, n24866, n24867, n24868,
         n24869, n24870, n24871, n24872, n24873, n24874, n24875, n24876,
         n24877, n24878, n24879, n24880, n24881, n24882, n24883, n24884,
         n24885, n24886, n24887, n24888, n24889, n24890, n24891, n24892,
         n24893, n24894, n24895, n24896, n24897, n24898, n24899, n24900,
         n24901, n24902, n24903, n24904, n24905, n24906, n24907, n24908,
         n24909, n24910, n24911, n24912, n24913, n24914, n24915, n24916,
         n24917, n24918, n24919, n24920, n24921, n24922, n24923, n24924,
         n24925, n24926, n24927, n24928, n24929, n24930, n24931, n24932,
         n24933, n24934, n24935, n24936, n24937, n24938, n24939, n24940,
         n24941, n24942, n24943, n24944, n24945, n24946, n24947, n24948,
         n24949, n24950, n24951, n24952, n24953, n24954, n24955, n24956,
         n24957, n24958, n24959, n24960, n24961, n24962, n24963, n24964,
         n24965, n24966, n24967, n24968, n24969, n24970, n24971, n24972,
         n24973, n24974, n24975, n24976, n24977, n24978, n24979, n24980,
         n24981, n24982, n24983, n24984, n24985, n24986, n24987, n24988,
         n24989, n24990, n24991, n24992, n24993, n24994, n24995, n24996,
         n24997, n24998, n24999, n25000, n25001, n25002, n25003, n25004,
         n25005, n25006, n25007, n25008, n25009, n25010, n25011, n25012,
         n25013, n25014, n25015, n25016, n25017, n25018, n25019, n25020,
         n25021, n25022, n25023, n25024, n25025, n25026, n25027, n25028,
         n25029, n25030, n25031, n25032, n25033, n25034, n25035, n25036,
         n25037, n25038, n25039, n25040, n25041, n25042, n25043, n25044,
         n25045, n25046, n25047, n25048, n25049, n25050, n25051, n25052,
         n25053, n25054, n25055, n25056, n25057, n25058, n25059, n25060,
         n25061, n25062, n25063, n25064, n25065, n25066, n25067, n25068,
         n25069, n25070, n25071, n25072, n25073, n25074, n25075, n25076,
         n25077, n25078, n25079, n25080, n25081, n25082, n25083, n25084,
         n25085, n25086, n25087, n25088, n25089, n25090, n25091, n25092,
         n25093, n25094, n25095, n25096, n25097, n25098, n25099, n25100,
         n25101, n25102, n25103, n25104, n25105, n25106, n25107, n25108,
         n25109, n25110, n25111, n25112, n25113, n25114, n25115, n25116,
         n25117, n25118, n25119, n25120, n25121, n25122, n25123, n25124,
         n25125, n25126, n25127, n25128, n25129, n25130, n25131, n25132,
         n25133, n25134, n25135, n25136, n25137, n25138, n25139, n25140,
         n25141, n25142, n25143, n25144, n25145, n25146, n25147, n25148,
         n25149, n25150, n25151, n25152, n25153, n25154, n25155, n25156,
         n25157, n25158, n25159, n25160, n25161, n25162, n25163, n25164,
         n25165, n25166, n25167, n25168, n25169, n25170, n25171, n25172,
         n25173, n25174, n25175, n25176, n25177, n25178, n25179, n25180,
         n25181, n25182, n25183, n25184, n25185, n25186, n25187, n25188,
         n25189, n25190, n25191, n25192, n25193, n25194, n25195, n25196,
         n25197, n25198, n25199, n25200, n25201, n25202, n25203, n25204,
         n25205, n25206, n25207, n25208, n25209, n25210, n25211, n25212,
         n25213, n25214, n25215, n25216, n25217, n25218, n25219, n25220,
         n25221, n25222, n25223, n25224, n25225, n25226, n25227, n25228,
         n25229, n25230, n25231, n25232, n25233, n25234, n25235, n25236,
         n25237, n25238, n25239, n25240, n25241, n25242, n25243, n25244,
         n25245, n25246, n25247, n25248, n25249, n25250, n25251, n25252,
         n25253, n25254, n25255, n25256, n25257, n25258, n25259, n25260,
         n25261, n25262, n25263, n25264, n25265, n25266, n25267, n25268,
         n25269, n25270, n25271, n25272, n25273, n25274, n25275, n25276,
         n25277, n25278, n25279, n25280, n25281, n25282, n25283, n25284,
         n25285, n25286, n25287, n25288, n25289, n25290, n25291, n25292,
         n25293, n25294, n25295, n25296, n25297, n25298, n25299, n25300,
         n25301, n25302, n25303, n25304, n25305, n25306, n25307, n25308,
         n25309, n25310, n25311, n25312, n25313, n25314, n25315, n25316,
         n25317, n25318, n25319, n25320, n25321, n25322, n25323, n25324,
         n25325, n25326, n25327, n25328, n25329, n25330, n25331, n25332,
         n25333, n25334, n25335, n25336, n25337, n25338, n25339, n25340,
         n25341, n25342, n25343, n25344, n25345, n25346, n25347, n25348,
         n25349, n25350, n25351, n25352, n25353, n25354, n25355, n25356,
         n25357, n25358, n25359, n25360, n25361, n25362, n25363, n25364,
         n25365, n25366, n25367, n25368, n25369, n25370, n25371, n25372,
         n25373, n25374, n25375, n25376, n25377, n25378, n25379, n25380,
         n25381, n25382, n25383, n25384, n25385, n25386, n25387, n25388,
         n25389, n25390, n25391, n25392, n25393, n25394, n25395, n25396,
         n25397, n25398, n25399, n25400, n25401, n25402, n25403, n25404,
         n25405, n25406, n25407, n25408, n25409, n25410, n25411, n25412,
         n25413, n25414, n25415, n25416, n25417, n25418, n25419, n25420,
         n25421, n25422, n25423, n25424, n25425, n25426, n25427, n25428,
         n25429, n25430, n25431, n25432, n25433, n25434, n25435, n25436,
         n25437, n25438, n25439, n25440, n25441, n25442, n25443, n25444,
         n25445, n25446, n25447, n25448, n25449, n25450, n25451, n25452,
         n25453, n25454, n25455, n25456, n25457, n25458, n25459, n25460,
         n25461, n25462, n25463, n25464, n25465, n25466, n25467, n25468,
         n25469, n25470, n25471, n25472, n25473, n25474, n25475, n25476,
         n25477, n25478, n25479, n25480, n25481, n25482, n25483, n25484,
         n25485, n25486, n25487, n25488, n25489, n25490, n25491, n25492,
         n25493, n25494, n25495, n25496, n25497, n25498, n25499, n25500,
         n25501, n25502, n25503, n25504, n25505, n25506, n25507, n25508,
         n25509, n25510, n25511, n25512, n25513, n25514, n25515, n25516,
         n25517, n25518, n25519, n25520, n25521, n25522, n25523, n25524,
         n25525, n25526, n25527, n25528, n25529, n25530, n25531, n25532,
         n25533, n25534, n25535, n25536, n25537, n25538, n25539, n25540,
         n25541, n25542, n25543, n25544, n25545, n25546, n25547, n25548,
         n25549, n25550, n25551, n25552, n25553, n25554, n25555, n25556,
         n25557, n25558, n25559, n25560, n25561, n25562, n25563, n25564,
         n25565, n25566, n25567, n25568, n25569, n25570, n25571, n25572,
         n25573, n25574, n25575, n25576, n25577, n25578, n25579, n25580,
         n25581, n25582, n25583, n25584, n25585, n25586, n25587, n25588,
         n25589, n25590, n25591, n25592, n25593, n25594, n25595, n25596,
         n25597, n25598, n25599, n25600, n25601, n25602, n25603, n25604,
         n25605, n25606, n25607, n25608, n25609, n25610, n25611, n25612,
         n25613, n25614, n25615, n25616, n25617, n25618, n25619, n25620,
         n25621, n25622, n25623, n25624, n25625, n25626, n25627, n25628,
         n25629, n25630, n25631, n25632, n25633, n25634, n25635, n25636,
         n25637, n25638, n25639, n25640, n25641, n25642, n25643, n25644,
         n25645, n25646, n25647, n25648, n25649, n25650, n25651, n25652,
         n25653, n25654, n25655, n25656, n25657, n25658, n25659, n25660,
         n25661, n25662, n25663, n25664, n25665, n25666, n25667, n25668,
         n25669, n25670, n25671, n25672, n25673, n25674, n25675, n25676,
         n25677, n25678, n25679, n25680, n25681, n25682, n25683, n25684,
         n25685, n25686, n25687, n25688, n25689, n25690, n25691, n25692,
         n25693, n25694, n25695, n25696, n25697, n25698, n25699, n25700,
         n25701, n25702, n25703, n25704, n25705, n25706, n25707, n25708,
         n25709, n25710, n25711, n25712, n25713, n25714, n25715, n25716,
         n25717, n25718, n25719, n25720, n25721, n25722, n25723, n25724,
         n25725, n25726, n25727, n25728, n25729, n25730, n25731, n25732,
         n25733, n25734, n25735, n25736, n25737, n25738, n25739, n25740,
         n25741, n25742, n25743, n25744, n25745, n25746, n25747, n25748,
         n25749, n25750, n25751, n25752, n25753, n25754, n25755, n25756,
         n25757, n25758, n25759, n25760, n25761, n25762, n25763, n25764,
         n25765, n25766, n25767, n25768, n25769, n25770, n25771, n25772,
         n25773, n25774, n25775, n25776, n25777, n25778, n25779, n25780,
         n25781, n25782, n25783, n25784, n25785, n25786, n25787, n25788,
         n25789, n25790, n25791, n25792, n25793, n25794, n25795, n25796,
         n25797, n25798, n25799, n25800, n25801, n25802, n25803, n25804,
         n25805, n25806, n25807, n25808, n25809, n25810, n25811, n25812,
         n25813, n25814, n25815, n25816, n25817, n25818, n25819, n25820,
         n25821, n25822, n25823, n25824, n25825, n25826, n25827, n25828,
         n25829, n25830, n25831, n25832, n25833, n25834, n25835, n25836,
         n25837, n25838, n25839, n25840, n25841, n25842, n25843, n25844,
         n25845, n25846, n25847, n25848, n25849, n25850, n25851, n25852,
         n25853, n25854, n25855, n25856, n25857, n25858, n25859, n25860,
         n25861, n25862, n25863, n25864, n25865, n25866, n25867, n25868,
         n25869, n25870, n25871, n25872, n25873, n25874, n25875, n25876,
         n25877, n25878, n25879, n25880, n25881, n25882, n25883, n25884,
         n25885, n25886, n25887, n25888, n25889, n25890, n25891, n25892,
         n25893, n25894, n25895, n25896, n25897, n25898, n25899, n25900,
         n25901, n25902, n25903, n25904, n25905, n25906, n25907, n25908,
         n25909, n25910, n25911, n25912, n25913, n25914, n25915, n25916,
         n25917, n25918, n25919, n25920, n25921, n25922, n25923, n25924,
         n25925, n25926, n25927, n25928, n25929, n25930, n25931, n25932,
         n25933, n25934, n25935, n25936, n25937, n25938, n25939, n25940,
         n25941, n25942, n25943, n25944, n25945, n25946, n25947, n25948,
         n25949, n25950, n25951, n25952, n25953, n25954, n25955, n25956,
         n25957, n25958, n25959, n25960, n25961, n25962, n25963, n25964,
         n25965, n25966, n25967, n25968, n25969, n25970, n25971, n25972,
         n25973, n25974, n25975, n25976, n25977, n25978, n25979, n25980,
         n25981, n25982, n25983, n25984, n25985, n25986, n25987, n25988,
         n25989, n25990, n25991, n25992, n25993, n25994, n25995, n25996,
         n25997, n25998, n25999, n26000, n26001, n26002, n26003, n26004,
         n26005, n26006, n26007, n26008, n26009, n26010, n26011, n26012,
         n26013, n26014, n26015, n26016, n26017, n26018, n26019, n26020,
         n26021, n26022, n26023, n26024, n26025, n26026, n26027, n26028,
         n26029, n26030, n26031, n26032, n26033, n26034, n26035, n26036,
         n26037, n26038, n26039, n26040, n26041, n26042, n26043, n26044,
         n26045, n26046, n26047, n26048, n26049, n26050, n26051, n26052,
         n26053, n26054, n26055, n26056, n26057, n26058, n26059, n26060,
         n26061, n26062, n26063, n26064, n26065, n26066, n26067, n26068,
         n26069, n26070, n26071, n26072, n26073, n26074, n26075, n26076,
         n26077, n26078, n26079, n26080, n26081, n26082, n26083, n26084,
         n26085, n26086, n26087, n26088, n26089, n26090, n26091, n26092,
         n26093, n26094, n26095, n26096, n26097, n26098, n26099, n26100,
         n26101, n26102, n26103, n26104, n26105, n26106, n26107, n26108,
         n26109, n26110, n26111, n26112, n26113, n26114, n26115, n26116,
         n26117, n26118, n26119, n26120, n26121, n26122, n26123, n26124,
         n26125, n26126, n26127, n26128, n26129, n26130, n26131, n26132,
         n26133, n26134, n26135, n26136, n26137, n26138, n26139, n26140,
         n26141, n26142, n26143, n26144, n26145, n26146, n26147, n26148,
         n26149, n26150, n26151, n26152, n26153, n26154, n26155, n26156,
         n26157, n26158, n26159, n26160, n26161, n26162, n26163, n26164,
         n26165, n26166, n26167, n26168, n26169, n26170, n26171, n26172,
         n26173, n26174, n26175, n26176, n26177, n26178, n26179, n26180,
         n26181, n26182, n26183, n26184, n26185, n26186, n26187, n26188,
         n26189, n26190, n26191, n26192, n26193, n26194, n26195, n26196,
         n26197, n26198, n26199, n26200, n26201, n26202, n26203, n26204,
         n26205, n26206, n26207, n26208, n26209, n26210, n26211, n26212,
         n26213, n26214, n26215, n26216, n26217, n26218, n26219, n26220,
         n26221, n26222, n26223, n26224, n26225, n26226, n26227, n26228,
         n26229, n26230, n26231, n26232, n26233, n26234, n26235, n26236,
         n26237, n26238, n26239, n26240, n26241, n26242, n26243, n26244,
         n26245, n26246, n26247, n26248, n26249, n26250, n26251, n26252,
         n26253, n26254, n26255, n26256, n26257, n26258, n26259, n26260,
         n26261, n26262, n26263, n26264, n26265, n26266, n26267, n26268,
         n26269, n26270, n26271, n26272, n26273, n26274, n26275, n26276,
         n26277, n26278, n26279, n26280, n26281, n26282, n26283, n26284,
         n26285, n26286, n26287, n26288, n26289, n26290, n26291, n26292,
         n26293, n26294, n26295, n26296, n26297, n26298, n26299, n26300,
         n26301, n26302, n26303, n26304, n26305, n26306, n26307, n26308,
         n26309, n26310, n26311, n26312, n26313, n26314, n26315, n26316,
         n26317, n26318, n26319, n26320, n26321, n26322, n26323, n26324,
         n26325, n26326, n26327, n26328, n26329, n26330, n26331, n26332,
         n26333, n26334, n26335, n26336, n26337, n26338, n26339, n26340,
         n26341, n26342, n26343, n26344, n26345, n26346, n26347, n26348,
         n26349, n26350, n26351, n26352, n26353, n26354, n26355, n26356,
         n26357, n26358, n26359, n26360, n26361, n26362, n26363, n26364,
         n26365, n26366, n26367, n26368, n26369, n26370, n26371, n26372,
         n26373, n26374, n26375, n26376, n26377, n26378, n26379, n26380,
         n26381, n26382, n26383, n26384, n26385, n26386, n26387, n26388,
         n26389, n26390, n26391, n26392, n26393, n26394, n26395, n26396,
         n26397, n26398, n26399, n26400, n26401, n26402, n26403, n26404,
         n26405, n26406, n26407, n26408, n26409, n26410, n26411, n26412,
         n26413, n26414, n26415, n26416, n26417, n26418, n26419, n26420,
         n26421, n26422, n26423, n26424, n26425, n26426, n26427, n26428,
         n26429, n26430, n26431, n26432, n26433, n26434, n26435, n26436,
         n26437, n26438, n26439, n26440, n26441, n26442, n26443, n26444,
         n26445, n26446, n26447, n26448, n26449, n26450, n26451, n26452,
         n26453, n26454, n26455, n26456, n26457, n26458, n26459, n26460,
         n26461, n26462, n26463, n26464, n26465, n26466, n26467, n26468,
         n26469, n26470, n26471, n26472, n26473, n26474, n26475, n26476,
         n26477, n26478, n26479, n26480, n26481, n26482, n26483, n26484,
         n26485, n26486, n26487, n26488, n26489, n26490, n26491, n26492,
         n26493, n26494, n26495, n26496, n26497, n26498, n26499, n26500,
         n26501, n26502, n26503, n26504, n26505, n26506, n26507, n26508,
         n26509, n26510, n26511, n26512, n26513, n26514, n26515, n26516,
         n26517, n26518, n26519, n26520, n26521, n26522, n26523, n26524,
         n26525, n26526, n26527, n26528, n26529, n26530, n26531, n26532,
         n26533, n26534, n26535, n26536, n26537, n26538, n26539, n26540,
         n26541, n26542, n26543, n26544, n26545, n26546, n26547, n26548,
         n26549, n26550, n26551, n26552, n26553, n26554, n26555, n26556,
         n26557, n26558, n26559, n26560, n26561, n26562, n26563, n26564,
         n26565, n26566, n26567, n26568, n26569, n26570, n26571, n26572,
         n26573, n26574, n26575, n26576, n26577, n26578, n26579, n26580,
         n26581, n26582, n26583, n26584, n26585, n26586, n26587, n26588,
         n26589, n26590, n26591, n26592, n26593, n26594, n26595, n26596,
         n26597, n26598, n26599, n26600, n26601, n26602, n26603, n26604,
         n26605, n26606, n26607, n26608, n26609, n26610, n26611, n26612,
         n26613, n26614, n26615, n26616, n26617, n26618, n26619, n26620,
         n26621, n26622, n26623, n26624, n26625, n26626, n26627, n26628,
         n26629, n26630, n26631, n26632, n26633, n26634, n26635, n26636,
         n26637, n26638, n26639, n26640, n26641, n26642, n26643, n26644,
         n26645, n26646, n26647, n26648, n26649, n26650, n26651, n26652,
         n26653, n26654, n26655, n26656, n26657, n26658, n26659, n26660,
         n26661, n26662, n26663, n26664, n26665, n26666, n26667, n26668,
         n26669, n26670, n26671, n26672, n26673, n26674, n26675, n26676,
         n26677, n26678, n26679, n26680, n26681, n26682, n26683, n26684,
         n26685, n26686, n26687, n26688, n26689, n26690, n26691, n26692,
         n26693, n26694, n26695, n26696, n26697, n26698, n26699, n26700,
         n26701, n26702, n26703, n26704, n26705, n26706, n26707, n26708,
         n26709, n26710, n26711, n26712, n26713, n26714, n26715, n26716,
         n26717, n26718, n26719, n26720, n26721, n26722, n26723, n26724,
         n26725, n26726, n26727, n26728, n26729, n26730, n26731, n26732,
         n26733, n26734, n26735, n26736, n26737, n26738, n26739, n26740,
         n26741, n26742, n26743, n26744, n26745, n26746, n26747, n26748,
         n26749, n26750, n26751, n26752, n26753, n26754, n26755, n26756,
         n26757, n26758, n26759, n26760, n26761, n26762, n26763, n26764,
         n26765, n26766, n26767, n26768, n26769, n26770, n26771, n26772,
         n26773, n26774, n26775, n26776, n26777, n26778, n26779, n26780,
         n26781, n26782, n26783, n26784, n26785, n26786, n26787, n26788,
         n26789, n26790, n26791, n26792, n26793, n26794, n26795, n26796,
         n26797, n26798, n26799, n26800, n26801, n26802, n26803, n26804,
         n26805, n26806, n26807, n26808, n26809, n26810, n26811, n26812,
         n26813, n26814, n26815, n26816, n26817, n26818, n26819, n26820,
         n26821, n26822, n26823, n26824, n26825, n26826, n26827, n26828,
         n26829, n26830, n26831, n26832, n26833, n26834, n26835, n26836,
         n26837, n26838, n26839, n26840, n26841, n26842, n26843, n26844,
         n26845, n26846, n26847, n26848, n26849, n26850, n26851, n26852,
         n26853, n26854, n26855, n26856, n26857, n26858, n26859, n26860,
         n26861, n26862, n26863, n26864, n26865, n26866, n26867, n26868,
         n26869, n26870, n26871, n26872, n26873, n26874, n26875, n26876,
         n26877, n26878, n26879, n26880, n26881, n26882, n26883, n26884,
         n26885, n26886, n26887, n26888, n26889, n26890, n26891, n26892,
         n26893, n26894, n26895, n26896, n26897, n26898, n26899, n26900,
         n26901, n26902, n26903, n26904, n26905, n26906, n26907, n26908,
         n26909, n26910, n26911, n26912, n26913, n26914, n26915, n26916,
         n26917, n26918, n26919, n26920, n26921, n26922, n26923, n26924,
         n26925, n26926, n26927, n26928, n26929, n26930, n26931, n26932,
         n26933, n26934, n26935, n26936, n26937, n26938, n26939, n26940,
         n26941, n26942, n26943, n26944, n26945, n26946, n26947, n26948,
         n26949, n26950, n26951, n26952, n26953, n26954, n26955, n26956,
         n26957, n26958, n26959, n26960, n26961, n26962, n26963, n26964,
         n26965, n26966, n26967, n26968, n26969, n26970, n26971, n26972,
         n26973, n26974, n26975, n26976, n26977, n26978, n26979, n26980,
         n26981, n26982, n26983, n26984, n26985, n26986, n26987, n26988,
         n26989, n26990, n26991, n26992, n26993, n26994, n26995, n26996,
         n26997, n26998, n26999, n27000, n27001, n27002, n27003, n27004,
         n27005, n27006, n27007, n27008, n27009, n27010, n27011, n27012,
         n27013, n27014, n27015, n27016, n27017, n27018, n27019, n27020,
         n27021, n27022, n27023, n27024, n27025, n27026, n27027, n27028,
         n27029, n27030, n27031, n27032, n27033, n27034, n27035, n27036,
         n27037, n27038, n27039, n27040, n27041, n27042, n27043, n27044,
         n27045, n27046, n27047, n27048, n27049, n27050, n27051, n27052,
         n27053, n27054, n27055, n27056, n27057, n27058, n27059, n27060,
         n27061, n27062, n27063, n27064, n27065, n27066, n27067, n27068,
         n27069, n27070, n27071, n27072, n27073, n27074, n27075, n27076,
         n27077, n27078, n27079, n27080, n27081, n27082, n27083, n27084,
         n27085, n27086, n27087, n27088, n27089, n27090, n27091, n27092,
         n27093, n27094, n27095, n27096, n27097, n27098, n27099, n27100,
         n27101, n27102, n27103, n27104, n27105, n27106, n27107, n27108,
         n27109, n27110, n27111, n27112, n27113, n27114, n27115, n27116,
         n27117, n27118, n27119, n27120, n27121, n27122, n27123, n27124,
         n27125, n27126, n27127, n27128, n27129, n27130, n27131, n27132,
         n27133, n27134, n27135, n27136, n27137, n27138, n27139, n27140,
         n27141, n27142, n27143, n27144, n27145, n27146, n27147, n27148,
         n27149, n27150, n27151, n27152, n27153, n27154, n27155, n27156,
         n27157, n27158, n27159, n27160, n27161, n27162, n27163, n27164,
         n27165, n27166, n27167, n27168, n27169, n27170, n27171, n27172,
         n27173, n27174, n27175, n27176, n27177, n27178, n27179, n27180,
         n27181, n27182, n27183, n27184, n27185, n27186, n27187, n27188,
         n27189, n27190, n27191, n27192, n27193, n27194, n27195, n27196,
         n27197, n27198, n27199, n27200, n27201, n27202, n27203, n27204,
         n27205, n27206, n27207, n27208, n27209, n27210, n27211, n27212,
         n27213, n27214, n27215, n27216, n27217, n27218, n27219, n27220,
         n27221, n27222, n27223, n27224, n27225, n27226, n27227, n27228,
         n27229, n27230, n27231, n27232, n27233, n27234, n27235, n27236,
         n27237, n27238, n27239, n27240, n27241, n27242, n27243, n27244,
         n27245, n27246, n27247, n27248, n27249, n27250, n27251, n27252,
         n27253, n27254, n27255, n27256, n27257, n27258, n27259, n27260,
         n27261, n27262, n27263, n27264, n27265, n27266, n27267, n27268,
         n27269, n27270, n27271, n27272, n27273, n27274, n27275, n27276,
         n27277, n27278, n27279, n27280, n27281, n27282, n27283, n27284,
         n27285, n27286, n27287, n27288, n27289, n27290, n27291, n27292,
         n27293, n27294, n27295, n27296, n27297, n27298, n27299, n27300,
         n27301, n27302, n27303, n27304, n27305, n27306, n27307, n27308,
         n27309, n27310, n27311, n27312, n27313, n27314, n27315, n27316,
         n27317, n27318, n27319, n27320, n27321, n27322, n27323, n27324,
         n27325, n27326, n27327, n27328, n27329, n27330, n27331, n27332,
         n27333, n27334, n27335, n27336, n27337, n27338, n27339, n27340,
         n27341, n27342, n27343, n27344, n27345, n27346, n27347, n27348,
         n27349, n27350, n27351, n27352, n27353, n27354, n27355, n27356,
         n27357, n27358, n27359, n27360, n27361, n27362, n27363, n27364,
         n27365, n27366, n27367, n27368, n27369, n27370, n27371, n27372,
         n27373, n27374, n27375, n27376, n27377, n27378, n27379, n27380,
         n27381, n27382, n27383, n27384, n27385, n27386, n27387, n27388,
         n27389, n27390, n27391, n27392, n27393, n27394, n27395, n27396,
         n27397, n27398, n27399, n27400, n27401, n27402, n27403, n27404,
         n27405, n27406, n27407, n27408, n27409, n27410, n27411, n27412,
         n27413, n27414, n27415, n27416, n27417, n27418, n27419, n27420,
         n27421, n27422, n27423, n27424, n27425, n27426, n27427, n27428,
         n27429, n27430, n27431, n27432, n27433, n27434, n27435, n27436,
         n27437, n27438, n27439, n27440, n27441, n27442, n27443, n27444,
         n27445, n27446, n27447, n27448, n27449, n27450, n27451, n27452,
         n27453, n27454, n27455, n27456, n27457, n27458, n27459, n27460,
         n27461, n27462, n27463, n27464, n27465, n27466, n27467, n27468,
         n27469, n27470, n27471, n27472, n27473, n27474, n27475, n27476,
         n27477, n27478, n27479, n27480, n27481, n27482, n27483, n27484,
         n27485, n27486, n27487, n27488, n27489, n27490, n27491, n27492,
         n27493, n27494, n27495, n27496, n27497, n27498, n27499, n27500,
         n27501, n27502, n27503, n27504, n27505, n27506, n27507, n27508,
         n27509, n27510, n27511, n27512, n27513, n27514, n27515, n27516,
         n27517, n27518, n27519, n27520, n27521, n27522, n27523, n27524,
         n27525, n27526, n27527, n27528, n27529, n27530, n27531, n27532,
         n27533, n27534, n27535, n27536, n27537, n27538, n27539, n27540,
         n27541, n27542, n27543, n27544, n27545, n27546, n27547, n27548,
         n27549, n27550, n27551, n27552, n27553, n27554, n27555, n27556,
         n27557, n27558, n27559, n27560, n27561, n27562, n27563, n27564,
         n27565, n27566, n27567, n27568, n27569, n27570, n27571, n27572,
         n27573, n27574, n27575, n27576, n27577, n27578, n27579, n27580,
         n27581, n27582, n27583, n27584, n27585, n27586, n27587, n27588,
         n27589, n27590, n27591, n27592, n27593, n27594, n27595, n27596,
         n27597, n27598, n27599, n27600, n27601, n27602, n27603, n27604,
         n27605, n27606, n27607, n27608, n27609, n27610, n27611, n27612,
         n27613, n27614, n27615, n27616, n27617, n27618, n27619, n27620,
         n27621, n27622, n27623, n27624, n27625, n27626, n27627, n27628,
         n27629, n27630, n27631, n27632, n27633, n27634, n27635, n27636,
         n27637, n27638, n27639, n27640, n27641, n27642, n27643, n27644,
         n27645, n27646, n27647, n27648, n27649, n27650, n27651, n27652,
         n27653, n27654, n27655, n27656, n27657, n27658, n27659, n27660,
         n27661, n27662, n27663, n27664, n27665, n27666, n27667, n27668,
         n27669, n27670, n27671, n27672, n27673, n27674, n27675, n27676,
         n27677, n27678, n27679, n27680, n27681, n27682, n27683, n27684,
         n27685, n27686, n27687, n27688, n27689, n27690, n27691, n27692,
         n27693, n27694, n27695, n27696, n27697, n27698, n27699, n27700,
         n27701, n27702, n27703, n27704, n27705, n27706, n27707, n27708,
         n27709, n27710, n27711, n27712, n27713, n27714, n27715, n27716,
         n27717, n27718, n27719, n27720, n27721, n27722, n27723, n27724,
         n27725, n27726, n27727, n27728, n27729, n27730, n27731, n27732,
         n27733, n27734, n27735, n27736, n27737, n27738, n27739, n27740,
         n27741, n27742, n27743, n27744, n27745, n27746, n27747, n27748,
         n27749, n27750, n27751, n27752, n27753, n27754, n27755, n27756,
         n27757, n27758, n27759, n27760, n27761, n27762, n27763, n27764,
         n27765, n27766, n27767, n27768, n27769, n27770, n27771, n27772,
         n27773, n27774, n27775, n27776, n27777, n27778, n27779, n27780,
         n27781, n27782, n27783, n27784, n27785, n27786, n27787, n27788,
         n27789, n27790, n27791, n27792, n27793, n27794, n27795, n27796,
         n27797, n27798, n27799, n27800, n27801, n27802, n27803, n27804,
         n27805, n27806, n27807, n27808, n27809, n27810, n27811, n27812,
         n27813, n27814, n27815, n27816, n27817, n27818, n27819, n27820,
         n27821, n27822, n27823, n27824, n27825, n27826, n27827, n27828,
         n27829, n27830, n27831, n27832, n27833, n27834, n27835, n27836,
         n27837, n27838, n27839, n27840, n27841, n27842, n27843, n27844,
         n27845, n27846, n27847, n27848, n27849, n27850, n27851, n27852,
         n27853, n27854, n27855, n27856, n27857, n27858, n27859, n27860,
         n27861, n27862, n27863, n27864, n27865, n27866, n27867, n27868,
         n27869, n27870, n27871, n27872, n27873, n27874, n27875, n27876,
         n27877, n27878, n27879, n27880, n27881, n27882, n27883, n27884,
         n27885, n27886, n27887, n27888, n27889, n27890, n27891, n27892,
         n27893, n27894, n27895, n27896, n27897, n27898, n27899, n27900,
         n27901, n27902, n27903, n27904, n27905, n27906, n27907, n27908,
         n27909, n27910, n27911, n27912, n27913, n27914, n27915, n27916,
         n27917, n27918, n27919, n27920, n27921, n27922, n27923, n27924,
         n27925, n27926, n27927, n27928, n27929, n27930, n27931, n27932,
         n27933, n27934, n27935, n27936, n27937, n27938, n27939, n27940,
         n27941, n27942, n27943, n27944, n27945, n27946, n27947, n27948,
         n27949, n27950, n27951, n27952, n27953, n27954, n27955, n27956,
         n27957, n27958, n27959, n27960, n27961, n27962, n27963, n27964,
         n27965, n27966, n27967, n27968, n27969, n27970, n27971, n27972,
         n27973, n27974, n27975, n27976, n27977, n27978, n27979, n27980,
         n27981, n27982, n27983, n27984, n27985, n27986, n27987, n27988,
         n27989, n27990, n27991, n27992, n27993, n27994, n27995, n27996,
         n27997, n27998, n27999, n28000, n28001, n28002, n28003, n28004,
         n28005, n28006, n28007, n28008, n28009, n28010, n28011, n28012,
         n28013, n28014, n28015, n28016, n28017, n28018, n28019, n28020,
         n28021, n28022, n28023, n28024, n28025, n28026, n28027, n28028,
         n28029, n28030, n28031, n28032, n28033, n28034, n28035, n28036,
         n28037, n28038, n28039, n28040, n28041, n28042, n28043, n28044,
         n28045, n28046, n28047, n28048, n28049, n28050, n28051, n28052,
         n28053, n28054, n28055, n28056, n28057, n28058, n28059, n28060,
         n28061, n28062, n28063, n28064, n28065, n28066, n28067, n28068,
         n28069, n28070, n28071, n28072, n28073, n28074, n28075, n28076,
         n28077, n28078, n28079, n28080, n28081, n28082, n28083, n28084,
         n28085, n28086, n28087, n28088, n28089, n28090, n28091, n28092,
         n28093, n28094, n28095, n28096, n28097, n28098, n28099, n28100,
         n28101, n28102, n28103, n28104, n28105, n28106, n28107, n28108,
         n28109, n28110, n28111, n28112, n28113, n28114, n28115, n28116,
         n28117, n28118, n28119, n28120, n28121, n28122, n28123, n28124,
         n28125, n28126, n28127, n28128, n28129, n28130, n28131, n28132,
         n28133, n28134, n28135, n28136, n28137, n28138, n28139, n28140,
         n28141, n28142, n28143, n28144, n28145, n28146, n28147, n28148,
         n28149, n28150, n28151, n28152, n28153, n28154, n28155, n28156,
         n28157, n28158, n28159, n28160, n28161, n28162, n28163, n28164,
         n28165, n28166, n28167, n28168, n28169, n28170, n28171, n28172,
         n28173, n28174, n28175, n28176, n28177, n28178, n28179, n28180,
         n28181, n28182, n28183, n28184, n28185, n28186, n28187, n28188,
         n28189, n28190, n28191, n28192, n28193, n28194, n28195, n28196,
         n28197, n28198, n28199, n28200, n28201, n28202, n28203, n28204,
         n28205, n28206, n28207, n28208, n28209, n28210, n28211, n28212,
         n28213, n28214, n28215, n28216, n28217, n28218, n28219, n28220,
         n28221, n28222, n28223, n28224, n28225, n28226, n28227, n28228,
         n28229, n28230, n28231, n28232, n28233, n28234, n28235, n28236,
         n28237, n28238, n28239, n28240, n28241, n28242, n28243, n28244,
         n28245, n28246, n28247, n28248, n28249, n28250, n28251, n28252,
         n28253, n28254, n28255, n28256, n28257, n28258, n28259, n28260,
         n28261, n28262, n28263, n28264, n28265, n28266, n28267, n28268,
         n28269, n28270, n28271, n28272, n28273, n28274, n28275, n28276,
         n28277, n28278, n28279, n28280, n28281, n28282, n28283, n28284,
         n28285, n28286, n28287, n28288, n28289, n28290, n28291, n28292,
         n28293, n28294, n28295, n28296, n28297, n28298, n28299, n28300,
         n28301, n28302, n28303, n28304, n28305, n28306, n28307, n28308,
         n28309, n28310, n28311, n28312, n28313, n28314, n28315, n28316,
         n28317, n28318, n28319, n28320, n28321, n28322, n28323, n28324,
         n28325, n28326, n28327, n28328, n28329, n28330, n28331, n28332,
         n28333, n28334, n28335, n28336, n28337, n28338, n28339, n28340,
         n28341, n28342, n28343, n28344, n28345, n28346, n28347, n28348,
         n28349, n28350, n28351, n28352, n28353, n28354, n28355, n28356,
         n28357, n28358, n28359, n28360, n28361, n28362, n28363, n28364,
         n28365, n28366, n28367, n28368, n28369, n28370, n28371, n28372,
         n28373, n28374, n28375, n28376, n28377, n28378, n28379, n28380,
         n28381, n28382, n28383, n28384, n28385, n28386, n28387, n28388,
         n28389, n28390, n28391, n28392, n28393, n28394, n28395, n28396,
         n28397, n28398, n28399, n28400, n28401, n28402, n28403, n28404,
         n28405, n28406, n28407, n28408, n28409, n28410, n28411, n28412,
         n28413, n28414, n28415, n28416, n28417, n28418, n28419, n28420,
         n28421, n28422, n28423, n28424, n28425, n28426, n28427, n28428,
         n28429, n28430, n28431, n28432, n28433, n28434, n28435, n28436,
         n28437, n28438, n28439, n28440, n28441, n28442, n28443, n28444,
         n28445, n28446, n28447, n28448, n28449, n28450, n28451, n28452,
         n28453, n28454, n28455, n28456, n28457, n28458, n28459, n28460,
         n28461, n28462, n28463, n28464, n28465, n28466, n28467, n28468,
         n28469, n28470, n28471, n28472, n28473, n28474, n28475, n28476,
         n28477, n28478, n28479, n28480, n28481, n28482, n28483, n28484,
         n28485, n28486, n28487, n28488, n28489, n28490, n28491, n28492,
         n28493, n28494, n28495, n28496, n28497, n28498, n28499, n28500,
         n28501, n28502, n28503, n28504, n28505, n28506, n28507, n28508,
         n28509, n28510, n28511, n28512, n28513, n28514, n28515, n28516,
         n28517, n28518, n28519, n28520, n28521, n28522, n28523, n28524,
         n28525, n28526, n28527, n28528, n28529, n28530, n28531, n28532,
         n28533, n28534, n28535, n28536, n28537, n28538, n28539, n28540,
         n28541, n28542, n28543, n28544, n28545, n28546, n28547, n28548,
         n28549, n28550, n28551, n28552, n28553, n28554, n28555, n28556,
         n28557, n28558, n28559, n28560, n28561, n28562, n28563, n28564,
         n28565, n28566, n28567, n28568, n28569, n28570, n28571, n28572,
         n28573, n28574, n28575, n28576, n28577, n28578, n28579, n28580,
         n28581, n28582, n28583, n28584, n28585, n28586, n28587, n28588,
         n28589, n28590, n28591, n28592, n28593, n28594, n28595, n28596,
         n28597, n28598, n28599, n28600, n28601, n28602, n28603, n28604,
         n28605, n28606, n28607, n28608, n28609, n28610, n28611, n28612,
         n28613, n28614, n28615, n28616, n28617, n28618, n28619, n28620,
         n28621, n28622, n28623, n28624, n28625, n28626, n28627, n28628,
         n28629, n28630, n28631, n28632, n28633, n28634, n28635, n28636,
         n28637, n28638, n28639, n28640, n28641, n28642, n28643, n28644,
         n28645, n28646, n28647, n28648, n28649, n28650, n28651, n28652,
         n28653, n28654, n28655, n28656, n28657, n28658, n28659, n28660,
         n28661, n28662, n28663, n28664, n28665, n28666, n28667, n28668,
         n28669, n28670, n28671, n28672, n28673, n28674, n28675, n28676,
         n28677, n28678, n28679, n28680, n28681, n28682, n28683, n28684,
         n28685, n28686, n28687, n28688, n28689, n28690, n28691, n28692,
         n28693, n28694, n28695, n28696, n28697, n28698, n28699, n28700,
         n28701, n28702, n28703, n28704, n28705, n28706, n28707, n28708,
         n28709, n28710, n28711, n28712, n28713, n28714, n28715, n28716,
         n28717, n28718, n28719, n28720, n28721, n28722, n28723, n28724,
         n28725, n28726, n28727, n28728, n28729, n28730, n28731, n28732,
         n28733, n28734, n28735, n28736, n28737, n28738, n28739, n28740,
         n28741, n28742, n28743, n28744, n28745, n28746, n28747, n28748,
         n28749, n28750, n28751, n28752, n28753, n28754, n28755, n28756,
         n28757, n28758, n28759, n28760, n28761, n28762, n28763, n28764,
         n28765, n28766, n28767, n28768, n28769, n28770, n28771, n28772,
         n28773, n28774, n28775, n28776, n28777, n28778, n28779, n28780,
         n28781, n28782, n28783, n28784, n28785, n28786, n28787, n28788,
         n28789, n28790, n28791, n28792, n28793, n28794, n28795, n28796,
         n28797, n28798, n28799, n28800, n28801, n28802, n28803, n28804,
         n28805, n28806, n28807, n28808, n28809, n28810, n28811, n28812,
         n28813, n28814, n28815, n28816, n28817, n28818, n28819, n28820,
         n28821, n28822, n28823, n28824, n28825, n28826, n28827, n28828,
         n28829, n28830, n28831, n28832, n28833, n28834, n28835, n28836,
         n28837, n28838, n28839, n28840, n28841, n28842, n28843, n28844,
         n28845, n28846, n28847, n28848, n28849, n28850, n28851, n28852,
         n28853, n28854, n28855, n28856, n28857, n28858, n28859, n28860,
         n28861, n28862, n28863, n28864, n28865, n28866, n28867, n28868,
         n28869, n28870, n28871, n28872, n28873, n28874, n28875, n28876,
         n28877, n28878, n28879, n28880, n28881, n28882, n28883, n28884,
         n28885, n28886, n28887, n28888, n28889, n28890, n28891, n28892,
         n28893, n28894, n28895, n28896, n28897, n28898, n28899, n28900,
         n28901, n28902, n28903, n28904, n28905, n28906, n28907, n28908,
         n28909, n28910, n28911, n28912, n28913, n28914, n28915, n28916,
         n28917, n28918, n28919, n28920, n28921, n28922, n28923, n28924,
         n28925, n28926, n28927, n28928, n28929, n28930, n28931, n28932,
         n28933, n28934, n28935, n28936, n28937, n28938, n28939, n28940,
         n28941, n28942, n28943, n28944, n28945, n28946, n28947, n28948,
         n28949, n28950, n28951, n28952, n28953, n28954, n28955, n28956,
         n28957, n28958, n28959, n28960, n28961, n28962, n28963, n28964,
         n28965, n28966, n28967, n28968, n28969, n28970, n28971, n28972,
         n28973, n28974, n28975, n28976, n28977, n28978, n28979, n28980,
         n28981, n28982, n28983, n28984, n28985, n28986, n28987, n28988,
         n28989, n28990, n28991, n28992, n28993, n28994, n28995, n28996,
         n28997, n28998, n28999, n29000, n29001, n29002, n29003, n29004,
         n29005, n29006, n29007, n29008, n29009, n29010, n29011, n29012,
         n29013, n29014, n29015, n29016, n29017, n29018, n29019, n29020,
         n29021, n29022, n29023, n29024, n29025, n29026, n29027, n29028,
         n29029, n29030, n29031, n29032, n29033, n29034, n29035, n29036,
         n29037, n29038, n29039, n29040, n29041, n29042, n29043, n29044,
         n29045, n29046, n29047, n29048, n29049, n29050, n29051, n29052,
         n29053, n29054, n29055, n29056, n29057, n29058, n29059, n29060,
         n29061, n29062, n29063, n29064, n29065, n29066, n29067, n29068,
         n29069, n29070, n29071, n29072, n29073, n29074, n29075, n29076,
         n29077, n29078, n29079, n29080, n29081, n29082, n29083, n29084,
         n29085, n29086, n29087, n29088, n29089, n29090, n29091, n29092,
         n29093, n29094, n29095, n29096, n29097, n29098, n29099, n29100,
         n29101, n29102, n29103, n29104, n29105, n29106, n29107, n29108,
         n29109, n29110, n29111, n29112, n29113, n29114, n29115, n29116,
         n29117, n29118, n29119, n29120, n29121, n29122, n29123, n29124,
         n29125, n29126, n29127, n29128, n29129, n29130, n29131, n29132,
         n29133, n29134, n29135, n29136, n29137, n29138, n29139, n29140,
         n29141, n29142, n29143, n29144, n29145, n29146, n29147, n29148,
         n29149, n29150, n29151, n29152, n29153, n29154, n29155, n29156,
         n29157, n29158, n29159, n29160, n29161, n29162, n29163, n29164,
         n29165, n29166, n29167, n29168, n29169, n29170, n29171, n29172,
         n29173, n29174, n29175, n29176, n29177, n29178, n29179, n29180,
         n29181, n29182, n29183, n29184, n29185, n29186, n29187, n29188,
         n29189, n29190, n29191, n29192, n29193, n29194, n29195, n29196,
         n29197, n29198, n29199, n29200, n29201, n29202, n29203, n29204,
         n29205, n29206, n29207, n29208, n29209, n29210, n29211, n29212,
         n29213, n29214, n29215, n29216, n29217, n29218, n29219, n29220,
         n29221, n29222, n29223, n29224, n29225, n29226, n29227, n29228,
         n29229, n29230, n29231, n29232, n29233, n29234, n29235, n29236,
         n29237, n29238, n29239, n29240, n29241, n29242, n29243, n29244,
         n29245, n29246, n29247, n29248, n29249, n29250, n29251, n29252,
         n29253, n29254, n29255, n29256, n29257, n29258, n29259, n29260,
         n29261, n29262, n29263, n29264, n29265, n29266, n29267, n29268,
         n29269, n29270, n29271, n29272, n29273, n29274, n29275, n29276,
         n29277, n29278, n29279, n29280, n29281, n29282, n29283, n29284,
         n29285, n29286, n29287, n29288, n29289, n29290, n29291, n29292,
         n29293, n29294, n29295, n29296, n29297, n29298, n29299, n29300,
         n29301, n29302, n29303, n29304, n29305, n29306, n29307, n29308,
         n29309, n29310, n29311, n29312, n29313, n29314, n29315, n29316,
         n29317, n29318, n29319, n29320, n29321, n29322, n29323, n29324,
         n29325, n29326, n29327, n29328, n29329, n29330, n29331, n29332,
         n29333, n29334, n29335, n29336, n29337, n29338, n29339, n29340,
         n29341, n29342, n29343, n29344, n29345, n29346, n29347, n29348,
         n29349, n29350, n29351, n29352, n29353, n29354, n29355, n29356,
         n29357, n29358, n29359, n29360, n29361, n29362, n29363, n29364,
         n29365, n29366, n29367, n29368, n29369, n29370, n29371, n29372,
         n29373, n29374, n29375, n29376, n29377, n29378, n29379, n29380,
         n29381, n29382, n29383, n29384, n29385, n29386, n29387, n29388,
         n29389, n29390, n29391, n29392, n29393, n29394, n29395, n29396,
         n29397, n29398, n29399, n29400, n29401, n29402, n29403, n29404,
         n29405, n29406, n29407, n29408, n29409, n29410, n29411, n29412,
         n29413, n29414, n29415, n29416, n29417, n29418, n29419, n29420,
         n29421, n29422, n29423, n29424, n29425, n29426, n29427, n29428,
         n29429, n29430, n29431, n29432, n29433, n29434, n29435, n29436,
         n29437, n29438, n29439, n29440, n29441, n29442, n29443, n29444,
         n29445, n29446, n29447, n29448, n29449, n29450, n29451, n29452,
         n29453, n29454, n29455, n29456, n29457, n29458, n29459, n29460,
         n29461, n29462, n29463, n29464, n29465, n29466, n29467, n29468,
         n29469, n29470, n29471, n29472, n29473, n29474, n29475, n29476,
         n29477, n29478, n29479, n29480, n29481, n29482, n29483, n29484,
         n29485, n29486, n29487, n29488, n29489, n29490, n29491, n29492,
         n29493, n29494, n29495, n29496, n29497, n29498, n29499, n29500,
         n29501, n29502, n29503, n29504, n29505, n29506, n29507, n29508,
         n29509, n29510, n29511, n29512, n29513, n29514, n29515, n29516,
         n29517, n29518, n29519, n29520, n29521, n29522, n29523, n29524,
         n29525, n29526, n29527, n29528, n29529, n29530, n29531, n29532,
         n29533, n29534, n29535, n29536, n29537, n29538, n29539, n29540,
         n29541, n29542, n29543, n29544, n29545, n29546, n29547, n29548,
         n29549, n29550, n29551, n29552, n29553, n29554, n29555, n29556,
         n29557, n29558, n29559, n29560, n29561, n29562, n29563, n29564,
         n29565, n29566, n29567, n29568, n29569, n29570, n29571, n29572,
         n29573, n29574, n29575, n29576, n29577, n29578, n29579, n29580,
         n29581, n29582, n29583, n29584, n29585, n29586, n29587, n29588,
         n29589, n29590, n29591, n29592;
  wire   [16383:0] ram;

  DFF_EN dout_reg_7_ ( .D(N29), .E(re), .CP(rclk), .Q(dout[7]) );
  DFF_EN dout_reg_6_ ( .D(N30), .E(re), .CP(rclk), .Q(dout[6]) );
  DFF_EN dout_reg_5_ ( .D(N31), .E(re), .CP(rclk), .Q(dout[5]) );
  DFF_EN dout_reg_4_ ( .D(N32), .E(re), .CP(rclk), .Q(dout[4]) );
  DFF_EN dout_reg_3_ ( .D(N33), .E(re), .CP(rclk), .Q(dout[3]) );
  DFF_EN dout_reg_2_ ( .D(N34), .E(re), .CP(rclk), .Q(dout[2]) );
  DFF_EN dout_reg_1_ ( .D(N35), .E(re), .CP(rclk), .Q(dout[1]) );
  DFF_EN dout_reg_0_ ( .D(N36), .E(re), .CP(rclk), .Q(dout[0]) );
  DFF ram_reg_40__7_ ( .D(n20304), .CP(wclk), .Q(ram[16063]) );
  DFF ram_reg_40__6_ ( .D(n20303), .CP(wclk), .Q(ram[16062]) );
  DFF ram_reg_40__5_ ( .D(n20302), .CP(wclk), .Q(ram[16061]) );
  DFF ram_reg_40__4_ ( .D(n20301), .CP(wclk), .Q(ram[16060]) );
  DFF ram_reg_40__3_ ( .D(n20300), .CP(wclk), .Q(ram[16059]) );
  DFF ram_reg_40__2_ ( .D(n20299), .CP(wclk), .Q(ram[16058]) );
  DFF ram_reg_40__1_ ( .D(n20298), .CP(wclk), .Q(ram[16057]) );
  DFF ram_reg_40__0_ ( .D(n20297), .CP(wclk), .Q(ram[16056]) );
  DFF ram_reg_56__7_ ( .D(n20176), .CP(wclk), .Q(ram[15935]) );
  DFF ram_reg_56__6_ ( .D(n20175), .CP(wclk), .Q(ram[15934]) );
  DFF ram_reg_56__5_ ( .D(n20174), .CP(wclk), .Q(ram[15933]) );
  DFF ram_reg_56__4_ ( .D(n20173), .CP(wclk), .Q(ram[15932]) );
  DFF ram_reg_56__3_ ( .D(n20172), .CP(wclk), .Q(ram[15931]) );
  DFF ram_reg_56__2_ ( .D(n20171), .CP(wclk), .Q(ram[15930]) );
  DFF ram_reg_56__1_ ( .D(n20170), .CP(wclk), .Q(ram[15929]) );
  DFF ram_reg_56__0_ ( .D(n20169), .CP(wclk), .Q(ram[15928]) );
  DFF ram_reg_136__7_ ( .D(n19536), .CP(wclk), .Q(ram[15295]) );
  DFF ram_reg_136__6_ ( .D(n19535), .CP(wclk), .Q(ram[15294]) );
  DFF ram_reg_136__5_ ( .D(n19534), .CP(wclk), .Q(ram[15293]) );
  DFF ram_reg_136__4_ ( .D(n19533), .CP(wclk), .Q(ram[15292]) );
  DFF ram_reg_136__3_ ( .D(n19532), .CP(wclk), .Q(ram[15291]) );
  DFF ram_reg_136__2_ ( .D(n19531), .CP(wclk), .Q(ram[15290]) );
  DFF ram_reg_136__1_ ( .D(n19530), .CP(wclk), .Q(ram[15289]) );
  DFF ram_reg_136__0_ ( .D(n19529), .CP(wclk), .Q(ram[15288]) );
  DFF ram_reg_140__7_ ( .D(n19504), .CP(wclk), .Q(ram[15263]) );
  DFF ram_reg_140__6_ ( .D(n19503), .CP(wclk), .Q(ram[15262]) );
  DFF ram_reg_140__5_ ( .D(n19502), .CP(wclk), .Q(ram[15261]) );
  DFF ram_reg_140__4_ ( .D(n19501), .CP(wclk), .Q(ram[15260]) );
  DFF ram_reg_140__3_ ( .D(n19500), .CP(wclk), .Q(ram[15259]) );
  DFF ram_reg_140__2_ ( .D(n19499), .CP(wclk), .Q(ram[15258]) );
  DFF ram_reg_140__1_ ( .D(n19498), .CP(wclk), .Q(ram[15257]) );
  DFF ram_reg_140__0_ ( .D(n19497), .CP(wclk), .Q(ram[15256]) );
  DFF ram_reg_152__7_ ( .D(n19408), .CP(wclk), .Q(ram[15167]) );
  DFF ram_reg_152__6_ ( .D(n19407), .CP(wclk), .Q(ram[15166]) );
  DFF ram_reg_152__5_ ( .D(n19406), .CP(wclk), .Q(ram[15165]) );
  DFF ram_reg_152__4_ ( .D(n19405), .CP(wclk), .Q(ram[15164]) );
  DFF ram_reg_152__3_ ( .D(n19404), .CP(wclk), .Q(ram[15163]) );
  DFF ram_reg_152__2_ ( .D(n19403), .CP(wclk), .Q(ram[15162]) );
  DFF ram_reg_152__1_ ( .D(n19402), .CP(wclk), .Q(ram[15161]) );
  DFF ram_reg_152__0_ ( .D(n19401), .CP(wclk), .Q(ram[15160]) );
  DFF ram_reg_160__7_ ( .D(n19344), .CP(wclk), .Q(ram[15103]) );
  DFF ram_reg_160__6_ ( .D(n19343), .CP(wclk), .Q(ram[15102]) );
  DFF ram_reg_160__5_ ( .D(n19342), .CP(wclk), .Q(ram[15101]) );
  DFF ram_reg_160__4_ ( .D(n19341), .CP(wclk), .Q(ram[15100]) );
  DFF ram_reg_160__3_ ( .D(n19340), .CP(wclk), .Q(ram[15099]) );
  DFF ram_reg_160__2_ ( .D(n19339), .CP(wclk), .Q(ram[15098]) );
  DFF ram_reg_160__1_ ( .D(n19338), .CP(wclk), .Q(ram[15097]) );
  DFF ram_reg_160__0_ ( .D(n19337), .CP(wclk), .Q(ram[15096]) );
  DFF ram_reg_168__7_ ( .D(n19280), .CP(wclk), .Q(ram[15039]) );
  DFF ram_reg_168__6_ ( .D(n19279), .CP(wclk), .Q(ram[15038]) );
  DFF ram_reg_168__5_ ( .D(n19278), .CP(wclk), .Q(ram[15037]) );
  DFF ram_reg_168__4_ ( .D(n19277), .CP(wclk), .Q(ram[15036]) );
  DFF ram_reg_168__3_ ( .D(n19276), .CP(wclk), .Q(ram[15035]) );
  DFF ram_reg_168__2_ ( .D(n19275), .CP(wclk), .Q(ram[15034]) );
  DFF ram_reg_168__1_ ( .D(n19274), .CP(wclk), .Q(ram[15033]) );
  DFF ram_reg_168__0_ ( .D(n19273), .CP(wclk), .Q(ram[15032]) );
  DFF ram_reg_172__7_ ( .D(n19248), .CP(wclk), .Q(ram[15007]) );
  DFF ram_reg_172__6_ ( .D(n19247), .CP(wclk), .Q(ram[15006]) );
  DFF ram_reg_172__5_ ( .D(n19246), .CP(wclk), .Q(ram[15005]) );
  DFF ram_reg_172__4_ ( .D(n19245), .CP(wclk), .Q(ram[15004]) );
  DFF ram_reg_172__3_ ( .D(n19244), .CP(wclk), .Q(ram[15003]) );
  DFF ram_reg_172__2_ ( .D(n19243), .CP(wclk), .Q(ram[15002]) );
  DFF ram_reg_172__1_ ( .D(n19242), .CP(wclk), .Q(ram[15001]) );
  DFF ram_reg_172__0_ ( .D(n19241), .CP(wclk), .Q(ram[15000]) );
  DFF ram_reg_176__7_ ( .D(n19216), .CP(wclk), .Q(ram[14975]) );
  DFF ram_reg_176__6_ ( .D(n19215), .CP(wclk), .Q(ram[14974]) );
  DFF ram_reg_176__5_ ( .D(n19214), .CP(wclk), .Q(ram[14973]) );
  DFF ram_reg_176__4_ ( .D(n19213), .CP(wclk), .Q(ram[14972]) );
  DFF ram_reg_176__3_ ( .D(n19212), .CP(wclk), .Q(ram[14971]) );
  DFF ram_reg_176__2_ ( .D(n19211), .CP(wclk), .Q(ram[14970]) );
  DFF ram_reg_176__1_ ( .D(n19210), .CP(wclk), .Q(ram[14969]) );
  DFF ram_reg_176__0_ ( .D(n19209), .CP(wclk), .Q(ram[14968]) );
  DFF ram_reg_184__7_ ( .D(n19152), .CP(wclk), .Q(ram[14911]) );
  DFF ram_reg_184__6_ ( .D(n19151), .CP(wclk), .Q(ram[14910]) );
  DFF ram_reg_184__5_ ( .D(n19150), .CP(wclk), .Q(ram[14909]) );
  DFF ram_reg_184__4_ ( .D(n19149), .CP(wclk), .Q(ram[14908]) );
  DFF ram_reg_184__3_ ( .D(n19148), .CP(wclk), .Q(ram[14907]) );
  DFF ram_reg_184__2_ ( .D(n19147), .CP(wclk), .Q(ram[14906]) );
  DFF ram_reg_184__1_ ( .D(n19146), .CP(wclk), .Q(ram[14905]) );
  DFF ram_reg_184__0_ ( .D(n19145), .CP(wclk), .Q(ram[14904]) );
  DFF ram_reg_188__7_ ( .D(n19120), .CP(wclk), .Q(ram[14879]) );
  DFF ram_reg_188__6_ ( .D(n19119), .CP(wclk), .Q(ram[14878]) );
  DFF ram_reg_188__5_ ( .D(n19118), .CP(wclk), .Q(ram[14877]) );
  DFF ram_reg_188__4_ ( .D(n19117), .CP(wclk), .Q(ram[14876]) );
  DFF ram_reg_188__3_ ( .D(n19116), .CP(wclk), .Q(ram[14875]) );
  DFF ram_reg_188__2_ ( .D(n19115), .CP(wclk), .Q(ram[14874]) );
  DFF ram_reg_188__1_ ( .D(n19114), .CP(wclk), .Q(ram[14873]) );
  DFF ram_reg_188__0_ ( .D(n19113), .CP(wclk), .Q(ram[14872]) );
  DFF ram_reg_200__7_ ( .D(n19024), .CP(wclk), .Q(ram[14783]) );
  DFF ram_reg_200__6_ ( .D(n19023), .CP(wclk), .Q(ram[14782]) );
  DFF ram_reg_200__5_ ( .D(n19022), .CP(wclk), .Q(ram[14781]) );
  DFF ram_reg_200__4_ ( .D(n19021), .CP(wclk), .Q(ram[14780]) );
  DFF ram_reg_200__3_ ( .D(n19020), .CP(wclk), .Q(ram[14779]) );
  DFF ram_reg_200__2_ ( .D(n19019), .CP(wclk), .Q(ram[14778]) );
  DFF ram_reg_200__1_ ( .D(n19018), .CP(wclk), .Q(ram[14777]) );
  DFF ram_reg_200__0_ ( .D(n19017), .CP(wclk), .Q(ram[14776]) );
  DFF ram_reg_232__7_ ( .D(n18768), .CP(wclk), .Q(ram[14527]) );
  DFF ram_reg_232__6_ ( .D(n18767), .CP(wclk), .Q(ram[14526]) );
  DFF ram_reg_232__5_ ( .D(n18766), .CP(wclk), .Q(ram[14525]) );
  DFF ram_reg_232__4_ ( .D(n18765), .CP(wclk), .Q(ram[14524]) );
  DFF ram_reg_232__3_ ( .D(n18764), .CP(wclk), .Q(ram[14523]) );
  DFF ram_reg_232__2_ ( .D(n18763), .CP(wclk), .Q(ram[14522]) );
  DFF ram_reg_232__1_ ( .D(n18762), .CP(wclk), .Q(ram[14521]) );
  DFF ram_reg_232__0_ ( .D(n18761), .CP(wclk), .Q(ram[14520]) );
  DFF ram_reg_236__7_ ( .D(n18736), .CP(wclk), .Q(ram[14495]) );
  DFF ram_reg_236__6_ ( .D(n18735), .CP(wclk), .Q(ram[14494]) );
  DFF ram_reg_236__5_ ( .D(n18734), .CP(wclk), .Q(ram[14493]) );
  DFF ram_reg_236__4_ ( .D(n18733), .CP(wclk), .Q(ram[14492]) );
  DFF ram_reg_236__3_ ( .D(n18732), .CP(wclk), .Q(ram[14491]) );
  DFF ram_reg_236__2_ ( .D(n18731), .CP(wclk), .Q(ram[14490]) );
  DFF ram_reg_236__1_ ( .D(n18730), .CP(wclk), .Q(ram[14489]) );
  DFF ram_reg_236__0_ ( .D(n18729), .CP(wclk), .Q(ram[14488]) );
  DFF ram_reg_248__7_ ( .D(n18640), .CP(wclk), .Q(ram[14399]) );
  DFF ram_reg_248__6_ ( .D(n18639), .CP(wclk), .Q(ram[14398]) );
  DFF ram_reg_248__5_ ( .D(n18638), .CP(wclk), .Q(ram[14397]) );
  DFF ram_reg_248__4_ ( .D(n18637), .CP(wclk), .Q(ram[14396]) );
  DFF ram_reg_248__3_ ( .D(n18636), .CP(wclk), .Q(ram[14395]) );
  DFF ram_reg_248__2_ ( .D(n18635), .CP(wclk), .Q(ram[14394]) );
  DFF ram_reg_248__1_ ( .D(n18634), .CP(wclk), .Q(ram[14393]) );
  DFF ram_reg_248__0_ ( .D(n18633), .CP(wclk), .Q(ram[14392]) );
  DFF ram_reg_252__7_ ( .D(n18608), .CP(wclk), .Q(ram[14367]) );
  DFF ram_reg_252__6_ ( .D(n18607), .CP(wclk), .Q(ram[14366]) );
  DFF ram_reg_252__5_ ( .D(n18606), .CP(wclk), .Q(ram[14365]) );
  DFF ram_reg_252__4_ ( .D(n18605), .CP(wclk), .Q(ram[14364]) );
  DFF ram_reg_252__3_ ( .D(n18604), .CP(wclk), .Q(ram[14363]) );
  DFF ram_reg_252__2_ ( .D(n18603), .CP(wclk), .Q(ram[14362]) );
  DFF ram_reg_252__1_ ( .D(n18602), .CP(wclk), .Q(ram[14361]) );
  DFF ram_reg_252__0_ ( .D(n18601), .CP(wclk), .Q(ram[14360]) );
  DFF ram_reg_296__7_ ( .D(n18256), .CP(wclk), .Q(ram[14015]) );
  DFF ram_reg_296__6_ ( .D(n18255), .CP(wclk), .Q(ram[14014]) );
  DFF ram_reg_296__5_ ( .D(n18254), .CP(wclk), .Q(ram[14013]) );
  DFF ram_reg_296__4_ ( .D(n18253), .CP(wclk), .Q(ram[14012]) );
  DFF ram_reg_296__3_ ( .D(n18252), .CP(wclk), .Q(ram[14011]) );
  DFF ram_reg_296__2_ ( .D(n18251), .CP(wclk), .Q(ram[14010]) );
  DFF ram_reg_296__1_ ( .D(n18250), .CP(wclk), .Q(ram[14009]) );
  DFF ram_reg_296__0_ ( .D(n18249), .CP(wclk), .Q(ram[14008]) );
  DFF ram_reg_312__7_ ( .D(n18128), .CP(wclk), .Q(ram[13887]) );
  DFF ram_reg_312__6_ ( .D(n18127), .CP(wclk), .Q(ram[13886]) );
  DFF ram_reg_312__5_ ( .D(n18126), .CP(wclk), .Q(ram[13885]) );
  DFF ram_reg_312__4_ ( .D(n18125), .CP(wclk), .Q(ram[13884]) );
  DFF ram_reg_312__3_ ( .D(n18124), .CP(wclk), .Q(ram[13883]) );
  DFF ram_reg_312__2_ ( .D(n18123), .CP(wclk), .Q(ram[13882]) );
  DFF ram_reg_312__1_ ( .D(n18122), .CP(wclk), .Q(ram[13881]) );
  DFF ram_reg_312__0_ ( .D(n18121), .CP(wclk), .Q(ram[13880]) );
  DFF ram_reg_316__7_ ( .D(n18096), .CP(wclk), .Q(ram[13855]) );
  DFF ram_reg_316__6_ ( .D(n18095), .CP(wclk), .Q(ram[13854]) );
  DFF ram_reg_316__5_ ( .D(n18094), .CP(wclk), .Q(ram[13853]) );
  DFF ram_reg_316__4_ ( .D(n18093), .CP(wclk), .Q(ram[13852]) );
  DFF ram_reg_316__3_ ( .D(n18092), .CP(wclk), .Q(ram[13851]) );
  DFF ram_reg_316__2_ ( .D(n18091), .CP(wclk), .Q(ram[13850]) );
  DFF ram_reg_316__1_ ( .D(n18090), .CP(wclk), .Q(ram[13849]) );
  DFF ram_reg_316__0_ ( .D(n18089), .CP(wclk), .Q(ram[13848]) );
  DFF ram_reg_392__7_ ( .D(n17488), .CP(wclk), .Q(ram[13247]) );
  DFF ram_reg_392__6_ ( .D(n17487), .CP(wclk), .Q(ram[13246]) );
  DFF ram_reg_392__5_ ( .D(n17486), .CP(wclk), .Q(ram[13245]) );
  DFF ram_reg_392__4_ ( .D(n17485), .CP(wclk), .Q(ram[13244]) );
  DFF ram_reg_392__3_ ( .D(n17484), .CP(wclk), .Q(ram[13243]) );
  DFF ram_reg_392__2_ ( .D(n17483), .CP(wclk), .Q(ram[13242]) );
  DFF ram_reg_392__1_ ( .D(n17482), .CP(wclk), .Q(ram[13241]) );
  DFF ram_reg_392__0_ ( .D(n17481), .CP(wclk), .Q(ram[13240]) );
  DFF ram_reg_396__7_ ( .D(n17456), .CP(wclk), .Q(ram[13215]) );
  DFF ram_reg_396__6_ ( .D(n17455), .CP(wclk), .Q(ram[13214]) );
  DFF ram_reg_396__5_ ( .D(n17454), .CP(wclk), .Q(ram[13213]) );
  DFF ram_reg_396__4_ ( .D(n17453), .CP(wclk), .Q(ram[13212]) );
  DFF ram_reg_396__3_ ( .D(n17452), .CP(wclk), .Q(ram[13211]) );
  DFF ram_reg_396__2_ ( .D(n17451), .CP(wclk), .Q(ram[13210]) );
  DFF ram_reg_396__1_ ( .D(n17450), .CP(wclk), .Q(ram[13209]) );
  DFF ram_reg_396__0_ ( .D(n17449), .CP(wclk), .Q(ram[13208]) );
  DFF ram_reg_408__7_ ( .D(n17360), .CP(wclk), .Q(ram[13119]) );
  DFF ram_reg_408__6_ ( .D(n17359), .CP(wclk), .Q(ram[13118]) );
  DFF ram_reg_408__5_ ( .D(n17358), .CP(wclk), .Q(ram[13117]) );
  DFF ram_reg_408__4_ ( .D(n17357), .CP(wclk), .Q(ram[13116]) );
  DFF ram_reg_408__3_ ( .D(n17356), .CP(wclk), .Q(ram[13115]) );
  DFF ram_reg_408__2_ ( .D(n17355), .CP(wclk), .Q(ram[13114]) );
  DFF ram_reg_408__1_ ( .D(n17354), .CP(wclk), .Q(ram[13113]) );
  DFF ram_reg_408__0_ ( .D(n17353), .CP(wclk), .Q(ram[13112]) );
  DFF ram_reg_412__7_ ( .D(n17328), .CP(wclk), .Q(ram[13087]) );
  DFF ram_reg_412__6_ ( .D(n17327), .CP(wclk), .Q(ram[13086]) );
  DFF ram_reg_412__5_ ( .D(n17326), .CP(wclk), .Q(ram[13085]) );
  DFF ram_reg_412__4_ ( .D(n17325), .CP(wclk), .Q(ram[13084]) );
  DFF ram_reg_412__3_ ( .D(n17324), .CP(wclk), .Q(ram[13083]) );
  DFF ram_reg_412__2_ ( .D(n17323), .CP(wclk), .Q(ram[13082]) );
  DFF ram_reg_412__1_ ( .D(n17322), .CP(wclk), .Q(ram[13081]) );
  DFF ram_reg_412__0_ ( .D(n17321), .CP(wclk), .Q(ram[13080]) );
  DFF ram_reg_416__7_ ( .D(n17296), .CP(wclk), .Q(ram[13055]) );
  DFF ram_reg_416__6_ ( .D(n17295), .CP(wclk), .Q(ram[13054]) );
  DFF ram_reg_416__5_ ( .D(n17294), .CP(wclk), .Q(ram[13053]) );
  DFF ram_reg_416__4_ ( .D(n17293), .CP(wclk), .Q(ram[13052]) );
  DFF ram_reg_416__3_ ( .D(n17292), .CP(wclk), .Q(ram[13051]) );
  DFF ram_reg_416__2_ ( .D(n17291), .CP(wclk), .Q(ram[13050]) );
  DFF ram_reg_416__1_ ( .D(n17290), .CP(wclk), .Q(ram[13049]) );
  DFF ram_reg_416__0_ ( .D(n17289), .CP(wclk), .Q(ram[13048]) );
  DFF ram_reg_424__7_ ( .D(n17232), .CP(wclk), .Q(ram[12991]) );
  DFF ram_reg_424__6_ ( .D(n17231), .CP(wclk), .Q(ram[12990]) );
  DFF ram_reg_424__5_ ( .D(n17230), .CP(wclk), .Q(ram[12989]) );
  DFF ram_reg_424__4_ ( .D(n17229), .CP(wclk), .Q(ram[12988]) );
  DFF ram_reg_424__3_ ( .D(n17228), .CP(wclk), .Q(ram[12987]) );
  DFF ram_reg_424__2_ ( .D(n17227), .CP(wclk), .Q(ram[12986]) );
  DFF ram_reg_424__1_ ( .D(n17226), .CP(wclk), .Q(ram[12985]) );
  DFF ram_reg_424__0_ ( .D(n17225), .CP(wclk), .Q(ram[12984]) );
  DFF ram_reg_428__7_ ( .D(n17200), .CP(wclk), .Q(ram[12959]) );
  DFF ram_reg_428__6_ ( .D(n17199), .CP(wclk), .Q(ram[12958]) );
  DFF ram_reg_428__5_ ( .D(n17198), .CP(wclk), .Q(ram[12957]) );
  DFF ram_reg_428__4_ ( .D(n17197), .CP(wclk), .Q(ram[12956]) );
  DFF ram_reg_428__3_ ( .D(n17196), .CP(wclk), .Q(ram[12955]) );
  DFF ram_reg_428__2_ ( .D(n17195), .CP(wclk), .Q(ram[12954]) );
  DFF ram_reg_428__1_ ( .D(n17194), .CP(wclk), .Q(ram[12953]) );
  DFF ram_reg_428__0_ ( .D(n17193), .CP(wclk), .Q(ram[12952]) );
  DFF ram_reg_432__7_ ( .D(n17168), .CP(wclk), .Q(ram[12927]) );
  DFF ram_reg_432__6_ ( .D(n17167), .CP(wclk), .Q(ram[12926]) );
  DFF ram_reg_432__5_ ( .D(n17166), .CP(wclk), .Q(ram[12925]) );
  DFF ram_reg_432__4_ ( .D(n17165), .CP(wclk), .Q(ram[12924]) );
  DFF ram_reg_432__3_ ( .D(n17164), .CP(wclk), .Q(ram[12923]) );
  DFF ram_reg_432__2_ ( .D(n17163), .CP(wclk), .Q(ram[12922]) );
  DFF ram_reg_432__1_ ( .D(n17162), .CP(wclk), .Q(ram[12921]) );
  DFF ram_reg_432__0_ ( .D(n17161), .CP(wclk), .Q(ram[12920]) );
  DFF ram_reg_440__7_ ( .D(n17104), .CP(wclk), .Q(ram[12863]) );
  DFF ram_reg_440__6_ ( .D(n17103), .CP(wclk), .Q(ram[12862]) );
  DFF ram_reg_440__5_ ( .D(n17102), .CP(wclk), .Q(ram[12861]) );
  DFF ram_reg_440__4_ ( .D(n17101), .CP(wclk), .Q(ram[12860]) );
  DFF ram_reg_440__3_ ( .D(n17100), .CP(wclk), .Q(ram[12859]) );
  DFF ram_reg_440__2_ ( .D(n17099), .CP(wclk), .Q(ram[12858]) );
  DFF ram_reg_440__1_ ( .D(n17098), .CP(wclk), .Q(ram[12857]) );
  DFF ram_reg_440__0_ ( .D(n17097), .CP(wclk), .Q(ram[12856]) );
  DFF ram_reg_444__7_ ( .D(n17072), .CP(wclk), .Q(ram[12831]) );
  DFF ram_reg_444__6_ ( .D(n17071), .CP(wclk), .Q(ram[12830]) );
  DFF ram_reg_444__5_ ( .D(n17070), .CP(wclk), .Q(ram[12829]) );
  DFF ram_reg_444__4_ ( .D(n17069), .CP(wclk), .Q(ram[12828]) );
  DFF ram_reg_444__3_ ( .D(n17068), .CP(wclk), .Q(ram[12827]) );
  DFF ram_reg_444__2_ ( .D(n17067), .CP(wclk), .Q(ram[12826]) );
  DFF ram_reg_444__1_ ( .D(n17066), .CP(wclk), .Q(ram[12825]) );
  DFF ram_reg_444__0_ ( .D(n17065), .CP(wclk), .Q(ram[12824]) );
  DFF ram_reg_456__7_ ( .D(n16976), .CP(wclk), .Q(ram[12735]) );
  DFF ram_reg_456__6_ ( .D(n16975), .CP(wclk), .Q(ram[12734]) );
  DFF ram_reg_456__5_ ( .D(n16974), .CP(wclk), .Q(ram[12733]) );
  DFF ram_reg_456__4_ ( .D(n16973), .CP(wclk), .Q(ram[12732]) );
  DFF ram_reg_456__3_ ( .D(n16972), .CP(wclk), .Q(ram[12731]) );
  DFF ram_reg_456__2_ ( .D(n16971), .CP(wclk), .Q(ram[12730]) );
  DFF ram_reg_456__1_ ( .D(n16970), .CP(wclk), .Q(ram[12729]) );
  DFF ram_reg_456__0_ ( .D(n16969), .CP(wclk), .Q(ram[12728]) );
  DFF ram_reg_460__7_ ( .D(n16944), .CP(wclk), .Q(ram[12703]) );
  DFF ram_reg_460__6_ ( .D(n16943), .CP(wclk), .Q(ram[12702]) );
  DFF ram_reg_460__5_ ( .D(n16942), .CP(wclk), .Q(ram[12701]) );
  DFF ram_reg_460__4_ ( .D(n16941), .CP(wclk), .Q(ram[12700]) );
  DFF ram_reg_460__3_ ( .D(n16940), .CP(wclk), .Q(ram[12699]) );
  DFF ram_reg_460__2_ ( .D(n16939), .CP(wclk), .Q(ram[12698]) );
  DFF ram_reg_460__1_ ( .D(n16938), .CP(wclk), .Q(ram[12697]) );
  DFF ram_reg_460__0_ ( .D(n16937), .CP(wclk), .Q(ram[12696]) );
  DFF ram_reg_472__7_ ( .D(n16848), .CP(wclk), .Q(ram[12607]) );
  DFF ram_reg_472__6_ ( .D(n16847), .CP(wclk), .Q(ram[12606]) );
  DFF ram_reg_472__5_ ( .D(n16846), .CP(wclk), .Q(ram[12605]) );
  DFF ram_reg_472__4_ ( .D(n16845), .CP(wclk), .Q(ram[12604]) );
  DFF ram_reg_472__3_ ( .D(n16844), .CP(wclk), .Q(ram[12603]) );
  DFF ram_reg_472__2_ ( .D(n16843), .CP(wclk), .Q(ram[12602]) );
  DFF ram_reg_472__1_ ( .D(n16842), .CP(wclk), .Q(ram[12601]) );
  DFF ram_reg_472__0_ ( .D(n16841), .CP(wclk), .Q(ram[12600]) );
  DFF ram_reg_488__7_ ( .D(n16720), .CP(wclk), .Q(ram[12479]) );
  DFF ram_reg_488__6_ ( .D(n16719), .CP(wclk), .Q(ram[12478]) );
  DFF ram_reg_488__5_ ( .D(n16718), .CP(wclk), .Q(ram[12477]) );
  DFF ram_reg_488__4_ ( .D(n16717), .CP(wclk), .Q(ram[12476]) );
  DFF ram_reg_488__3_ ( .D(n16716), .CP(wclk), .Q(ram[12475]) );
  DFF ram_reg_488__2_ ( .D(n16715), .CP(wclk), .Q(ram[12474]) );
  DFF ram_reg_488__1_ ( .D(n16714), .CP(wclk), .Q(ram[12473]) );
  DFF ram_reg_488__0_ ( .D(n16713), .CP(wclk), .Q(ram[12472]) );
  DFF ram_reg_492__7_ ( .D(n16688), .CP(wclk), .Q(ram[12447]) );
  DFF ram_reg_492__6_ ( .D(n16687), .CP(wclk), .Q(ram[12446]) );
  DFF ram_reg_492__5_ ( .D(n16686), .CP(wclk), .Q(ram[12445]) );
  DFF ram_reg_492__4_ ( .D(n16685), .CP(wclk), .Q(ram[12444]) );
  DFF ram_reg_492__3_ ( .D(n16684), .CP(wclk), .Q(ram[12443]) );
  DFF ram_reg_492__2_ ( .D(n16683), .CP(wclk), .Q(ram[12442]) );
  DFF ram_reg_492__1_ ( .D(n16682), .CP(wclk), .Q(ram[12441]) );
  DFF ram_reg_492__0_ ( .D(n16681), .CP(wclk), .Q(ram[12440]) );
  DFF ram_reg_496__7_ ( .D(n16656), .CP(wclk), .Q(ram[12415]) );
  DFF ram_reg_496__6_ ( .D(n16655), .CP(wclk), .Q(ram[12414]) );
  DFF ram_reg_496__5_ ( .D(n16654), .CP(wclk), .Q(ram[12413]) );
  DFF ram_reg_496__4_ ( .D(n16653), .CP(wclk), .Q(ram[12412]) );
  DFF ram_reg_496__3_ ( .D(n16652), .CP(wclk), .Q(ram[12411]) );
  DFF ram_reg_496__2_ ( .D(n16651), .CP(wclk), .Q(ram[12410]) );
  DFF ram_reg_496__1_ ( .D(n16650), .CP(wclk), .Q(ram[12409]) );
  DFF ram_reg_496__0_ ( .D(n16649), .CP(wclk), .Q(ram[12408]) );
  DFF ram_reg_504__7_ ( .D(n16592), .CP(wclk), .Q(ram[12351]) );
  DFF ram_reg_504__6_ ( .D(n16591), .CP(wclk), .Q(ram[12350]) );
  DFF ram_reg_504__5_ ( .D(n16590), .CP(wclk), .Q(ram[12349]) );
  DFF ram_reg_504__4_ ( .D(n16589), .CP(wclk), .Q(ram[12348]) );
  DFF ram_reg_504__3_ ( .D(n16588), .CP(wclk), .Q(ram[12347]) );
  DFF ram_reg_504__2_ ( .D(n16587), .CP(wclk), .Q(ram[12346]) );
  DFF ram_reg_504__1_ ( .D(n16586), .CP(wclk), .Q(ram[12345]) );
  DFF ram_reg_504__0_ ( .D(n16585), .CP(wclk), .Q(ram[12344]) );
  DFF ram_reg_508__7_ ( .D(n16560), .CP(wclk), .Q(ram[12319]) );
  DFF ram_reg_508__6_ ( .D(n16559), .CP(wclk), .Q(ram[12318]) );
  DFF ram_reg_508__5_ ( .D(n16558), .CP(wclk), .Q(ram[12317]) );
  DFF ram_reg_508__4_ ( .D(n16557), .CP(wclk), .Q(ram[12316]) );
  DFF ram_reg_508__3_ ( .D(n16556), .CP(wclk), .Q(ram[12315]) );
  DFF ram_reg_508__2_ ( .D(n16555), .CP(wclk), .Q(ram[12314]) );
  DFF ram_reg_508__1_ ( .D(n16554), .CP(wclk), .Q(ram[12313]) );
  DFF ram_reg_508__0_ ( .D(n16553), .CP(wclk), .Q(ram[12312]) );
  DFF ram_reg_520__7_ ( .D(n16464), .CP(wclk), .Q(ram[12223]) );
  DFF ram_reg_520__6_ ( .D(n16463), .CP(wclk), .Q(ram[12222]) );
  DFF ram_reg_520__5_ ( .D(n16462), .CP(wclk), .Q(ram[12221]) );
  DFF ram_reg_520__4_ ( .D(n16461), .CP(wclk), .Q(ram[12220]) );
  DFF ram_reg_520__3_ ( .D(n16460), .CP(wclk), .Q(ram[12219]) );
  DFF ram_reg_520__2_ ( .D(n16459), .CP(wclk), .Q(ram[12218]) );
  DFF ram_reg_520__1_ ( .D(n16458), .CP(wclk), .Q(ram[12217]) );
  DFF ram_reg_520__0_ ( .D(n16457), .CP(wclk), .Q(ram[12216]) );
  DFF ram_reg_536__7_ ( .D(n16336), .CP(wclk), .Q(ram[12095]) );
  DFF ram_reg_536__6_ ( .D(n16335), .CP(wclk), .Q(ram[12094]) );
  DFF ram_reg_536__5_ ( .D(n16334), .CP(wclk), .Q(ram[12093]) );
  DFF ram_reg_536__4_ ( .D(n16333), .CP(wclk), .Q(ram[12092]) );
  DFF ram_reg_536__3_ ( .D(n16332), .CP(wclk), .Q(ram[12091]) );
  DFF ram_reg_536__2_ ( .D(n16331), .CP(wclk), .Q(ram[12090]) );
  DFF ram_reg_536__1_ ( .D(n16330), .CP(wclk), .Q(ram[12089]) );
  DFF ram_reg_536__0_ ( .D(n16329), .CP(wclk), .Q(ram[12088]) );
  DFF ram_reg_552__7_ ( .D(n16208), .CP(wclk), .Q(ram[11967]) );
  DFF ram_reg_552__6_ ( .D(n16207), .CP(wclk), .Q(ram[11966]) );
  DFF ram_reg_552__5_ ( .D(n16206), .CP(wclk), .Q(ram[11965]) );
  DFF ram_reg_552__4_ ( .D(n16205), .CP(wclk), .Q(ram[11964]) );
  DFF ram_reg_552__3_ ( .D(n16204), .CP(wclk), .Q(ram[11963]) );
  DFF ram_reg_552__2_ ( .D(n16203), .CP(wclk), .Q(ram[11962]) );
  DFF ram_reg_552__1_ ( .D(n16202), .CP(wclk), .Q(ram[11961]) );
  DFF ram_reg_552__0_ ( .D(n16201), .CP(wclk), .Q(ram[11960]) );
  DFF ram_reg_556__7_ ( .D(n16176), .CP(wclk), .Q(ram[11935]) );
  DFF ram_reg_556__6_ ( .D(n16175), .CP(wclk), .Q(ram[11934]) );
  DFF ram_reg_556__5_ ( .D(n16174), .CP(wclk), .Q(ram[11933]) );
  DFF ram_reg_556__4_ ( .D(n16173), .CP(wclk), .Q(ram[11932]) );
  DFF ram_reg_556__3_ ( .D(n16172), .CP(wclk), .Q(ram[11931]) );
  DFF ram_reg_556__2_ ( .D(n16171), .CP(wclk), .Q(ram[11930]) );
  DFF ram_reg_556__1_ ( .D(n16170), .CP(wclk), .Q(ram[11929]) );
  DFF ram_reg_556__0_ ( .D(n16169), .CP(wclk), .Q(ram[11928]) );
  DFF ram_reg_568__7_ ( .D(n16080), .CP(wclk), .Q(ram[11839]) );
  DFF ram_reg_568__6_ ( .D(n16079), .CP(wclk), .Q(ram[11838]) );
  DFF ram_reg_568__5_ ( .D(n16078), .CP(wclk), .Q(ram[11837]) );
  DFF ram_reg_568__4_ ( .D(n16077), .CP(wclk), .Q(ram[11836]) );
  DFF ram_reg_568__3_ ( .D(n16076), .CP(wclk), .Q(ram[11835]) );
  DFF ram_reg_568__2_ ( .D(n16075), .CP(wclk), .Q(ram[11834]) );
  DFF ram_reg_568__1_ ( .D(n16074), .CP(wclk), .Q(ram[11833]) );
  DFF ram_reg_568__0_ ( .D(n16073), .CP(wclk), .Q(ram[11832]) );
  DFF ram_reg_572__7_ ( .D(n16048), .CP(wclk), .Q(ram[11807]) );
  DFF ram_reg_572__6_ ( .D(n16047), .CP(wclk), .Q(ram[11806]) );
  DFF ram_reg_572__5_ ( .D(n16046), .CP(wclk), .Q(ram[11805]) );
  DFF ram_reg_572__4_ ( .D(n16045), .CP(wclk), .Q(ram[11804]) );
  DFF ram_reg_572__3_ ( .D(n16044), .CP(wclk), .Q(ram[11803]) );
  DFF ram_reg_572__2_ ( .D(n16043), .CP(wclk), .Q(ram[11802]) );
  DFF ram_reg_572__1_ ( .D(n16042), .CP(wclk), .Q(ram[11801]) );
  DFF ram_reg_572__0_ ( .D(n16041), .CP(wclk), .Q(ram[11800]) );
  DFF ram_reg_632__7_ ( .D(n15568), .CP(wclk), .Q(ram[11327]) );
  DFF ram_reg_632__6_ ( .D(n15567), .CP(wclk), .Q(ram[11326]) );
  DFF ram_reg_632__5_ ( .D(n15566), .CP(wclk), .Q(ram[11325]) );
  DFF ram_reg_632__4_ ( .D(n15565), .CP(wclk), .Q(ram[11324]) );
  DFF ram_reg_632__3_ ( .D(n15564), .CP(wclk), .Q(ram[11323]) );
  DFF ram_reg_632__2_ ( .D(n15563), .CP(wclk), .Q(ram[11322]) );
  DFF ram_reg_632__1_ ( .D(n15562), .CP(wclk), .Q(ram[11321]) );
  DFF ram_reg_632__0_ ( .D(n15561), .CP(wclk), .Q(ram[11320]) );
  DFF ram_reg_640__7_ ( .D(n15504), .CP(wclk), .Q(ram[11263]) );
  DFF ram_reg_640__6_ ( .D(n15503), .CP(wclk), .Q(ram[11262]) );
  DFF ram_reg_640__5_ ( .D(n15502), .CP(wclk), .Q(ram[11261]) );
  DFF ram_reg_640__4_ ( .D(n15501), .CP(wclk), .Q(ram[11260]) );
  DFF ram_reg_640__3_ ( .D(n15500), .CP(wclk), .Q(ram[11259]) );
  DFF ram_reg_640__2_ ( .D(n15499), .CP(wclk), .Q(ram[11258]) );
  DFF ram_reg_640__1_ ( .D(n15498), .CP(wclk), .Q(ram[11257]) );
  DFF ram_reg_640__0_ ( .D(n15497), .CP(wclk), .Q(ram[11256]) );
  DFF ram_reg_648__7_ ( .D(n15440), .CP(wclk), .Q(ram[11199]) );
  DFF ram_reg_648__6_ ( .D(n15439), .CP(wclk), .Q(ram[11198]) );
  DFF ram_reg_648__5_ ( .D(n15438), .CP(wclk), .Q(ram[11197]) );
  DFF ram_reg_648__4_ ( .D(n15437), .CP(wclk), .Q(ram[11196]) );
  DFF ram_reg_648__3_ ( .D(n15436), .CP(wclk), .Q(ram[11195]) );
  DFF ram_reg_648__2_ ( .D(n15435), .CP(wclk), .Q(ram[11194]) );
  DFF ram_reg_648__1_ ( .D(n15434), .CP(wclk), .Q(ram[11193]) );
  DFF ram_reg_648__0_ ( .D(n15433), .CP(wclk), .Q(ram[11192]) );
  DFF ram_reg_652__7_ ( .D(n15408), .CP(wclk), .Q(ram[11167]) );
  DFF ram_reg_652__6_ ( .D(n15407), .CP(wclk), .Q(ram[11166]) );
  DFF ram_reg_652__5_ ( .D(n15406), .CP(wclk), .Q(ram[11165]) );
  DFF ram_reg_652__4_ ( .D(n15405), .CP(wclk), .Q(ram[11164]) );
  DFF ram_reg_652__3_ ( .D(n15404), .CP(wclk), .Q(ram[11163]) );
  DFF ram_reg_652__2_ ( .D(n15403), .CP(wclk), .Q(ram[11162]) );
  DFF ram_reg_652__1_ ( .D(n15402), .CP(wclk), .Q(ram[11161]) );
  DFF ram_reg_652__0_ ( .D(n15401), .CP(wclk), .Q(ram[11160]) );
  DFF ram_reg_656__7_ ( .D(n15376), .CP(wclk), .Q(ram[11135]) );
  DFF ram_reg_656__6_ ( .D(n15375), .CP(wclk), .Q(ram[11134]) );
  DFF ram_reg_656__5_ ( .D(n15374), .CP(wclk), .Q(ram[11133]) );
  DFF ram_reg_656__4_ ( .D(n15373), .CP(wclk), .Q(ram[11132]) );
  DFF ram_reg_656__3_ ( .D(n15372), .CP(wclk), .Q(ram[11131]) );
  DFF ram_reg_656__2_ ( .D(n15371), .CP(wclk), .Q(ram[11130]) );
  DFF ram_reg_656__1_ ( .D(n15370), .CP(wclk), .Q(ram[11129]) );
  DFF ram_reg_656__0_ ( .D(n15369), .CP(wclk), .Q(ram[11128]) );
  DFF ram_reg_664__7_ ( .D(n15312), .CP(wclk), .Q(ram[11071]) );
  DFF ram_reg_664__6_ ( .D(n15311), .CP(wclk), .Q(ram[11070]) );
  DFF ram_reg_664__5_ ( .D(n15310), .CP(wclk), .Q(ram[11069]) );
  DFF ram_reg_664__4_ ( .D(n15309), .CP(wclk), .Q(ram[11068]) );
  DFF ram_reg_664__3_ ( .D(n15308), .CP(wclk), .Q(ram[11067]) );
  DFF ram_reg_664__2_ ( .D(n15307), .CP(wclk), .Q(ram[11066]) );
  DFF ram_reg_664__1_ ( .D(n15306), .CP(wclk), .Q(ram[11065]) );
  DFF ram_reg_664__0_ ( .D(n15305), .CP(wclk), .Q(ram[11064]) );
  DFF ram_reg_668__7_ ( .D(n15280), .CP(wclk), .Q(ram[11039]) );
  DFF ram_reg_668__6_ ( .D(n15279), .CP(wclk), .Q(ram[11038]) );
  DFF ram_reg_668__5_ ( .D(n15278), .CP(wclk), .Q(ram[11037]) );
  DFF ram_reg_668__4_ ( .D(n15277), .CP(wclk), .Q(ram[11036]) );
  DFF ram_reg_668__3_ ( .D(n15276), .CP(wclk), .Q(ram[11035]) );
  DFF ram_reg_668__2_ ( .D(n15275), .CP(wclk), .Q(ram[11034]) );
  DFF ram_reg_668__1_ ( .D(n15274), .CP(wclk), .Q(ram[11033]) );
  DFF ram_reg_668__0_ ( .D(n15273), .CP(wclk), .Q(ram[11032]) );
  DFF ram_reg_672__7_ ( .D(n15248), .CP(wclk), .Q(ram[11007]) );
  DFF ram_reg_672__6_ ( .D(n15247), .CP(wclk), .Q(ram[11006]) );
  DFF ram_reg_672__5_ ( .D(n15246), .CP(wclk), .Q(ram[11005]) );
  DFF ram_reg_672__4_ ( .D(n15245), .CP(wclk), .Q(ram[11004]) );
  DFF ram_reg_672__3_ ( .D(n15244), .CP(wclk), .Q(ram[11003]) );
  DFF ram_reg_672__2_ ( .D(n15243), .CP(wclk), .Q(ram[11002]) );
  DFF ram_reg_672__1_ ( .D(n15242), .CP(wclk), .Q(ram[11001]) );
  DFF ram_reg_672__0_ ( .D(n15241), .CP(wclk), .Q(ram[11000]) );
  DFF ram_reg_680__7_ ( .D(n15184), .CP(wclk), .Q(ram[10943]) );
  DFF ram_reg_680__6_ ( .D(n15183), .CP(wclk), .Q(ram[10942]) );
  DFF ram_reg_680__5_ ( .D(n15182), .CP(wclk), .Q(ram[10941]) );
  DFF ram_reg_680__4_ ( .D(n15181), .CP(wclk), .Q(ram[10940]) );
  DFF ram_reg_680__3_ ( .D(n15180), .CP(wclk), .Q(ram[10939]) );
  DFF ram_reg_680__2_ ( .D(n15179), .CP(wclk), .Q(ram[10938]) );
  DFF ram_reg_680__1_ ( .D(n15178), .CP(wclk), .Q(ram[10937]) );
  DFF ram_reg_680__0_ ( .D(n15177), .CP(wclk), .Q(ram[10936]) );
  DFF ram_reg_684__7_ ( .D(n15152), .CP(wclk), .Q(ram[10911]) );
  DFF ram_reg_684__6_ ( .D(n15151), .CP(wclk), .Q(ram[10910]) );
  DFF ram_reg_684__5_ ( .D(n15150), .CP(wclk), .Q(ram[10909]) );
  DFF ram_reg_684__4_ ( .D(n15149), .CP(wclk), .Q(ram[10908]) );
  DFF ram_reg_684__3_ ( .D(n15148), .CP(wclk), .Q(ram[10907]) );
  DFF ram_reg_684__2_ ( .D(n15147), .CP(wclk), .Q(ram[10906]) );
  DFF ram_reg_684__1_ ( .D(n15146), .CP(wclk), .Q(ram[10905]) );
  DFF ram_reg_684__0_ ( .D(n15145), .CP(wclk), .Q(ram[10904]) );
  DFF ram_reg_688__7_ ( .D(n15120), .CP(wclk), .Q(ram[10879]) );
  DFF ram_reg_688__6_ ( .D(n15119), .CP(wclk), .Q(ram[10878]) );
  DFF ram_reg_688__5_ ( .D(n15118), .CP(wclk), .Q(ram[10877]) );
  DFF ram_reg_688__4_ ( .D(n15117), .CP(wclk), .Q(ram[10876]) );
  DFF ram_reg_688__3_ ( .D(n15116), .CP(wclk), .Q(ram[10875]) );
  DFF ram_reg_688__2_ ( .D(n15115), .CP(wclk), .Q(ram[10874]) );
  DFF ram_reg_688__1_ ( .D(n15114), .CP(wclk), .Q(ram[10873]) );
  DFF ram_reg_688__0_ ( .D(n15113), .CP(wclk), .Q(ram[10872]) );
  DFF ram_reg_692__7_ ( .D(n15088), .CP(wclk), .Q(ram[10847]) );
  DFF ram_reg_692__6_ ( .D(n15087), .CP(wclk), .Q(ram[10846]) );
  DFF ram_reg_692__5_ ( .D(n15086), .CP(wclk), .Q(ram[10845]) );
  DFF ram_reg_692__4_ ( .D(n15085), .CP(wclk), .Q(ram[10844]) );
  DFF ram_reg_692__3_ ( .D(n15084), .CP(wclk), .Q(ram[10843]) );
  DFF ram_reg_692__2_ ( .D(n15083), .CP(wclk), .Q(ram[10842]) );
  DFF ram_reg_692__1_ ( .D(n15082), .CP(wclk), .Q(ram[10841]) );
  DFF ram_reg_692__0_ ( .D(n15081), .CP(wclk), .Q(ram[10840]) );
  DFF ram_reg_696__7_ ( .D(n15056), .CP(wclk), .Q(ram[10815]) );
  DFF ram_reg_696__6_ ( .D(n15055), .CP(wclk), .Q(ram[10814]) );
  DFF ram_reg_696__5_ ( .D(n15054), .CP(wclk), .Q(ram[10813]) );
  DFF ram_reg_696__4_ ( .D(n15053), .CP(wclk), .Q(ram[10812]) );
  DFF ram_reg_696__3_ ( .D(n15052), .CP(wclk), .Q(ram[10811]) );
  DFF ram_reg_696__2_ ( .D(n15051), .CP(wclk), .Q(ram[10810]) );
  DFF ram_reg_696__1_ ( .D(n15050), .CP(wclk), .Q(ram[10809]) );
  DFF ram_reg_696__0_ ( .D(n15049), .CP(wclk), .Q(ram[10808]) );
  DFF ram_reg_700__7_ ( .D(n15024), .CP(wclk), .Q(ram[10783]) );
  DFF ram_reg_700__6_ ( .D(n15023), .CP(wclk), .Q(ram[10782]) );
  DFF ram_reg_700__5_ ( .D(n15022), .CP(wclk), .Q(ram[10781]) );
  DFF ram_reg_700__4_ ( .D(n15021), .CP(wclk), .Q(ram[10780]) );
  DFF ram_reg_700__3_ ( .D(n15020), .CP(wclk), .Q(ram[10779]) );
  DFF ram_reg_700__2_ ( .D(n15019), .CP(wclk), .Q(ram[10778]) );
  DFF ram_reg_700__1_ ( .D(n15018), .CP(wclk), .Q(ram[10777]) );
  DFF ram_reg_700__0_ ( .D(n15017), .CP(wclk), .Q(ram[10776]) );
  DFF ram_reg_712__7_ ( .D(n14928), .CP(wclk), .Q(ram[10687]) );
  DFF ram_reg_712__6_ ( .D(n14927), .CP(wclk), .Q(ram[10686]) );
  DFF ram_reg_712__5_ ( .D(n14926), .CP(wclk), .Q(ram[10685]) );
  DFF ram_reg_712__4_ ( .D(n14925), .CP(wclk), .Q(ram[10684]) );
  DFF ram_reg_712__3_ ( .D(n14924), .CP(wclk), .Q(ram[10683]) );
  DFF ram_reg_712__2_ ( .D(n14923), .CP(wclk), .Q(ram[10682]) );
  DFF ram_reg_712__1_ ( .D(n14922), .CP(wclk), .Q(ram[10681]) );
  DFF ram_reg_712__0_ ( .D(n14921), .CP(wclk), .Q(ram[10680]) );
  DFF ram_reg_716__7_ ( .D(n14896), .CP(wclk), .Q(ram[10655]) );
  DFF ram_reg_716__6_ ( .D(n14895), .CP(wclk), .Q(ram[10654]) );
  DFF ram_reg_716__5_ ( .D(n14894), .CP(wclk), .Q(ram[10653]) );
  DFF ram_reg_716__4_ ( .D(n14893), .CP(wclk), .Q(ram[10652]) );
  DFF ram_reg_716__3_ ( .D(n14892), .CP(wclk), .Q(ram[10651]) );
  DFF ram_reg_716__2_ ( .D(n14891), .CP(wclk), .Q(ram[10650]) );
  DFF ram_reg_716__1_ ( .D(n14890), .CP(wclk), .Q(ram[10649]) );
  DFF ram_reg_716__0_ ( .D(n14889), .CP(wclk), .Q(ram[10648]) );
  DFF ram_reg_728__7_ ( .D(n14800), .CP(wclk), .Q(ram[10559]) );
  DFF ram_reg_728__6_ ( .D(n14799), .CP(wclk), .Q(ram[10558]) );
  DFF ram_reg_728__5_ ( .D(n14798), .CP(wclk), .Q(ram[10557]) );
  DFF ram_reg_728__4_ ( .D(n14797), .CP(wclk), .Q(ram[10556]) );
  DFF ram_reg_728__3_ ( .D(n14796), .CP(wclk), .Q(ram[10555]) );
  DFF ram_reg_728__2_ ( .D(n14795), .CP(wclk), .Q(ram[10554]) );
  DFF ram_reg_728__1_ ( .D(n14794), .CP(wclk), .Q(ram[10553]) );
  DFF ram_reg_728__0_ ( .D(n14793), .CP(wclk), .Q(ram[10552]) );
  DFF ram_reg_732__7_ ( .D(n14768), .CP(wclk), .Q(ram[10527]) );
  DFF ram_reg_732__6_ ( .D(n14767), .CP(wclk), .Q(ram[10526]) );
  DFF ram_reg_732__5_ ( .D(n14766), .CP(wclk), .Q(ram[10525]) );
  DFF ram_reg_732__4_ ( .D(n14765), .CP(wclk), .Q(ram[10524]) );
  DFF ram_reg_732__3_ ( .D(n14764), .CP(wclk), .Q(ram[10523]) );
  DFF ram_reg_732__2_ ( .D(n14763), .CP(wclk), .Q(ram[10522]) );
  DFF ram_reg_732__1_ ( .D(n14762), .CP(wclk), .Q(ram[10521]) );
  DFF ram_reg_732__0_ ( .D(n14761), .CP(wclk), .Q(ram[10520]) );
  DFF ram_reg_736__7_ ( .D(n14736), .CP(wclk), .Q(ram[10495]) );
  DFF ram_reg_736__6_ ( .D(n14735), .CP(wclk), .Q(ram[10494]) );
  DFF ram_reg_736__5_ ( .D(n14734), .CP(wclk), .Q(ram[10493]) );
  DFF ram_reg_736__4_ ( .D(n14733), .CP(wclk), .Q(ram[10492]) );
  DFF ram_reg_736__3_ ( .D(n14732), .CP(wclk), .Q(ram[10491]) );
  DFF ram_reg_736__2_ ( .D(n14731), .CP(wclk), .Q(ram[10490]) );
  DFF ram_reg_736__1_ ( .D(n14730), .CP(wclk), .Q(ram[10489]) );
  DFF ram_reg_736__0_ ( .D(n14729), .CP(wclk), .Q(ram[10488]) );
  DFF ram_reg_744__7_ ( .D(n14672), .CP(wclk), .Q(ram[10431]) );
  DFF ram_reg_744__6_ ( .D(n14671), .CP(wclk), .Q(ram[10430]) );
  DFF ram_reg_744__5_ ( .D(n14670), .CP(wclk), .Q(ram[10429]) );
  DFF ram_reg_744__4_ ( .D(n14669), .CP(wclk), .Q(ram[10428]) );
  DFF ram_reg_744__3_ ( .D(n14668), .CP(wclk), .Q(ram[10427]) );
  DFF ram_reg_744__2_ ( .D(n14667), .CP(wclk), .Q(ram[10426]) );
  DFF ram_reg_744__1_ ( .D(n14666), .CP(wclk), .Q(ram[10425]) );
  DFF ram_reg_744__0_ ( .D(n14665), .CP(wclk), .Q(ram[10424]) );
  DFF ram_reg_748__7_ ( .D(n14640), .CP(wclk), .Q(ram[10399]) );
  DFF ram_reg_748__6_ ( .D(n14639), .CP(wclk), .Q(ram[10398]) );
  DFF ram_reg_748__5_ ( .D(n14638), .CP(wclk), .Q(ram[10397]) );
  DFF ram_reg_748__4_ ( .D(n14637), .CP(wclk), .Q(ram[10396]) );
  DFF ram_reg_748__3_ ( .D(n14636), .CP(wclk), .Q(ram[10395]) );
  DFF ram_reg_748__2_ ( .D(n14635), .CP(wclk), .Q(ram[10394]) );
  DFF ram_reg_748__1_ ( .D(n14634), .CP(wclk), .Q(ram[10393]) );
  DFF ram_reg_748__0_ ( .D(n14633), .CP(wclk), .Q(ram[10392]) );
  DFF ram_reg_752__7_ ( .D(n14608), .CP(wclk), .Q(ram[10367]) );
  DFF ram_reg_752__6_ ( .D(n14607), .CP(wclk), .Q(ram[10366]) );
  DFF ram_reg_752__5_ ( .D(n14606), .CP(wclk), .Q(ram[10365]) );
  DFF ram_reg_752__4_ ( .D(n14605), .CP(wclk), .Q(ram[10364]) );
  DFF ram_reg_752__3_ ( .D(n14604), .CP(wclk), .Q(ram[10363]) );
  DFF ram_reg_752__2_ ( .D(n14603), .CP(wclk), .Q(ram[10362]) );
  DFF ram_reg_752__1_ ( .D(n14602), .CP(wclk), .Q(ram[10361]) );
  DFF ram_reg_752__0_ ( .D(n14601), .CP(wclk), .Q(ram[10360]) );
  DFF ram_reg_760__7_ ( .D(n14544), .CP(wclk), .Q(ram[10303]) );
  DFF ram_reg_760__6_ ( .D(n14543), .CP(wclk), .Q(ram[10302]) );
  DFF ram_reg_760__5_ ( .D(n14542), .CP(wclk), .Q(ram[10301]) );
  DFF ram_reg_760__4_ ( .D(n14541), .CP(wclk), .Q(ram[10300]) );
  DFF ram_reg_760__3_ ( .D(n14540), .CP(wclk), .Q(ram[10299]) );
  DFF ram_reg_760__2_ ( .D(n14539), .CP(wclk), .Q(ram[10298]) );
  DFF ram_reg_760__1_ ( .D(n14538), .CP(wclk), .Q(ram[10297]) );
  DFF ram_reg_760__0_ ( .D(n14537), .CP(wclk), .Q(ram[10296]) );
  DFF ram_reg_764__7_ ( .D(n14512), .CP(wclk), .Q(ram[10271]) );
  DFF ram_reg_764__6_ ( .D(n14511), .CP(wclk), .Q(ram[10270]) );
  DFF ram_reg_764__5_ ( .D(n14510), .CP(wclk), .Q(ram[10269]) );
  DFF ram_reg_764__4_ ( .D(n14509), .CP(wclk), .Q(ram[10268]) );
  DFF ram_reg_764__3_ ( .D(n14508), .CP(wclk), .Q(ram[10267]) );
  DFF ram_reg_764__2_ ( .D(n14507), .CP(wclk), .Q(ram[10266]) );
  DFF ram_reg_764__1_ ( .D(n14506), .CP(wclk), .Q(ram[10265]) );
  DFF ram_reg_764__0_ ( .D(n14505), .CP(wclk), .Q(ram[10264]) );
  DFF ram_reg_776__7_ ( .D(n14416), .CP(wclk), .Q(ram[10175]) );
  DFF ram_reg_776__6_ ( .D(n14415), .CP(wclk), .Q(ram[10174]) );
  DFF ram_reg_776__5_ ( .D(n14414), .CP(wclk), .Q(ram[10173]) );
  DFF ram_reg_776__4_ ( .D(n14413), .CP(wclk), .Q(ram[10172]) );
  DFF ram_reg_776__3_ ( .D(n14412), .CP(wclk), .Q(ram[10171]) );
  DFF ram_reg_776__2_ ( .D(n14411), .CP(wclk), .Q(ram[10170]) );
  DFF ram_reg_776__1_ ( .D(n14410), .CP(wclk), .Q(ram[10169]) );
  DFF ram_reg_776__0_ ( .D(n14409), .CP(wclk), .Q(ram[10168]) );
  DFF ram_reg_780__7_ ( .D(n14384), .CP(wclk), .Q(ram[10143]) );
  DFF ram_reg_780__6_ ( .D(n14383), .CP(wclk), .Q(ram[10142]) );
  DFF ram_reg_780__5_ ( .D(n14382), .CP(wclk), .Q(ram[10141]) );
  DFF ram_reg_780__4_ ( .D(n14381), .CP(wclk), .Q(ram[10140]) );
  DFF ram_reg_780__3_ ( .D(n14380), .CP(wclk), .Q(ram[10139]) );
  DFF ram_reg_780__2_ ( .D(n14379), .CP(wclk), .Q(ram[10138]) );
  DFF ram_reg_780__1_ ( .D(n14378), .CP(wclk), .Q(ram[10137]) );
  DFF ram_reg_780__0_ ( .D(n14377), .CP(wclk), .Q(ram[10136]) );
  DFF ram_reg_792__7_ ( .D(n14288), .CP(wclk), .Q(ram[10047]) );
  DFF ram_reg_792__6_ ( .D(n14287), .CP(wclk), .Q(ram[10046]) );
  DFF ram_reg_792__5_ ( .D(n14286), .CP(wclk), .Q(ram[10045]) );
  DFF ram_reg_792__4_ ( .D(n14285), .CP(wclk), .Q(ram[10044]) );
  DFF ram_reg_792__3_ ( .D(n14284), .CP(wclk), .Q(ram[10043]) );
  DFF ram_reg_792__2_ ( .D(n14283), .CP(wclk), .Q(ram[10042]) );
  DFF ram_reg_792__1_ ( .D(n14282), .CP(wclk), .Q(ram[10041]) );
  DFF ram_reg_792__0_ ( .D(n14281), .CP(wclk), .Q(ram[10040]) );
  DFF ram_reg_808__7_ ( .D(n14160), .CP(wclk), .Q(ram[9919]) );
  DFF ram_reg_808__6_ ( .D(n14159), .CP(wclk), .Q(ram[9918]) );
  DFF ram_reg_808__5_ ( .D(n14158), .CP(wclk), .Q(ram[9917]) );
  DFF ram_reg_808__4_ ( .D(n14157), .CP(wclk), .Q(ram[9916]) );
  DFF ram_reg_808__3_ ( .D(n14156), .CP(wclk), .Q(ram[9915]) );
  DFF ram_reg_808__2_ ( .D(n14155), .CP(wclk), .Q(ram[9914]) );
  DFF ram_reg_808__1_ ( .D(n14154), .CP(wclk), .Q(ram[9913]) );
  DFF ram_reg_808__0_ ( .D(n14153), .CP(wclk), .Q(ram[9912]) );
  DFF ram_reg_812__7_ ( .D(n14128), .CP(wclk), .Q(ram[9887]) );
  DFF ram_reg_812__6_ ( .D(n14127), .CP(wclk), .Q(ram[9886]) );
  DFF ram_reg_812__5_ ( .D(n14126), .CP(wclk), .Q(ram[9885]) );
  DFF ram_reg_812__4_ ( .D(n14125), .CP(wclk), .Q(ram[9884]) );
  DFF ram_reg_812__3_ ( .D(n14124), .CP(wclk), .Q(ram[9883]) );
  DFF ram_reg_812__2_ ( .D(n14123), .CP(wclk), .Q(ram[9882]) );
  DFF ram_reg_812__1_ ( .D(n14122), .CP(wclk), .Q(ram[9881]) );
  DFF ram_reg_812__0_ ( .D(n14121), .CP(wclk), .Q(ram[9880]) );
  DFF ram_reg_816__7_ ( .D(n14096), .CP(wclk), .Q(ram[9855]) );
  DFF ram_reg_816__6_ ( .D(n14095), .CP(wclk), .Q(ram[9854]) );
  DFF ram_reg_816__5_ ( .D(n14094), .CP(wclk), .Q(ram[9853]) );
  DFF ram_reg_816__4_ ( .D(n14093), .CP(wclk), .Q(ram[9852]) );
  DFF ram_reg_816__3_ ( .D(n14092), .CP(wclk), .Q(ram[9851]) );
  DFF ram_reg_816__2_ ( .D(n14091), .CP(wclk), .Q(ram[9850]) );
  DFF ram_reg_816__1_ ( .D(n14090), .CP(wclk), .Q(ram[9849]) );
  DFF ram_reg_816__0_ ( .D(n14089), .CP(wclk), .Q(ram[9848]) );
  DFF ram_reg_824__7_ ( .D(n14032), .CP(wclk), .Q(ram[9791]) );
  DFF ram_reg_824__6_ ( .D(n14031), .CP(wclk), .Q(ram[9790]) );
  DFF ram_reg_824__5_ ( .D(n14030), .CP(wclk), .Q(ram[9789]) );
  DFF ram_reg_824__4_ ( .D(n14029), .CP(wclk), .Q(ram[9788]) );
  DFF ram_reg_824__3_ ( .D(n14028), .CP(wclk), .Q(ram[9787]) );
  DFF ram_reg_824__2_ ( .D(n14027), .CP(wclk), .Q(ram[9786]) );
  DFF ram_reg_824__1_ ( .D(n14026), .CP(wclk), .Q(ram[9785]) );
  DFF ram_reg_824__0_ ( .D(n14025), .CP(wclk), .Q(ram[9784]) );
  DFF ram_reg_828__7_ ( .D(n14000), .CP(wclk), .Q(ram[9759]) );
  DFF ram_reg_828__6_ ( .D(n13999), .CP(wclk), .Q(ram[9758]) );
  DFF ram_reg_828__5_ ( .D(n13998), .CP(wclk), .Q(ram[9757]) );
  DFF ram_reg_828__4_ ( .D(n13997), .CP(wclk), .Q(ram[9756]) );
  DFF ram_reg_828__3_ ( .D(n13996), .CP(wclk), .Q(ram[9755]) );
  DFF ram_reg_828__2_ ( .D(n13995), .CP(wclk), .Q(ram[9754]) );
  DFF ram_reg_828__1_ ( .D(n13994), .CP(wclk), .Q(ram[9753]) );
  DFF ram_reg_828__0_ ( .D(n13993), .CP(wclk), .Q(ram[9752]) );
  DFF ram_reg_872__7_ ( .D(n13648), .CP(wclk), .Q(ram[9407]) );
  DFF ram_reg_872__6_ ( .D(n13647), .CP(wclk), .Q(ram[9406]) );
  DFF ram_reg_872__5_ ( .D(n13646), .CP(wclk), .Q(ram[9405]) );
  DFF ram_reg_872__4_ ( .D(n13645), .CP(wclk), .Q(ram[9404]) );
  DFF ram_reg_872__3_ ( .D(n13644), .CP(wclk), .Q(ram[9403]) );
  DFF ram_reg_872__2_ ( .D(n13643), .CP(wclk), .Q(ram[9402]) );
  DFF ram_reg_872__1_ ( .D(n13642), .CP(wclk), .Q(ram[9401]) );
  DFF ram_reg_872__0_ ( .D(n13641), .CP(wclk), .Q(ram[9400]) );
  DFF ram_reg_888__7_ ( .D(n13520), .CP(wclk), .Q(ram[9279]) );
  DFF ram_reg_888__6_ ( .D(n13519), .CP(wclk), .Q(ram[9278]) );
  DFF ram_reg_888__5_ ( .D(n13518), .CP(wclk), .Q(ram[9277]) );
  DFF ram_reg_888__4_ ( .D(n13517), .CP(wclk), .Q(ram[9276]) );
  DFF ram_reg_888__3_ ( .D(n13516), .CP(wclk), .Q(ram[9275]) );
  DFF ram_reg_888__2_ ( .D(n13515), .CP(wclk), .Q(ram[9274]) );
  DFF ram_reg_888__1_ ( .D(n13514), .CP(wclk), .Q(ram[9273]) );
  DFF ram_reg_888__0_ ( .D(n13513), .CP(wclk), .Q(ram[9272]) );
  DFF ram_reg_896__7_ ( .D(n13456), .CP(wclk), .Q(ram[9215]) );
  DFF ram_reg_896__6_ ( .D(n13455), .CP(wclk), .Q(ram[9214]) );
  DFF ram_reg_896__5_ ( .D(n13454), .CP(wclk), .Q(ram[9213]) );
  DFF ram_reg_896__4_ ( .D(n13453), .CP(wclk), .Q(ram[9212]) );
  DFF ram_reg_896__3_ ( .D(n13452), .CP(wclk), .Q(ram[9211]) );
  DFF ram_reg_896__2_ ( .D(n13451), .CP(wclk), .Q(ram[9210]) );
  DFF ram_reg_896__1_ ( .D(n13450), .CP(wclk), .Q(ram[9209]) );
  DFF ram_reg_896__0_ ( .D(n13449), .CP(wclk), .Q(ram[9208]) );
  DFF ram_reg_904__7_ ( .D(n13392), .CP(wclk), .Q(ram[9151]) );
  DFF ram_reg_904__6_ ( .D(n13391), .CP(wclk), .Q(ram[9150]) );
  DFF ram_reg_904__5_ ( .D(n13390), .CP(wclk), .Q(ram[9149]) );
  DFF ram_reg_904__4_ ( .D(n13389), .CP(wclk), .Q(ram[9148]) );
  DFF ram_reg_904__3_ ( .D(n13388), .CP(wclk), .Q(ram[9147]) );
  DFF ram_reg_904__2_ ( .D(n13387), .CP(wclk), .Q(ram[9146]) );
  DFF ram_reg_904__1_ ( .D(n13386), .CP(wclk), .Q(ram[9145]) );
  DFF ram_reg_904__0_ ( .D(n13385), .CP(wclk), .Q(ram[9144]) );
  DFF ram_reg_908__7_ ( .D(n13360), .CP(wclk), .Q(ram[9119]) );
  DFF ram_reg_908__6_ ( .D(n13359), .CP(wclk), .Q(ram[9118]) );
  DFF ram_reg_908__5_ ( .D(n13358), .CP(wclk), .Q(ram[9117]) );
  DFF ram_reg_908__4_ ( .D(n13357), .CP(wclk), .Q(ram[9116]) );
  DFF ram_reg_908__3_ ( .D(n13356), .CP(wclk), .Q(ram[9115]) );
  DFF ram_reg_908__2_ ( .D(n13355), .CP(wclk), .Q(ram[9114]) );
  DFF ram_reg_908__1_ ( .D(n13354), .CP(wclk), .Q(ram[9113]) );
  DFF ram_reg_908__0_ ( .D(n13353), .CP(wclk), .Q(ram[9112]) );
  DFF ram_reg_912__7_ ( .D(n13328), .CP(wclk), .Q(ram[9087]) );
  DFF ram_reg_912__6_ ( .D(n13327), .CP(wclk), .Q(ram[9086]) );
  DFF ram_reg_912__5_ ( .D(n13326), .CP(wclk), .Q(ram[9085]) );
  DFF ram_reg_912__4_ ( .D(n13325), .CP(wclk), .Q(ram[9084]) );
  DFF ram_reg_912__3_ ( .D(n13324), .CP(wclk), .Q(ram[9083]) );
  DFF ram_reg_912__2_ ( .D(n13323), .CP(wclk), .Q(ram[9082]) );
  DFF ram_reg_912__1_ ( .D(n13322), .CP(wclk), .Q(ram[9081]) );
  DFF ram_reg_912__0_ ( .D(n13321), .CP(wclk), .Q(ram[9080]) );
  DFF ram_reg_920__7_ ( .D(n13264), .CP(wclk), .Q(ram[9023]) );
  DFF ram_reg_920__6_ ( .D(n13263), .CP(wclk), .Q(ram[9022]) );
  DFF ram_reg_920__5_ ( .D(n13262), .CP(wclk), .Q(ram[9021]) );
  DFF ram_reg_920__4_ ( .D(n13261), .CP(wclk), .Q(ram[9020]) );
  DFF ram_reg_920__3_ ( .D(n13260), .CP(wclk), .Q(ram[9019]) );
  DFF ram_reg_920__2_ ( .D(n13259), .CP(wclk), .Q(ram[9018]) );
  DFF ram_reg_920__1_ ( .D(n13258), .CP(wclk), .Q(ram[9017]) );
  DFF ram_reg_920__0_ ( .D(n13257), .CP(wclk), .Q(ram[9016]) );
  DFF ram_reg_924__7_ ( .D(n13232), .CP(wclk), .Q(ram[8991]) );
  DFF ram_reg_924__6_ ( .D(n13231), .CP(wclk), .Q(ram[8990]) );
  DFF ram_reg_924__5_ ( .D(n13230), .CP(wclk), .Q(ram[8989]) );
  DFF ram_reg_924__4_ ( .D(n13229), .CP(wclk), .Q(ram[8988]) );
  DFF ram_reg_924__3_ ( .D(n13228), .CP(wclk), .Q(ram[8987]) );
  DFF ram_reg_924__2_ ( .D(n13227), .CP(wclk), .Q(ram[8986]) );
  DFF ram_reg_924__1_ ( .D(n13226), .CP(wclk), .Q(ram[8985]) );
  DFF ram_reg_924__0_ ( .D(n13225), .CP(wclk), .Q(ram[8984]) );
  DFF ram_reg_928__7_ ( .D(n13200), .CP(wclk), .Q(ram[8959]) );
  DFF ram_reg_928__6_ ( .D(n13199), .CP(wclk), .Q(ram[8958]) );
  DFF ram_reg_928__5_ ( .D(n13198), .CP(wclk), .Q(ram[8957]) );
  DFF ram_reg_928__4_ ( .D(n13197), .CP(wclk), .Q(ram[8956]) );
  DFF ram_reg_928__3_ ( .D(n13196), .CP(wclk), .Q(ram[8955]) );
  DFF ram_reg_928__2_ ( .D(n13195), .CP(wclk), .Q(ram[8954]) );
  DFF ram_reg_928__1_ ( .D(n13194), .CP(wclk), .Q(ram[8953]) );
  DFF ram_reg_928__0_ ( .D(n13193), .CP(wclk), .Q(ram[8952]) );
  DFF ram_reg_932__7_ ( .D(n13168), .CP(wclk), .Q(ram[8927]) );
  DFF ram_reg_932__6_ ( .D(n13167), .CP(wclk), .Q(ram[8926]) );
  DFF ram_reg_932__5_ ( .D(n13166), .CP(wclk), .Q(ram[8925]) );
  DFF ram_reg_932__4_ ( .D(n13165), .CP(wclk), .Q(ram[8924]) );
  DFF ram_reg_932__3_ ( .D(n13164), .CP(wclk), .Q(ram[8923]) );
  DFF ram_reg_932__2_ ( .D(n13163), .CP(wclk), .Q(ram[8922]) );
  DFF ram_reg_932__1_ ( .D(n13162), .CP(wclk), .Q(ram[8921]) );
  DFF ram_reg_932__0_ ( .D(n13161), .CP(wclk), .Q(ram[8920]) );
  DFF ram_reg_936__7_ ( .D(n13136), .CP(wclk), .Q(ram[8895]) );
  DFF ram_reg_936__6_ ( .D(n13135), .CP(wclk), .Q(ram[8894]) );
  DFF ram_reg_936__5_ ( .D(n13134), .CP(wclk), .Q(ram[8893]) );
  DFF ram_reg_936__4_ ( .D(n13133), .CP(wclk), .Q(ram[8892]) );
  DFF ram_reg_936__3_ ( .D(n13132), .CP(wclk), .Q(ram[8891]) );
  DFF ram_reg_936__2_ ( .D(n13131), .CP(wclk), .Q(ram[8890]) );
  DFF ram_reg_936__1_ ( .D(n13130), .CP(wclk), .Q(ram[8889]) );
  DFF ram_reg_936__0_ ( .D(n13129), .CP(wclk), .Q(ram[8888]) );
  DFF ram_reg_940__7_ ( .D(n13104), .CP(wclk), .Q(ram[8863]) );
  DFF ram_reg_940__6_ ( .D(n13103), .CP(wclk), .Q(ram[8862]) );
  DFF ram_reg_940__5_ ( .D(n13102), .CP(wclk), .Q(ram[8861]) );
  DFF ram_reg_940__4_ ( .D(n13101), .CP(wclk), .Q(ram[8860]) );
  DFF ram_reg_940__3_ ( .D(n13100), .CP(wclk), .Q(ram[8859]) );
  DFF ram_reg_940__2_ ( .D(n13099), .CP(wclk), .Q(ram[8858]) );
  DFF ram_reg_940__1_ ( .D(n13098), .CP(wclk), .Q(ram[8857]) );
  DFF ram_reg_940__0_ ( .D(n13097), .CP(wclk), .Q(ram[8856]) );
  DFF ram_reg_944__7_ ( .D(n13072), .CP(wclk), .Q(ram[8831]) );
  DFF ram_reg_944__6_ ( .D(n13071), .CP(wclk), .Q(ram[8830]) );
  DFF ram_reg_944__5_ ( .D(n13070), .CP(wclk), .Q(ram[8829]) );
  DFF ram_reg_944__4_ ( .D(n13069), .CP(wclk), .Q(ram[8828]) );
  DFF ram_reg_944__3_ ( .D(n13068), .CP(wclk), .Q(ram[8827]) );
  DFF ram_reg_944__2_ ( .D(n13067), .CP(wclk), .Q(ram[8826]) );
  DFF ram_reg_944__1_ ( .D(n13066), .CP(wclk), .Q(ram[8825]) );
  DFF ram_reg_944__0_ ( .D(n13065), .CP(wclk), .Q(ram[8824]) );
  DFF ram_reg_948__7_ ( .D(n13040), .CP(wclk), .Q(ram[8799]) );
  DFF ram_reg_948__6_ ( .D(n13039), .CP(wclk), .Q(ram[8798]) );
  DFF ram_reg_948__5_ ( .D(n13038), .CP(wclk), .Q(ram[8797]) );
  DFF ram_reg_948__4_ ( .D(n13037), .CP(wclk), .Q(ram[8796]) );
  DFF ram_reg_948__3_ ( .D(n13036), .CP(wclk), .Q(ram[8795]) );
  DFF ram_reg_948__2_ ( .D(n13035), .CP(wclk), .Q(ram[8794]) );
  DFF ram_reg_948__1_ ( .D(n13034), .CP(wclk), .Q(ram[8793]) );
  DFF ram_reg_948__0_ ( .D(n13033), .CP(wclk), .Q(ram[8792]) );
  DFF ram_reg_952__7_ ( .D(n13008), .CP(wclk), .Q(ram[8767]) );
  DFF ram_reg_952__6_ ( .D(n13007), .CP(wclk), .Q(ram[8766]) );
  DFF ram_reg_952__5_ ( .D(n13006), .CP(wclk), .Q(ram[8765]) );
  DFF ram_reg_952__4_ ( .D(n13005), .CP(wclk), .Q(ram[8764]) );
  DFF ram_reg_952__3_ ( .D(n13004), .CP(wclk), .Q(ram[8763]) );
  DFF ram_reg_952__2_ ( .D(n13003), .CP(wclk), .Q(ram[8762]) );
  DFF ram_reg_952__1_ ( .D(n13002), .CP(wclk), .Q(ram[8761]) );
  DFF ram_reg_952__0_ ( .D(n13001), .CP(wclk), .Q(ram[8760]) );
  DFF ram_reg_956__7_ ( .D(n12976), .CP(wclk), .Q(ram[8735]) );
  DFF ram_reg_956__6_ ( .D(n12975), .CP(wclk), .Q(ram[8734]) );
  DFF ram_reg_956__5_ ( .D(n12974), .CP(wclk), .Q(ram[8733]) );
  DFF ram_reg_956__4_ ( .D(n12973), .CP(wclk), .Q(ram[8732]) );
  DFF ram_reg_956__3_ ( .D(n12972), .CP(wclk), .Q(ram[8731]) );
  DFF ram_reg_956__2_ ( .D(n12971), .CP(wclk), .Q(ram[8730]) );
  DFF ram_reg_956__1_ ( .D(n12970), .CP(wclk), .Q(ram[8729]) );
  DFF ram_reg_956__0_ ( .D(n12969), .CP(wclk), .Q(ram[8728]) );
  DFF ram_reg_960__7_ ( .D(n12944), .CP(wclk), .Q(ram[8703]) );
  DFF ram_reg_960__6_ ( .D(n12943), .CP(wclk), .Q(ram[8702]) );
  DFF ram_reg_960__5_ ( .D(n12942), .CP(wclk), .Q(ram[8701]) );
  DFF ram_reg_960__4_ ( .D(n12941), .CP(wclk), .Q(ram[8700]) );
  DFF ram_reg_960__3_ ( .D(n12940), .CP(wclk), .Q(ram[8699]) );
  DFF ram_reg_960__2_ ( .D(n12939), .CP(wclk), .Q(ram[8698]) );
  DFF ram_reg_960__1_ ( .D(n12938), .CP(wclk), .Q(ram[8697]) );
  DFF ram_reg_960__0_ ( .D(n12937), .CP(wclk), .Q(ram[8696]) );
  DFF ram_reg_968__7_ ( .D(n12880), .CP(wclk), .Q(ram[8639]) );
  DFF ram_reg_968__6_ ( .D(n12879), .CP(wclk), .Q(ram[8638]) );
  DFF ram_reg_968__5_ ( .D(n12878), .CP(wclk), .Q(ram[8637]) );
  DFF ram_reg_968__4_ ( .D(n12877), .CP(wclk), .Q(ram[8636]) );
  DFF ram_reg_968__3_ ( .D(n12876), .CP(wclk), .Q(ram[8635]) );
  DFF ram_reg_968__2_ ( .D(n12875), .CP(wclk), .Q(ram[8634]) );
  DFF ram_reg_968__1_ ( .D(n12874), .CP(wclk), .Q(ram[8633]) );
  DFF ram_reg_968__0_ ( .D(n12873), .CP(wclk), .Q(ram[8632]) );
  DFF ram_reg_972__7_ ( .D(n12848), .CP(wclk), .Q(ram[8607]) );
  DFF ram_reg_972__6_ ( .D(n12847), .CP(wclk), .Q(ram[8606]) );
  DFF ram_reg_972__5_ ( .D(n12846), .CP(wclk), .Q(ram[8605]) );
  DFF ram_reg_972__4_ ( .D(n12845), .CP(wclk), .Q(ram[8604]) );
  DFF ram_reg_972__3_ ( .D(n12844), .CP(wclk), .Q(ram[8603]) );
  DFF ram_reg_972__2_ ( .D(n12843), .CP(wclk), .Q(ram[8602]) );
  DFF ram_reg_972__1_ ( .D(n12842), .CP(wclk), .Q(ram[8601]) );
  DFF ram_reg_972__0_ ( .D(n12841), .CP(wclk), .Q(ram[8600]) );
  DFF ram_reg_984__7_ ( .D(n12752), .CP(wclk), .Q(ram[8511]) );
  DFF ram_reg_984__6_ ( .D(n12751), .CP(wclk), .Q(ram[8510]) );
  DFF ram_reg_984__5_ ( .D(n12750), .CP(wclk), .Q(ram[8509]) );
  DFF ram_reg_984__4_ ( .D(n12749), .CP(wclk), .Q(ram[8508]) );
  DFF ram_reg_984__3_ ( .D(n12748), .CP(wclk), .Q(ram[8507]) );
  DFF ram_reg_984__2_ ( .D(n12747), .CP(wclk), .Q(ram[8506]) );
  DFF ram_reg_984__1_ ( .D(n12746), .CP(wclk), .Q(ram[8505]) );
  DFF ram_reg_984__0_ ( .D(n12745), .CP(wclk), .Q(ram[8504]) );
  DFF ram_reg_988__7_ ( .D(n12720), .CP(wclk), .Q(ram[8479]) );
  DFF ram_reg_988__6_ ( .D(n12719), .CP(wclk), .Q(ram[8478]) );
  DFF ram_reg_988__5_ ( .D(n12718), .CP(wclk), .Q(ram[8477]) );
  DFF ram_reg_988__4_ ( .D(n12717), .CP(wclk), .Q(ram[8476]) );
  DFF ram_reg_988__3_ ( .D(n12716), .CP(wclk), .Q(ram[8475]) );
  DFF ram_reg_988__2_ ( .D(n12715), .CP(wclk), .Q(ram[8474]) );
  DFF ram_reg_988__1_ ( .D(n12714), .CP(wclk), .Q(ram[8473]) );
  DFF ram_reg_988__0_ ( .D(n12713), .CP(wclk), .Q(ram[8472]) );
  DFF ram_reg_992__7_ ( .D(n12688), .CP(wclk), .Q(ram[8447]) );
  DFF ram_reg_992__6_ ( .D(n12687), .CP(wclk), .Q(ram[8446]) );
  DFF ram_reg_992__5_ ( .D(n12686), .CP(wclk), .Q(ram[8445]) );
  DFF ram_reg_992__4_ ( .D(n12685), .CP(wclk), .Q(ram[8444]) );
  DFF ram_reg_992__3_ ( .D(n12684), .CP(wclk), .Q(ram[8443]) );
  DFF ram_reg_992__2_ ( .D(n12683), .CP(wclk), .Q(ram[8442]) );
  DFF ram_reg_992__1_ ( .D(n12682), .CP(wclk), .Q(ram[8441]) );
  DFF ram_reg_992__0_ ( .D(n12681), .CP(wclk), .Q(ram[8440]) );
  DFF ram_reg_1000__7_ ( .D(n12624), .CP(wclk), .Q(ram[8383]) );
  DFF ram_reg_1000__6_ ( .D(n12623), .CP(wclk), .Q(ram[8382]) );
  DFF ram_reg_1000__5_ ( .D(n12622), .CP(wclk), .Q(ram[8381]) );
  DFF ram_reg_1000__4_ ( .D(n12621), .CP(wclk), .Q(ram[8380]) );
  DFF ram_reg_1000__3_ ( .D(n12620), .CP(wclk), .Q(ram[8379]) );
  DFF ram_reg_1000__2_ ( .D(n12619), .CP(wclk), .Q(ram[8378]) );
  DFF ram_reg_1000__1_ ( .D(n12618), .CP(wclk), .Q(ram[8377]) );
  DFF ram_reg_1000__0_ ( .D(n12617), .CP(wclk), .Q(ram[8376]) );
  DFF ram_reg_1004__7_ ( .D(n12592), .CP(wclk), .Q(ram[8351]) );
  DFF ram_reg_1004__6_ ( .D(n12591), .CP(wclk), .Q(ram[8350]) );
  DFF ram_reg_1004__5_ ( .D(n12590), .CP(wclk), .Q(ram[8349]) );
  DFF ram_reg_1004__4_ ( .D(n12589), .CP(wclk), .Q(ram[8348]) );
  DFF ram_reg_1004__3_ ( .D(n12588), .CP(wclk), .Q(ram[8347]) );
  DFF ram_reg_1004__2_ ( .D(n12587), .CP(wclk), .Q(ram[8346]) );
  DFF ram_reg_1004__1_ ( .D(n12586), .CP(wclk), .Q(ram[8345]) );
  DFF ram_reg_1004__0_ ( .D(n12585), .CP(wclk), .Q(ram[8344]) );
  DFF ram_reg_1008__7_ ( .D(n12560), .CP(wclk), .Q(ram[8319]) );
  DFF ram_reg_1008__6_ ( .D(n12559), .CP(wclk), .Q(ram[8318]) );
  DFF ram_reg_1008__5_ ( .D(n12558), .CP(wclk), .Q(ram[8317]) );
  DFF ram_reg_1008__4_ ( .D(n12557), .CP(wclk), .Q(ram[8316]) );
  DFF ram_reg_1008__3_ ( .D(n12556), .CP(wclk), .Q(ram[8315]) );
  DFF ram_reg_1008__2_ ( .D(n12555), .CP(wclk), .Q(ram[8314]) );
  DFF ram_reg_1008__1_ ( .D(n12554), .CP(wclk), .Q(ram[8313]) );
  DFF ram_reg_1008__0_ ( .D(n12553), .CP(wclk), .Q(ram[8312]) );
  DFF ram_reg_1016__7_ ( .D(n12496), .CP(wclk), .Q(ram[8255]) );
  DFF ram_reg_1016__6_ ( .D(n12495), .CP(wclk), .Q(ram[8254]) );
  DFF ram_reg_1016__5_ ( .D(n12494), .CP(wclk), .Q(ram[8253]) );
  DFF ram_reg_1016__4_ ( .D(n12493), .CP(wclk), .Q(ram[8252]) );
  DFF ram_reg_1016__3_ ( .D(n12492), .CP(wclk), .Q(ram[8251]) );
  DFF ram_reg_1016__2_ ( .D(n12491), .CP(wclk), .Q(ram[8250]) );
  DFF ram_reg_1016__1_ ( .D(n12490), .CP(wclk), .Q(ram[8249]) );
  DFF ram_reg_1016__0_ ( .D(n12489), .CP(wclk), .Q(ram[8248]) );
  DFF ram_reg_1020__7_ ( .D(n12464), .CP(wclk), .Q(ram[8223]) );
  DFF ram_reg_1020__6_ ( .D(n12463), .CP(wclk), .Q(ram[8222]) );
  DFF ram_reg_1020__5_ ( .D(n12462), .CP(wclk), .Q(ram[8221]) );
  DFF ram_reg_1020__4_ ( .D(n12461), .CP(wclk), .Q(ram[8220]) );
  DFF ram_reg_1020__3_ ( .D(n12460), .CP(wclk), .Q(ram[8219]) );
  DFF ram_reg_1020__2_ ( .D(n12459), .CP(wclk), .Q(ram[8218]) );
  DFF ram_reg_1020__1_ ( .D(n12458), .CP(wclk), .Q(ram[8217]) );
  DFF ram_reg_1020__0_ ( .D(n12457), .CP(wclk), .Q(ram[8216]) );
  DFF ram_reg_1032__7_ ( .D(n12368), .CP(wclk), .Q(ram[8127]) );
  DFF ram_reg_1032__6_ ( .D(n12367), .CP(wclk), .Q(ram[8126]) );
  DFF ram_reg_1032__5_ ( .D(n12366), .CP(wclk), .Q(ram[8125]) );
  DFF ram_reg_1032__4_ ( .D(n12365), .CP(wclk), .Q(ram[8124]) );
  DFF ram_reg_1032__3_ ( .D(n12364), .CP(wclk), .Q(ram[8123]) );
  DFF ram_reg_1032__2_ ( .D(n12363), .CP(wclk), .Q(ram[8122]) );
  DFF ram_reg_1032__1_ ( .D(n12362), .CP(wclk), .Q(ram[8121]) );
  DFF ram_reg_1032__0_ ( .D(n12361), .CP(wclk), .Q(ram[8120]) );
  DFF ram_reg_1064__7_ ( .D(n12112), .CP(wclk), .Q(ram[7871]) );
  DFF ram_reg_1064__6_ ( .D(n12111), .CP(wclk), .Q(ram[7870]) );
  DFF ram_reg_1064__5_ ( .D(n12110), .CP(wclk), .Q(ram[7869]) );
  DFF ram_reg_1064__4_ ( .D(n12109), .CP(wclk), .Q(ram[7868]) );
  DFF ram_reg_1064__3_ ( .D(n12108), .CP(wclk), .Q(ram[7867]) );
  DFF ram_reg_1064__2_ ( .D(n12107), .CP(wclk), .Q(ram[7866]) );
  DFF ram_reg_1064__1_ ( .D(n12106), .CP(wclk), .Q(ram[7865]) );
  DFF ram_reg_1064__0_ ( .D(n12105), .CP(wclk), .Q(ram[7864]) );
  DFF ram_reg_1068__7_ ( .D(n12080), .CP(wclk), .Q(ram[7839]) );
  DFF ram_reg_1068__6_ ( .D(n12079), .CP(wclk), .Q(ram[7838]) );
  DFF ram_reg_1068__5_ ( .D(n12078), .CP(wclk), .Q(ram[7837]) );
  DFF ram_reg_1068__4_ ( .D(n12077), .CP(wclk), .Q(ram[7836]) );
  DFF ram_reg_1068__3_ ( .D(n12076), .CP(wclk), .Q(ram[7835]) );
  DFF ram_reg_1068__2_ ( .D(n12075), .CP(wclk), .Q(ram[7834]) );
  DFF ram_reg_1068__1_ ( .D(n12074), .CP(wclk), .Q(ram[7833]) );
  DFF ram_reg_1068__0_ ( .D(n12073), .CP(wclk), .Q(ram[7832]) );
  DFF ram_reg_1080__7_ ( .D(n11984), .CP(wclk), .Q(ram[7743]) );
  DFF ram_reg_1080__6_ ( .D(n11983), .CP(wclk), .Q(ram[7742]) );
  DFF ram_reg_1080__5_ ( .D(n11982), .CP(wclk), .Q(ram[7741]) );
  DFF ram_reg_1080__4_ ( .D(n11981), .CP(wclk), .Q(ram[7740]) );
  DFF ram_reg_1080__3_ ( .D(n11980), .CP(wclk), .Q(ram[7739]) );
  DFF ram_reg_1080__2_ ( .D(n11979), .CP(wclk), .Q(ram[7738]) );
  DFF ram_reg_1080__1_ ( .D(n11978), .CP(wclk), .Q(ram[7737]) );
  DFF ram_reg_1080__0_ ( .D(n11977), .CP(wclk), .Q(ram[7736]) );
  DFF ram_reg_1084__7_ ( .D(n11952), .CP(wclk), .Q(ram[7711]) );
  DFF ram_reg_1084__6_ ( .D(n11951), .CP(wclk), .Q(ram[7710]) );
  DFF ram_reg_1084__5_ ( .D(n11950), .CP(wclk), .Q(ram[7709]) );
  DFF ram_reg_1084__4_ ( .D(n11949), .CP(wclk), .Q(ram[7708]) );
  DFF ram_reg_1084__3_ ( .D(n11948), .CP(wclk), .Q(ram[7707]) );
  DFF ram_reg_1084__2_ ( .D(n11947), .CP(wclk), .Q(ram[7706]) );
  DFF ram_reg_1084__1_ ( .D(n11946), .CP(wclk), .Q(ram[7705]) );
  DFF ram_reg_1084__0_ ( .D(n11945), .CP(wclk), .Q(ram[7704]) );
  DFF ram_reg_1152__7_ ( .D(n11408), .CP(wclk), .Q(ram[7167]) );
  DFF ram_reg_1152__6_ ( .D(n11407), .CP(wclk), .Q(ram[7166]) );
  DFF ram_reg_1152__5_ ( .D(n11406), .CP(wclk), .Q(ram[7165]) );
  DFF ram_reg_1152__4_ ( .D(n11405), .CP(wclk), .Q(ram[7164]) );
  DFF ram_reg_1152__3_ ( .D(n11404), .CP(wclk), .Q(ram[7163]) );
  DFF ram_reg_1152__2_ ( .D(n11403), .CP(wclk), .Q(ram[7162]) );
  DFF ram_reg_1152__1_ ( .D(n11402), .CP(wclk), .Q(ram[7161]) );
  DFF ram_reg_1152__0_ ( .D(n11401), .CP(wclk), .Q(ram[7160]) );
  DFF ram_reg_1160__7_ ( .D(n11344), .CP(wclk), .Q(ram[7103]) );
  DFF ram_reg_1160__6_ ( .D(n11343), .CP(wclk), .Q(ram[7102]) );
  DFF ram_reg_1160__5_ ( .D(n11342), .CP(wclk), .Q(ram[7101]) );
  DFF ram_reg_1160__4_ ( .D(n11341), .CP(wclk), .Q(ram[7100]) );
  DFF ram_reg_1160__3_ ( .D(n11340), .CP(wclk), .Q(ram[7099]) );
  DFF ram_reg_1160__2_ ( .D(n11339), .CP(wclk), .Q(ram[7098]) );
  DFF ram_reg_1160__1_ ( .D(n11338), .CP(wclk), .Q(ram[7097]) );
  DFF ram_reg_1160__0_ ( .D(n11337), .CP(wclk), .Q(ram[7096]) );
  DFF ram_reg_1164__7_ ( .D(n11312), .CP(wclk), .Q(ram[7071]) );
  DFF ram_reg_1164__6_ ( .D(n11311), .CP(wclk), .Q(ram[7070]) );
  DFF ram_reg_1164__5_ ( .D(n11310), .CP(wclk), .Q(ram[7069]) );
  DFF ram_reg_1164__4_ ( .D(n11309), .CP(wclk), .Q(ram[7068]) );
  DFF ram_reg_1164__3_ ( .D(n11308), .CP(wclk), .Q(ram[7067]) );
  DFF ram_reg_1164__2_ ( .D(n11307), .CP(wclk), .Q(ram[7066]) );
  DFF ram_reg_1164__1_ ( .D(n11306), .CP(wclk), .Q(ram[7065]) );
  DFF ram_reg_1164__0_ ( .D(n11305), .CP(wclk), .Q(ram[7064]) );
  DFF ram_reg_1176__7_ ( .D(n11216), .CP(wclk), .Q(ram[6975]) );
  DFF ram_reg_1176__6_ ( .D(n11215), .CP(wclk), .Q(ram[6974]) );
  DFF ram_reg_1176__5_ ( .D(n11214), .CP(wclk), .Q(ram[6973]) );
  DFF ram_reg_1176__4_ ( .D(n11213), .CP(wclk), .Q(ram[6972]) );
  DFF ram_reg_1176__3_ ( .D(n11212), .CP(wclk), .Q(ram[6971]) );
  DFF ram_reg_1176__2_ ( .D(n11211), .CP(wclk), .Q(ram[6970]) );
  DFF ram_reg_1176__1_ ( .D(n11210), .CP(wclk), .Q(ram[6969]) );
  DFF ram_reg_1176__0_ ( .D(n11209), .CP(wclk), .Q(ram[6968]) );
  DFF ram_reg_1180__7_ ( .D(n11184), .CP(wclk), .Q(ram[6943]) );
  DFF ram_reg_1180__6_ ( .D(n11183), .CP(wclk), .Q(ram[6942]) );
  DFF ram_reg_1180__5_ ( .D(n11182), .CP(wclk), .Q(ram[6941]) );
  DFF ram_reg_1180__4_ ( .D(n11181), .CP(wclk), .Q(ram[6940]) );
  DFF ram_reg_1180__3_ ( .D(n11180), .CP(wclk), .Q(ram[6939]) );
  DFF ram_reg_1180__2_ ( .D(n11179), .CP(wclk), .Q(ram[6938]) );
  DFF ram_reg_1180__1_ ( .D(n11178), .CP(wclk), .Q(ram[6937]) );
  DFF ram_reg_1180__0_ ( .D(n11177), .CP(wclk), .Q(ram[6936]) );
  DFF ram_reg_1184__7_ ( .D(n11152), .CP(wclk), .Q(ram[6911]) );
  DFF ram_reg_1184__6_ ( .D(n11151), .CP(wclk), .Q(ram[6910]) );
  DFF ram_reg_1184__5_ ( .D(n11150), .CP(wclk), .Q(ram[6909]) );
  DFF ram_reg_1184__4_ ( .D(n11149), .CP(wclk), .Q(ram[6908]) );
  DFF ram_reg_1184__3_ ( .D(n11148), .CP(wclk), .Q(ram[6907]) );
  DFF ram_reg_1184__2_ ( .D(n11147), .CP(wclk), .Q(ram[6906]) );
  DFF ram_reg_1184__1_ ( .D(n11146), .CP(wclk), .Q(ram[6905]) );
  DFF ram_reg_1184__0_ ( .D(n11145), .CP(wclk), .Q(ram[6904]) );
  DFF ram_reg_1192__7_ ( .D(n11088), .CP(wclk), .Q(ram[6847]) );
  DFF ram_reg_1192__6_ ( .D(n11087), .CP(wclk), .Q(ram[6846]) );
  DFF ram_reg_1192__5_ ( .D(n11086), .CP(wclk), .Q(ram[6845]) );
  DFF ram_reg_1192__4_ ( .D(n11085), .CP(wclk), .Q(ram[6844]) );
  DFF ram_reg_1192__3_ ( .D(n11084), .CP(wclk), .Q(ram[6843]) );
  DFF ram_reg_1192__2_ ( .D(n11083), .CP(wclk), .Q(ram[6842]) );
  DFF ram_reg_1192__1_ ( .D(n11082), .CP(wclk), .Q(ram[6841]) );
  DFF ram_reg_1192__0_ ( .D(n11081), .CP(wclk), .Q(ram[6840]) );
  DFF ram_reg_1196__7_ ( .D(n11056), .CP(wclk), .Q(ram[6815]) );
  DFF ram_reg_1196__6_ ( .D(n11055), .CP(wclk), .Q(ram[6814]) );
  DFF ram_reg_1196__5_ ( .D(n11054), .CP(wclk), .Q(ram[6813]) );
  DFF ram_reg_1196__4_ ( .D(n11053), .CP(wclk), .Q(ram[6812]) );
  DFF ram_reg_1196__3_ ( .D(n11052), .CP(wclk), .Q(ram[6811]) );
  DFF ram_reg_1196__2_ ( .D(n11051), .CP(wclk), .Q(ram[6810]) );
  DFF ram_reg_1196__1_ ( .D(n11050), .CP(wclk), .Q(ram[6809]) );
  DFF ram_reg_1196__0_ ( .D(n11049), .CP(wclk), .Q(ram[6808]) );
  DFF ram_reg_1200__7_ ( .D(n11024), .CP(wclk), .Q(ram[6783]) );
  DFF ram_reg_1200__6_ ( .D(n11023), .CP(wclk), .Q(ram[6782]) );
  DFF ram_reg_1200__5_ ( .D(n11022), .CP(wclk), .Q(ram[6781]) );
  DFF ram_reg_1200__4_ ( .D(n11021), .CP(wclk), .Q(ram[6780]) );
  DFF ram_reg_1200__3_ ( .D(n11020), .CP(wclk), .Q(ram[6779]) );
  DFF ram_reg_1200__2_ ( .D(n11019), .CP(wclk), .Q(ram[6778]) );
  DFF ram_reg_1200__1_ ( .D(n11018), .CP(wclk), .Q(ram[6777]) );
  DFF ram_reg_1200__0_ ( .D(n11017), .CP(wclk), .Q(ram[6776]) );
  DFF ram_reg_1208__7_ ( .D(n10960), .CP(wclk), .Q(ram[6719]) );
  DFF ram_reg_1208__6_ ( .D(n10959), .CP(wclk), .Q(ram[6718]) );
  DFF ram_reg_1208__5_ ( .D(n10958), .CP(wclk), .Q(ram[6717]) );
  DFF ram_reg_1208__4_ ( .D(n10957), .CP(wclk), .Q(ram[6716]) );
  DFF ram_reg_1208__3_ ( .D(n10956), .CP(wclk), .Q(ram[6715]) );
  DFF ram_reg_1208__2_ ( .D(n10955), .CP(wclk), .Q(ram[6714]) );
  DFF ram_reg_1208__1_ ( .D(n10954), .CP(wclk), .Q(ram[6713]) );
  DFF ram_reg_1208__0_ ( .D(n10953), .CP(wclk), .Q(ram[6712]) );
  DFF ram_reg_1212__7_ ( .D(n10928), .CP(wclk), .Q(ram[6687]) );
  DFF ram_reg_1212__6_ ( .D(n10927), .CP(wclk), .Q(ram[6686]) );
  DFF ram_reg_1212__5_ ( .D(n10926), .CP(wclk), .Q(ram[6685]) );
  DFF ram_reg_1212__4_ ( .D(n10925), .CP(wclk), .Q(ram[6684]) );
  DFF ram_reg_1212__3_ ( .D(n10924), .CP(wclk), .Q(ram[6683]) );
  DFF ram_reg_1212__2_ ( .D(n10923), .CP(wclk), .Q(ram[6682]) );
  DFF ram_reg_1212__1_ ( .D(n10922), .CP(wclk), .Q(ram[6681]) );
  DFF ram_reg_1212__0_ ( .D(n10921), .CP(wclk), .Q(ram[6680]) );
  DFF ram_reg_1224__7_ ( .D(n10832), .CP(wclk), .Q(ram[6591]) );
  DFF ram_reg_1224__6_ ( .D(n10831), .CP(wclk), .Q(ram[6590]) );
  DFF ram_reg_1224__5_ ( .D(n10830), .CP(wclk), .Q(ram[6589]) );
  DFF ram_reg_1224__4_ ( .D(n10829), .CP(wclk), .Q(ram[6588]) );
  DFF ram_reg_1224__3_ ( .D(n10828), .CP(wclk), .Q(ram[6587]) );
  DFF ram_reg_1224__2_ ( .D(n10827), .CP(wclk), .Q(ram[6586]) );
  DFF ram_reg_1224__1_ ( .D(n10826), .CP(wclk), .Q(ram[6585]) );
  DFF ram_reg_1224__0_ ( .D(n10825), .CP(wclk), .Q(ram[6584]) );
  DFF ram_reg_1228__7_ ( .D(n10800), .CP(wclk), .Q(ram[6559]) );
  DFF ram_reg_1228__6_ ( .D(n10799), .CP(wclk), .Q(ram[6558]) );
  DFF ram_reg_1228__5_ ( .D(n10798), .CP(wclk), .Q(ram[6557]) );
  DFF ram_reg_1228__4_ ( .D(n10797), .CP(wclk), .Q(ram[6556]) );
  DFF ram_reg_1228__3_ ( .D(n10796), .CP(wclk), .Q(ram[6555]) );
  DFF ram_reg_1228__2_ ( .D(n10795), .CP(wclk), .Q(ram[6554]) );
  DFF ram_reg_1228__1_ ( .D(n10794), .CP(wclk), .Q(ram[6553]) );
  DFF ram_reg_1228__0_ ( .D(n10793), .CP(wclk), .Q(ram[6552]) );
  DFF ram_reg_1240__7_ ( .D(n10704), .CP(wclk), .Q(ram[6463]) );
  DFF ram_reg_1240__6_ ( .D(n10703), .CP(wclk), .Q(ram[6462]) );
  DFF ram_reg_1240__5_ ( .D(n10702), .CP(wclk), .Q(ram[6461]) );
  DFF ram_reg_1240__4_ ( .D(n10701), .CP(wclk), .Q(ram[6460]) );
  DFF ram_reg_1240__3_ ( .D(n10700), .CP(wclk), .Q(ram[6459]) );
  DFF ram_reg_1240__2_ ( .D(n10699), .CP(wclk), .Q(ram[6458]) );
  DFF ram_reg_1240__1_ ( .D(n10698), .CP(wclk), .Q(ram[6457]) );
  DFF ram_reg_1240__0_ ( .D(n10697), .CP(wclk), .Q(ram[6456]) );
  DFF ram_reg_1248__7_ ( .D(n10640), .CP(wclk), .Q(ram[6399]) );
  DFF ram_reg_1248__6_ ( .D(n10639), .CP(wclk), .Q(ram[6398]) );
  DFF ram_reg_1248__5_ ( .D(n10638), .CP(wclk), .Q(ram[6397]) );
  DFF ram_reg_1248__4_ ( .D(n10637), .CP(wclk), .Q(ram[6396]) );
  DFF ram_reg_1248__3_ ( .D(n10636), .CP(wclk), .Q(ram[6395]) );
  DFF ram_reg_1248__2_ ( .D(n10635), .CP(wclk), .Q(ram[6394]) );
  DFF ram_reg_1248__1_ ( .D(n10634), .CP(wclk), .Q(ram[6393]) );
  DFF ram_reg_1248__0_ ( .D(n10633), .CP(wclk), .Q(ram[6392]) );
  DFF ram_reg_1256__7_ ( .D(n10576), .CP(wclk), .Q(ram[6335]) );
  DFF ram_reg_1256__6_ ( .D(n10575), .CP(wclk), .Q(ram[6334]) );
  DFF ram_reg_1256__5_ ( .D(n10574), .CP(wclk), .Q(ram[6333]) );
  DFF ram_reg_1256__4_ ( .D(n10573), .CP(wclk), .Q(ram[6332]) );
  DFF ram_reg_1256__3_ ( .D(n10572), .CP(wclk), .Q(ram[6331]) );
  DFF ram_reg_1256__2_ ( .D(n10571), .CP(wclk), .Q(ram[6330]) );
  DFF ram_reg_1256__1_ ( .D(n10570), .CP(wclk), .Q(ram[6329]) );
  DFF ram_reg_1256__0_ ( .D(n10569), .CP(wclk), .Q(ram[6328]) );
  DFF ram_reg_1260__7_ ( .D(n10544), .CP(wclk), .Q(ram[6303]) );
  DFF ram_reg_1260__6_ ( .D(n10543), .CP(wclk), .Q(ram[6302]) );
  DFF ram_reg_1260__5_ ( .D(n10542), .CP(wclk), .Q(ram[6301]) );
  DFF ram_reg_1260__4_ ( .D(n10541), .CP(wclk), .Q(ram[6300]) );
  DFF ram_reg_1260__3_ ( .D(n10540), .CP(wclk), .Q(ram[6299]) );
  DFF ram_reg_1260__2_ ( .D(n10539), .CP(wclk), .Q(ram[6298]) );
  DFF ram_reg_1260__1_ ( .D(n10538), .CP(wclk), .Q(ram[6297]) );
  DFF ram_reg_1260__0_ ( .D(n10537), .CP(wclk), .Q(ram[6296]) );
  DFF ram_reg_1264__7_ ( .D(n10512), .CP(wclk), .Q(ram[6271]) );
  DFF ram_reg_1264__6_ ( .D(n10511), .CP(wclk), .Q(ram[6270]) );
  DFF ram_reg_1264__5_ ( .D(n10510), .CP(wclk), .Q(ram[6269]) );
  DFF ram_reg_1264__4_ ( .D(n10509), .CP(wclk), .Q(ram[6268]) );
  DFF ram_reg_1264__3_ ( .D(n10508), .CP(wclk), .Q(ram[6267]) );
  DFF ram_reg_1264__2_ ( .D(n10507), .CP(wclk), .Q(ram[6266]) );
  DFF ram_reg_1264__1_ ( .D(n10506), .CP(wclk), .Q(ram[6265]) );
  DFF ram_reg_1264__0_ ( .D(n10505), .CP(wclk), .Q(ram[6264]) );
  DFF ram_reg_1272__7_ ( .D(n10448), .CP(wclk), .Q(ram[6207]) );
  DFF ram_reg_1272__6_ ( .D(n10447), .CP(wclk), .Q(ram[6206]) );
  DFF ram_reg_1272__5_ ( .D(n10446), .CP(wclk), .Q(ram[6205]) );
  DFF ram_reg_1272__4_ ( .D(n10445), .CP(wclk), .Q(ram[6204]) );
  DFF ram_reg_1272__3_ ( .D(n10444), .CP(wclk), .Q(ram[6203]) );
  DFF ram_reg_1272__2_ ( .D(n10443), .CP(wclk), .Q(ram[6202]) );
  DFF ram_reg_1272__1_ ( .D(n10442), .CP(wclk), .Q(ram[6201]) );
  DFF ram_reg_1272__0_ ( .D(n10441), .CP(wclk), .Q(ram[6200]) );
  DFF ram_reg_1276__7_ ( .D(n10416), .CP(wclk), .Q(ram[6175]) );
  DFF ram_reg_1276__6_ ( .D(n10415), .CP(wclk), .Q(ram[6174]) );
  DFF ram_reg_1276__5_ ( .D(n10414), .CP(wclk), .Q(ram[6173]) );
  DFF ram_reg_1276__4_ ( .D(n10413), .CP(wclk), .Q(ram[6172]) );
  DFF ram_reg_1276__3_ ( .D(n10412), .CP(wclk), .Q(ram[6171]) );
  DFF ram_reg_1276__2_ ( .D(n10411), .CP(wclk), .Q(ram[6170]) );
  DFF ram_reg_1276__1_ ( .D(n10410), .CP(wclk), .Q(ram[6169]) );
  DFF ram_reg_1276__0_ ( .D(n10409), .CP(wclk), .Q(ram[6168]) );
  DFF ram_reg_1288__7_ ( .D(n10320), .CP(wclk), .Q(ram[6079]) );
  DFF ram_reg_1288__6_ ( .D(n10319), .CP(wclk), .Q(ram[6078]) );
  DFF ram_reg_1288__5_ ( .D(n10318), .CP(wclk), .Q(ram[6077]) );
  DFF ram_reg_1288__4_ ( .D(n10317), .CP(wclk), .Q(ram[6076]) );
  DFF ram_reg_1288__3_ ( .D(n10316), .CP(wclk), .Q(ram[6075]) );
  DFF ram_reg_1288__2_ ( .D(n10315), .CP(wclk), .Q(ram[6074]) );
  DFF ram_reg_1288__1_ ( .D(n10314), .CP(wclk), .Q(ram[6073]) );
  DFF ram_reg_1288__0_ ( .D(n10313), .CP(wclk), .Q(ram[6072]) );
  DFF ram_reg_1292__7_ ( .D(n10288), .CP(wclk), .Q(ram[6047]) );
  DFF ram_reg_1292__6_ ( .D(n10287), .CP(wclk), .Q(ram[6046]) );
  DFF ram_reg_1292__5_ ( .D(n10286), .CP(wclk), .Q(ram[6045]) );
  DFF ram_reg_1292__4_ ( .D(n10285), .CP(wclk), .Q(ram[6044]) );
  DFF ram_reg_1292__3_ ( .D(n10284), .CP(wclk), .Q(ram[6043]) );
  DFF ram_reg_1292__2_ ( .D(n10283), .CP(wclk), .Q(ram[6042]) );
  DFF ram_reg_1292__1_ ( .D(n10282), .CP(wclk), .Q(ram[6041]) );
  DFF ram_reg_1292__0_ ( .D(n10281), .CP(wclk), .Q(ram[6040]) );
  DFF ram_reg_1304__7_ ( .D(n10192), .CP(wclk), .Q(ram[5951]) );
  DFF ram_reg_1304__6_ ( .D(n10191), .CP(wclk), .Q(ram[5950]) );
  DFF ram_reg_1304__5_ ( .D(n10190), .CP(wclk), .Q(ram[5949]) );
  DFF ram_reg_1304__4_ ( .D(n10189), .CP(wclk), .Q(ram[5948]) );
  DFF ram_reg_1304__3_ ( .D(n10188), .CP(wclk), .Q(ram[5947]) );
  DFF ram_reg_1304__2_ ( .D(n10187), .CP(wclk), .Q(ram[5946]) );
  DFF ram_reg_1304__1_ ( .D(n10186), .CP(wclk), .Q(ram[5945]) );
  DFF ram_reg_1304__0_ ( .D(n10185), .CP(wclk), .Q(ram[5944]) );
  DFF ram_reg_1308__7_ ( .D(n10160), .CP(wclk), .Q(ram[5919]) );
  DFF ram_reg_1308__6_ ( .D(n10159), .CP(wclk), .Q(ram[5918]) );
  DFF ram_reg_1308__5_ ( .D(n10158), .CP(wclk), .Q(ram[5917]) );
  DFF ram_reg_1308__4_ ( .D(n10157), .CP(wclk), .Q(ram[5916]) );
  DFF ram_reg_1308__3_ ( .D(n10156), .CP(wclk), .Q(ram[5915]) );
  DFF ram_reg_1308__2_ ( .D(n10155), .CP(wclk), .Q(ram[5914]) );
  DFF ram_reg_1308__1_ ( .D(n10154), .CP(wclk), .Q(ram[5913]) );
  DFF ram_reg_1308__0_ ( .D(n10153), .CP(wclk), .Q(ram[5912]) );
  DFF ram_reg_1312__7_ ( .D(n10128), .CP(wclk), .Q(ram[5887]) );
  DFF ram_reg_1312__6_ ( .D(n10127), .CP(wclk), .Q(ram[5886]) );
  DFF ram_reg_1312__5_ ( .D(n10126), .CP(wclk), .Q(ram[5885]) );
  DFF ram_reg_1312__4_ ( .D(n10125), .CP(wclk), .Q(ram[5884]) );
  DFF ram_reg_1312__3_ ( .D(n10124), .CP(wclk), .Q(ram[5883]) );
  DFF ram_reg_1312__2_ ( .D(n10123), .CP(wclk), .Q(ram[5882]) );
  DFF ram_reg_1312__1_ ( .D(n10122), .CP(wclk), .Q(ram[5881]) );
  DFF ram_reg_1312__0_ ( .D(n10121), .CP(wclk), .Q(ram[5880]) );
  DFF ram_reg_1320__7_ ( .D(n10064), .CP(wclk), .Q(ram[5823]) );
  DFF ram_reg_1320__6_ ( .D(n10063), .CP(wclk), .Q(ram[5822]) );
  DFF ram_reg_1320__5_ ( .D(n10062), .CP(wclk), .Q(ram[5821]) );
  DFF ram_reg_1320__4_ ( .D(n10061), .CP(wclk), .Q(ram[5820]) );
  DFF ram_reg_1320__3_ ( .D(n10060), .CP(wclk), .Q(ram[5819]) );
  DFF ram_reg_1320__2_ ( .D(n10059), .CP(wclk), .Q(ram[5818]) );
  DFF ram_reg_1320__1_ ( .D(n10058), .CP(wclk), .Q(ram[5817]) );
  DFF ram_reg_1320__0_ ( .D(n10057), .CP(wclk), .Q(ram[5816]) );
  DFF ram_reg_1324__7_ ( .D(n10032), .CP(wclk), .Q(ram[5791]) );
  DFF ram_reg_1324__6_ ( .D(n10031), .CP(wclk), .Q(ram[5790]) );
  DFF ram_reg_1324__5_ ( .D(n10030), .CP(wclk), .Q(ram[5789]) );
  DFF ram_reg_1324__4_ ( .D(n10029), .CP(wclk), .Q(ram[5788]) );
  DFF ram_reg_1324__3_ ( .D(n10028), .CP(wclk), .Q(ram[5787]) );
  DFF ram_reg_1324__2_ ( .D(n10027), .CP(wclk), .Q(ram[5786]) );
  DFF ram_reg_1324__1_ ( .D(n10026), .CP(wclk), .Q(ram[5785]) );
  DFF ram_reg_1324__0_ ( .D(n10025), .CP(wclk), .Q(ram[5784]) );
  DFF ram_reg_1328__7_ ( .D(n10000), .CP(wclk), .Q(ram[5759]) );
  DFF ram_reg_1328__6_ ( .D(n9999), .CP(wclk), .Q(ram[5758]) );
  DFF ram_reg_1328__5_ ( .D(n9998), .CP(wclk), .Q(ram[5757]) );
  DFF ram_reg_1328__4_ ( .D(n9997), .CP(wclk), .Q(ram[5756]) );
  DFF ram_reg_1328__3_ ( .D(n9996), .CP(wclk), .Q(ram[5755]) );
  DFF ram_reg_1328__2_ ( .D(n9995), .CP(wclk), .Q(ram[5754]) );
  DFF ram_reg_1328__1_ ( .D(n9994), .CP(wclk), .Q(ram[5753]) );
  DFF ram_reg_1328__0_ ( .D(n9993), .CP(wclk), .Q(ram[5752]) );
  DFF ram_reg_1336__7_ ( .D(n9936), .CP(wclk), .Q(ram[5695]) );
  DFF ram_reg_1336__6_ ( .D(n9935), .CP(wclk), .Q(ram[5694]) );
  DFF ram_reg_1336__5_ ( .D(n9934), .CP(wclk), .Q(ram[5693]) );
  DFF ram_reg_1336__4_ ( .D(n9933), .CP(wclk), .Q(ram[5692]) );
  DFF ram_reg_1336__3_ ( .D(n9932), .CP(wclk), .Q(ram[5691]) );
  DFF ram_reg_1336__2_ ( .D(n9931), .CP(wclk), .Q(ram[5690]) );
  DFF ram_reg_1336__1_ ( .D(n9930), .CP(wclk), .Q(ram[5689]) );
  DFF ram_reg_1336__0_ ( .D(n9929), .CP(wclk), .Q(ram[5688]) );
  DFF ram_reg_1340__7_ ( .D(n9904), .CP(wclk), .Q(ram[5663]) );
  DFF ram_reg_1340__6_ ( .D(n9903), .CP(wclk), .Q(ram[5662]) );
  DFF ram_reg_1340__5_ ( .D(n9902), .CP(wclk), .Q(ram[5661]) );
  DFF ram_reg_1340__4_ ( .D(n9901), .CP(wclk), .Q(ram[5660]) );
  DFF ram_reg_1340__3_ ( .D(n9900), .CP(wclk), .Q(ram[5659]) );
  DFF ram_reg_1340__2_ ( .D(n9899), .CP(wclk), .Q(ram[5658]) );
  DFF ram_reg_1340__1_ ( .D(n9898), .CP(wclk), .Q(ram[5657]) );
  DFF ram_reg_1340__0_ ( .D(n9897), .CP(wclk), .Q(ram[5656]) );
  DFF ram_reg_1352__7_ ( .D(n9808), .CP(wclk), .Q(ram[5567]) );
  DFF ram_reg_1352__6_ ( .D(n9807), .CP(wclk), .Q(ram[5566]) );
  DFF ram_reg_1352__5_ ( .D(n9806), .CP(wclk), .Q(ram[5565]) );
  DFF ram_reg_1352__4_ ( .D(n9805), .CP(wclk), .Q(ram[5564]) );
  DFF ram_reg_1352__3_ ( .D(n9804), .CP(wclk), .Q(ram[5563]) );
  DFF ram_reg_1352__2_ ( .D(n9803), .CP(wclk), .Q(ram[5562]) );
  DFF ram_reg_1352__1_ ( .D(n9802), .CP(wclk), .Q(ram[5561]) );
  DFF ram_reg_1352__0_ ( .D(n9801), .CP(wclk), .Q(ram[5560]) );
  DFF ram_reg_1384__7_ ( .D(n9552), .CP(wclk), .Q(ram[5311]) );
  DFF ram_reg_1384__6_ ( .D(n9551), .CP(wclk), .Q(ram[5310]) );
  DFF ram_reg_1384__5_ ( .D(n9550), .CP(wclk), .Q(ram[5309]) );
  DFF ram_reg_1384__4_ ( .D(n9549), .CP(wclk), .Q(ram[5308]) );
  DFF ram_reg_1384__3_ ( .D(n9548), .CP(wclk), .Q(ram[5307]) );
  DFF ram_reg_1384__2_ ( .D(n9547), .CP(wclk), .Q(ram[5306]) );
  DFF ram_reg_1384__1_ ( .D(n9546), .CP(wclk), .Q(ram[5305]) );
  DFF ram_reg_1384__0_ ( .D(n9545), .CP(wclk), .Q(ram[5304]) );
  DFF ram_reg_1388__7_ ( .D(n9520), .CP(wclk), .Q(ram[5279]) );
  DFF ram_reg_1388__6_ ( .D(n9519), .CP(wclk), .Q(ram[5278]) );
  DFF ram_reg_1388__5_ ( .D(n9518), .CP(wclk), .Q(ram[5277]) );
  DFF ram_reg_1388__4_ ( .D(n9517), .CP(wclk), .Q(ram[5276]) );
  DFF ram_reg_1388__3_ ( .D(n9516), .CP(wclk), .Q(ram[5275]) );
  DFF ram_reg_1388__2_ ( .D(n9515), .CP(wclk), .Q(ram[5274]) );
  DFF ram_reg_1388__1_ ( .D(n9514), .CP(wclk), .Q(ram[5273]) );
  DFF ram_reg_1388__0_ ( .D(n9513), .CP(wclk), .Q(ram[5272]) );
  DFF ram_reg_1400__7_ ( .D(n9424), .CP(wclk), .Q(ram[5183]) );
  DFF ram_reg_1400__6_ ( .D(n9423), .CP(wclk), .Q(ram[5182]) );
  DFF ram_reg_1400__5_ ( .D(n9422), .CP(wclk), .Q(ram[5181]) );
  DFF ram_reg_1400__4_ ( .D(n9421), .CP(wclk), .Q(ram[5180]) );
  DFF ram_reg_1400__3_ ( .D(n9420), .CP(wclk), .Q(ram[5179]) );
  DFF ram_reg_1400__2_ ( .D(n9419), .CP(wclk), .Q(ram[5178]) );
  DFF ram_reg_1400__1_ ( .D(n9418), .CP(wclk), .Q(ram[5177]) );
  DFF ram_reg_1400__0_ ( .D(n9417), .CP(wclk), .Q(ram[5176]) );
  DFF ram_reg_1404__7_ ( .D(n9392), .CP(wclk), .Q(ram[5151]) );
  DFF ram_reg_1404__6_ ( .D(n9391), .CP(wclk), .Q(ram[5150]) );
  DFF ram_reg_1404__5_ ( .D(n9390), .CP(wclk), .Q(ram[5149]) );
  DFF ram_reg_1404__4_ ( .D(n9389), .CP(wclk), .Q(ram[5148]) );
  DFF ram_reg_1404__3_ ( .D(n9388), .CP(wclk), .Q(ram[5147]) );
  DFF ram_reg_1404__2_ ( .D(n9387), .CP(wclk), .Q(ram[5146]) );
  DFF ram_reg_1404__1_ ( .D(n9386), .CP(wclk), .Q(ram[5145]) );
  DFF ram_reg_1404__0_ ( .D(n9385), .CP(wclk), .Q(ram[5144]) );
  DFF ram_reg_1408__7_ ( .D(n9360), .CP(wclk), .Q(ram[5119]) );
  DFF ram_reg_1408__6_ ( .D(n9359), .CP(wclk), .Q(ram[5118]) );
  DFF ram_reg_1408__5_ ( .D(n9358), .CP(wclk), .Q(ram[5117]) );
  DFF ram_reg_1408__4_ ( .D(n9357), .CP(wclk), .Q(ram[5116]) );
  DFF ram_reg_1408__3_ ( .D(n9356), .CP(wclk), .Q(ram[5115]) );
  DFF ram_reg_1408__2_ ( .D(n9355), .CP(wclk), .Q(ram[5114]) );
  DFF ram_reg_1408__1_ ( .D(n9354), .CP(wclk), .Q(ram[5113]) );
  DFF ram_reg_1408__0_ ( .D(n9353), .CP(wclk), .Q(ram[5112]) );
  DFF ram_reg_1412__7_ ( .D(n9328), .CP(wclk), .Q(ram[5087]) );
  DFF ram_reg_1412__6_ ( .D(n9327), .CP(wclk), .Q(ram[5086]) );
  DFF ram_reg_1412__5_ ( .D(n9326), .CP(wclk), .Q(ram[5085]) );
  DFF ram_reg_1412__4_ ( .D(n9325), .CP(wclk), .Q(ram[5084]) );
  DFF ram_reg_1412__3_ ( .D(n9324), .CP(wclk), .Q(ram[5083]) );
  DFF ram_reg_1412__2_ ( .D(n9323), .CP(wclk), .Q(ram[5082]) );
  DFF ram_reg_1412__1_ ( .D(n9322), .CP(wclk), .Q(ram[5081]) );
  DFF ram_reg_1412__0_ ( .D(n9321), .CP(wclk), .Q(ram[5080]) );
  DFF ram_reg_1416__7_ ( .D(n9296), .CP(wclk), .Q(ram[5055]) );
  DFF ram_reg_1416__6_ ( .D(n9295), .CP(wclk), .Q(ram[5054]) );
  DFF ram_reg_1416__5_ ( .D(n9294), .CP(wclk), .Q(ram[5053]) );
  DFF ram_reg_1416__4_ ( .D(n9293), .CP(wclk), .Q(ram[5052]) );
  DFF ram_reg_1416__3_ ( .D(n9292), .CP(wclk), .Q(ram[5051]) );
  DFF ram_reg_1416__2_ ( .D(n9291), .CP(wclk), .Q(ram[5050]) );
  DFF ram_reg_1416__1_ ( .D(n9290), .CP(wclk), .Q(ram[5049]) );
  DFF ram_reg_1416__0_ ( .D(n9289), .CP(wclk), .Q(ram[5048]) );
  DFF ram_reg_1420__7_ ( .D(n9264), .CP(wclk), .Q(ram[5023]) );
  DFF ram_reg_1420__6_ ( .D(n9263), .CP(wclk), .Q(ram[5022]) );
  DFF ram_reg_1420__5_ ( .D(n9262), .CP(wclk), .Q(ram[5021]) );
  DFF ram_reg_1420__4_ ( .D(n9261), .CP(wclk), .Q(ram[5020]) );
  DFF ram_reg_1420__3_ ( .D(n9260), .CP(wclk), .Q(ram[5019]) );
  DFF ram_reg_1420__2_ ( .D(n9259), .CP(wclk), .Q(ram[5018]) );
  DFF ram_reg_1420__1_ ( .D(n9258), .CP(wclk), .Q(ram[5017]) );
  DFF ram_reg_1420__0_ ( .D(n9257), .CP(wclk), .Q(ram[5016]) );
  DFF ram_reg_1424__7_ ( .D(n9232), .CP(wclk), .Q(ram[4991]) );
  DFF ram_reg_1424__6_ ( .D(n9231), .CP(wclk), .Q(ram[4990]) );
  DFF ram_reg_1424__5_ ( .D(n9230), .CP(wclk), .Q(ram[4989]) );
  DFF ram_reg_1424__4_ ( .D(n9229), .CP(wclk), .Q(ram[4988]) );
  DFF ram_reg_1424__3_ ( .D(n9228), .CP(wclk), .Q(ram[4987]) );
  DFF ram_reg_1424__2_ ( .D(n9227), .CP(wclk), .Q(ram[4986]) );
  DFF ram_reg_1424__1_ ( .D(n9226), .CP(wclk), .Q(ram[4985]) );
  DFF ram_reg_1424__0_ ( .D(n9225), .CP(wclk), .Q(ram[4984]) );
  DFF ram_reg_1432__7_ ( .D(n9168), .CP(wclk), .Q(ram[4927]) );
  DFF ram_reg_1432__6_ ( .D(n9167), .CP(wclk), .Q(ram[4926]) );
  DFF ram_reg_1432__5_ ( .D(n9166), .CP(wclk), .Q(ram[4925]) );
  DFF ram_reg_1432__4_ ( .D(n9165), .CP(wclk), .Q(ram[4924]) );
  DFF ram_reg_1432__3_ ( .D(n9164), .CP(wclk), .Q(ram[4923]) );
  DFF ram_reg_1432__2_ ( .D(n9163), .CP(wclk), .Q(ram[4922]) );
  DFF ram_reg_1432__1_ ( .D(n9162), .CP(wclk), .Q(ram[4921]) );
  DFF ram_reg_1432__0_ ( .D(n9161), .CP(wclk), .Q(ram[4920]) );
  DFF ram_reg_1436__7_ ( .D(n9136), .CP(wclk), .Q(ram[4895]) );
  DFF ram_reg_1436__6_ ( .D(n9135), .CP(wclk), .Q(ram[4894]) );
  DFF ram_reg_1436__5_ ( .D(n9134), .CP(wclk), .Q(ram[4893]) );
  DFF ram_reg_1436__4_ ( .D(n9133), .CP(wclk), .Q(ram[4892]) );
  DFF ram_reg_1436__3_ ( .D(n9132), .CP(wclk), .Q(ram[4891]) );
  DFF ram_reg_1436__2_ ( .D(n9131), .CP(wclk), .Q(ram[4890]) );
  DFF ram_reg_1436__1_ ( .D(n9130), .CP(wclk), .Q(ram[4889]) );
  DFF ram_reg_1436__0_ ( .D(n9129), .CP(wclk), .Q(ram[4888]) );
  DFF ram_reg_1440__7_ ( .D(n9104), .CP(wclk), .Q(ram[4863]) );
  DFF ram_reg_1440__6_ ( .D(n9103), .CP(wclk), .Q(ram[4862]) );
  DFF ram_reg_1440__5_ ( .D(n9102), .CP(wclk), .Q(ram[4861]) );
  DFF ram_reg_1440__4_ ( .D(n9101), .CP(wclk), .Q(ram[4860]) );
  DFF ram_reg_1440__3_ ( .D(n9100), .CP(wclk), .Q(ram[4859]) );
  DFF ram_reg_1440__2_ ( .D(n9099), .CP(wclk), .Q(ram[4858]) );
  DFF ram_reg_1440__1_ ( .D(n9098), .CP(wclk), .Q(ram[4857]) );
  DFF ram_reg_1440__0_ ( .D(n9097), .CP(wclk), .Q(ram[4856]) );
  DFF ram_reg_1444__7_ ( .D(n9072), .CP(wclk), .Q(ram[4831]) );
  DFF ram_reg_1444__6_ ( .D(n9071), .CP(wclk), .Q(ram[4830]) );
  DFF ram_reg_1444__5_ ( .D(n9070), .CP(wclk), .Q(ram[4829]) );
  DFF ram_reg_1444__4_ ( .D(n9069), .CP(wclk), .Q(ram[4828]) );
  DFF ram_reg_1444__3_ ( .D(n9068), .CP(wclk), .Q(ram[4827]) );
  DFF ram_reg_1444__2_ ( .D(n9067), .CP(wclk), .Q(ram[4826]) );
  DFF ram_reg_1444__1_ ( .D(n9066), .CP(wclk), .Q(ram[4825]) );
  DFF ram_reg_1444__0_ ( .D(n9065), .CP(wclk), .Q(ram[4824]) );
  DFF ram_reg_1448__7_ ( .D(n9040), .CP(wclk), .Q(ram[4799]) );
  DFF ram_reg_1448__6_ ( .D(n9039), .CP(wclk), .Q(ram[4798]) );
  DFF ram_reg_1448__5_ ( .D(n9038), .CP(wclk), .Q(ram[4797]) );
  DFF ram_reg_1448__4_ ( .D(n9037), .CP(wclk), .Q(ram[4796]) );
  DFF ram_reg_1448__3_ ( .D(n9036), .CP(wclk), .Q(ram[4795]) );
  DFF ram_reg_1448__2_ ( .D(n9035), .CP(wclk), .Q(ram[4794]) );
  DFF ram_reg_1448__1_ ( .D(n9034), .CP(wclk), .Q(ram[4793]) );
  DFF ram_reg_1448__0_ ( .D(n9033), .CP(wclk), .Q(ram[4792]) );
  DFF ram_reg_1452__7_ ( .D(n9008), .CP(wclk), .Q(ram[4767]) );
  DFF ram_reg_1452__6_ ( .D(n9007), .CP(wclk), .Q(ram[4766]) );
  DFF ram_reg_1452__5_ ( .D(n9006), .CP(wclk), .Q(ram[4765]) );
  DFF ram_reg_1452__4_ ( .D(n9005), .CP(wclk), .Q(ram[4764]) );
  DFF ram_reg_1452__3_ ( .D(n9004), .CP(wclk), .Q(ram[4763]) );
  DFF ram_reg_1452__2_ ( .D(n9003), .CP(wclk), .Q(ram[4762]) );
  DFF ram_reg_1452__1_ ( .D(n9002), .CP(wclk), .Q(ram[4761]) );
  DFF ram_reg_1452__0_ ( .D(n9001), .CP(wclk), .Q(ram[4760]) );
  DFF ram_reg_1456__7_ ( .D(n8976), .CP(wclk), .Q(ram[4735]) );
  DFF ram_reg_1456__6_ ( .D(n8975), .CP(wclk), .Q(ram[4734]) );
  DFF ram_reg_1456__5_ ( .D(n8974), .CP(wclk), .Q(ram[4733]) );
  DFF ram_reg_1456__4_ ( .D(n8973), .CP(wclk), .Q(ram[4732]) );
  DFF ram_reg_1456__3_ ( .D(n8972), .CP(wclk), .Q(ram[4731]) );
  DFF ram_reg_1456__2_ ( .D(n8971), .CP(wclk), .Q(ram[4730]) );
  DFF ram_reg_1456__1_ ( .D(n8970), .CP(wclk), .Q(ram[4729]) );
  DFF ram_reg_1456__0_ ( .D(n8969), .CP(wclk), .Q(ram[4728]) );
  DFF ram_reg_1460__7_ ( .D(n8944), .CP(wclk), .Q(ram[4703]) );
  DFF ram_reg_1460__6_ ( .D(n8943), .CP(wclk), .Q(ram[4702]) );
  DFF ram_reg_1460__5_ ( .D(n8942), .CP(wclk), .Q(ram[4701]) );
  DFF ram_reg_1460__4_ ( .D(n8941), .CP(wclk), .Q(ram[4700]) );
  DFF ram_reg_1460__3_ ( .D(n8940), .CP(wclk), .Q(ram[4699]) );
  DFF ram_reg_1460__2_ ( .D(n8939), .CP(wclk), .Q(ram[4698]) );
  DFF ram_reg_1460__1_ ( .D(n8938), .CP(wclk), .Q(ram[4697]) );
  DFF ram_reg_1460__0_ ( .D(n8937), .CP(wclk), .Q(ram[4696]) );
  DFF ram_reg_1464__7_ ( .D(n8912), .CP(wclk), .Q(ram[4671]) );
  DFF ram_reg_1464__6_ ( .D(n8911), .CP(wclk), .Q(ram[4670]) );
  DFF ram_reg_1464__5_ ( .D(n8910), .CP(wclk), .Q(ram[4669]) );
  DFF ram_reg_1464__4_ ( .D(n8909), .CP(wclk), .Q(ram[4668]) );
  DFF ram_reg_1464__3_ ( .D(n8908), .CP(wclk), .Q(ram[4667]) );
  DFF ram_reg_1464__2_ ( .D(n8907), .CP(wclk), .Q(ram[4666]) );
  DFF ram_reg_1464__1_ ( .D(n8906), .CP(wclk), .Q(ram[4665]) );
  DFF ram_reg_1464__0_ ( .D(n8905), .CP(wclk), .Q(ram[4664]) );
  DFF ram_reg_1468__7_ ( .D(n8880), .CP(wclk), .Q(ram[4639]) );
  DFF ram_reg_1468__6_ ( .D(n8879), .CP(wclk), .Q(ram[4638]) );
  DFF ram_reg_1468__5_ ( .D(n8878), .CP(wclk), .Q(ram[4637]) );
  DFF ram_reg_1468__4_ ( .D(n8877), .CP(wclk), .Q(ram[4636]) );
  DFF ram_reg_1468__3_ ( .D(n8876), .CP(wclk), .Q(ram[4635]) );
  DFF ram_reg_1468__2_ ( .D(n8875), .CP(wclk), .Q(ram[4634]) );
  DFF ram_reg_1468__1_ ( .D(n8874), .CP(wclk), .Q(ram[4633]) );
  DFF ram_reg_1468__0_ ( .D(n8873), .CP(wclk), .Q(ram[4632]) );
  DFF ram_reg_1472__7_ ( .D(n8848), .CP(wclk), .Q(ram[4607]) );
  DFF ram_reg_1472__6_ ( .D(n8847), .CP(wclk), .Q(ram[4606]) );
  DFF ram_reg_1472__5_ ( .D(n8846), .CP(wclk), .Q(ram[4605]) );
  DFF ram_reg_1472__4_ ( .D(n8845), .CP(wclk), .Q(ram[4604]) );
  DFF ram_reg_1472__3_ ( .D(n8844), .CP(wclk), .Q(ram[4603]) );
  DFF ram_reg_1472__2_ ( .D(n8843), .CP(wclk), .Q(ram[4602]) );
  DFF ram_reg_1472__1_ ( .D(n8842), .CP(wclk), .Q(ram[4601]) );
  DFF ram_reg_1472__0_ ( .D(n8841), .CP(wclk), .Q(ram[4600]) );
  DFF ram_reg_1480__7_ ( .D(n8784), .CP(wclk), .Q(ram[4543]) );
  DFF ram_reg_1480__6_ ( .D(n8783), .CP(wclk), .Q(ram[4542]) );
  DFF ram_reg_1480__5_ ( .D(n8782), .CP(wclk), .Q(ram[4541]) );
  DFF ram_reg_1480__4_ ( .D(n8781), .CP(wclk), .Q(ram[4540]) );
  DFF ram_reg_1480__3_ ( .D(n8780), .CP(wclk), .Q(ram[4539]) );
  DFF ram_reg_1480__2_ ( .D(n8779), .CP(wclk), .Q(ram[4538]) );
  DFF ram_reg_1480__1_ ( .D(n8778), .CP(wclk), .Q(ram[4537]) );
  DFF ram_reg_1480__0_ ( .D(n8777), .CP(wclk), .Q(ram[4536]) );
  DFF ram_reg_1484__7_ ( .D(n8752), .CP(wclk), .Q(ram[4511]) );
  DFF ram_reg_1484__6_ ( .D(n8751), .CP(wclk), .Q(ram[4510]) );
  DFF ram_reg_1484__5_ ( .D(n8750), .CP(wclk), .Q(ram[4509]) );
  DFF ram_reg_1484__4_ ( .D(n8749), .CP(wclk), .Q(ram[4508]) );
  DFF ram_reg_1484__3_ ( .D(n8748), .CP(wclk), .Q(ram[4507]) );
  DFF ram_reg_1484__2_ ( .D(n8747), .CP(wclk), .Q(ram[4506]) );
  DFF ram_reg_1484__1_ ( .D(n8746), .CP(wclk), .Q(ram[4505]) );
  DFF ram_reg_1484__0_ ( .D(n8745), .CP(wclk), .Q(ram[4504]) );
  DFF ram_reg_1488__7_ ( .D(n8720), .CP(wclk), .Q(ram[4479]) );
  DFF ram_reg_1488__6_ ( .D(n8719), .CP(wclk), .Q(ram[4478]) );
  DFF ram_reg_1488__5_ ( .D(n8718), .CP(wclk), .Q(ram[4477]) );
  DFF ram_reg_1488__4_ ( .D(n8717), .CP(wclk), .Q(ram[4476]) );
  DFF ram_reg_1488__3_ ( .D(n8716), .CP(wclk), .Q(ram[4475]) );
  DFF ram_reg_1488__2_ ( .D(n8715), .CP(wclk), .Q(ram[4474]) );
  DFF ram_reg_1488__1_ ( .D(n8714), .CP(wclk), .Q(ram[4473]) );
  DFF ram_reg_1488__0_ ( .D(n8713), .CP(wclk), .Q(ram[4472]) );
  DFF ram_reg_1496__7_ ( .D(n8656), .CP(wclk), .Q(ram[4415]) );
  DFF ram_reg_1496__6_ ( .D(n8655), .CP(wclk), .Q(ram[4414]) );
  DFF ram_reg_1496__5_ ( .D(n8654), .CP(wclk), .Q(ram[4413]) );
  DFF ram_reg_1496__4_ ( .D(n8653), .CP(wclk), .Q(ram[4412]) );
  DFF ram_reg_1496__3_ ( .D(n8652), .CP(wclk), .Q(ram[4411]) );
  DFF ram_reg_1496__2_ ( .D(n8651), .CP(wclk), .Q(ram[4410]) );
  DFF ram_reg_1496__1_ ( .D(n8650), .CP(wclk), .Q(ram[4409]) );
  DFF ram_reg_1496__0_ ( .D(n8649), .CP(wclk), .Q(ram[4408]) );
  DFF ram_reg_1500__7_ ( .D(n8624), .CP(wclk), .Q(ram[4383]) );
  DFF ram_reg_1500__6_ ( .D(n8623), .CP(wclk), .Q(ram[4382]) );
  DFF ram_reg_1500__5_ ( .D(n8622), .CP(wclk), .Q(ram[4381]) );
  DFF ram_reg_1500__4_ ( .D(n8621), .CP(wclk), .Q(ram[4380]) );
  DFF ram_reg_1500__3_ ( .D(n8620), .CP(wclk), .Q(ram[4379]) );
  DFF ram_reg_1500__2_ ( .D(n8619), .CP(wclk), .Q(ram[4378]) );
  DFF ram_reg_1500__1_ ( .D(n8618), .CP(wclk), .Q(ram[4377]) );
  DFF ram_reg_1500__0_ ( .D(n8617), .CP(wclk), .Q(ram[4376]) );
  DFF ram_reg_1504__7_ ( .D(n8592), .CP(wclk), .Q(ram[4351]) );
  DFF ram_reg_1504__6_ ( .D(n8591), .CP(wclk), .Q(ram[4350]) );
  DFF ram_reg_1504__5_ ( .D(n8590), .CP(wclk), .Q(ram[4349]) );
  DFF ram_reg_1504__4_ ( .D(n8589), .CP(wclk), .Q(ram[4348]) );
  DFF ram_reg_1504__3_ ( .D(n8588), .CP(wclk), .Q(ram[4347]) );
  DFF ram_reg_1504__2_ ( .D(n8587), .CP(wclk), .Q(ram[4346]) );
  DFF ram_reg_1504__1_ ( .D(n8586), .CP(wclk), .Q(ram[4345]) );
  DFF ram_reg_1504__0_ ( .D(n8585), .CP(wclk), .Q(ram[4344]) );
  DFF ram_reg_1508__7_ ( .D(n8560), .CP(wclk), .Q(ram[4319]) );
  DFF ram_reg_1508__6_ ( .D(n8559), .CP(wclk), .Q(ram[4318]) );
  DFF ram_reg_1508__5_ ( .D(n8558), .CP(wclk), .Q(ram[4317]) );
  DFF ram_reg_1508__4_ ( .D(n8557), .CP(wclk), .Q(ram[4316]) );
  DFF ram_reg_1508__3_ ( .D(n8556), .CP(wclk), .Q(ram[4315]) );
  DFF ram_reg_1508__2_ ( .D(n8555), .CP(wclk), .Q(ram[4314]) );
  DFF ram_reg_1508__1_ ( .D(n8554), .CP(wclk), .Q(ram[4313]) );
  DFF ram_reg_1508__0_ ( .D(n8553), .CP(wclk), .Q(ram[4312]) );
  DFF ram_reg_1512__7_ ( .D(n8528), .CP(wclk), .Q(ram[4287]) );
  DFF ram_reg_1512__6_ ( .D(n8527), .CP(wclk), .Q(ram[4286]) );
  DFF ram_reg_1512__5_ ( .D(n8526), .CP(wclk), .Q(ram[4285]) );
  DFF ram_reg_1512__4_ ( .D(n8525), .CP(wclk), .Q(ram[4284]) );
  DFF ram_reg_1512__3_ ( .D(n8524), .CP(wclk), .Q(ram[4283]) );
  DFF ram_reg_1512__2_ ( .D(n8523), .CP(wclk), .Q(ram[4282]) );
  DFF ram_reg_1512__1_ ( .D(n8522), .CP(wclk), .Q(ram[4281]) );
  DFF ram_reg_1512__0_ ( .D(n8521), .CP(wclk), .Q(ram[4280]) );
  DFF ram_reg_1516__7_ ( .D(n8496), .CP(wclk), .Q(ram[4255]) );
  DFF ram_reg_1516__6_ ( .D(n8495), .CP(wclk), .Q(ram[4254]) );
  DFF ram_reg_1516__5_ ( .D(n8494), .CP(wclk), .Q(ram[4253]) );
  DFF ram_reg_1516__4_ ( .D(n8493), .CP(wclk), .Q(ram[4252]) );
  DFF ram_reg_1516__3_ ( .D(n8492), .CP(wclk), .Q(ram[4251]) );
  DFF ram_reg_1516__2_ ( .D(n8491), .CP(wclk), .Q(ram[4250]) );
  DFF ram_reg_1516__1_ ( .D(n8490), .CP(wclk), .Q(ram[4249]) );
  DFF ram_reg_1516__0_ ( .D(n8489), .CP(wclk), .Q(ram[4248]) );
  DFF ram_reg_1520__7_ ( .D(n8464), .CP(wclk), .Q(ram[4223]) );
  DFF ram_reg_1520__6_ ( .D(n8463), .CP(wclk), .Q(ram[4222]) );
  DFF ram_reg_1520__5_ ( .D(n8462), .CP(wclk), .Q(ram[4221]) );
  DFF ram_reg_1520__4_ ( .D(n8461), .CP(wclk), .Q(ram[4220]) );
  DFF ram_reg_1520__3_ ( .D(n8460), .CP(wclk), .Q(ram[4219]) );
  DFF ram_reg_1520__2_ ( .D(n8459), .CP(wclk), .Q(ram[4218]) );
  DFF ram_reg_1520__1_ ( .D(n8458), .CP(wclk), .Q(ram[4217]) );
  DFF ram_reg_1520__0_ ( .D(n8457), .CP(wclk), .Q(ram[4216]) );
  DFF ram_reg_1524__7_ ( .D(n8432), .CP(wclk), .Q(ram[4191]) );
  DFF ram_reg_1524__6_ ( .D(n8431), .CP(wclk), .Q(ram[4190]) );
  DFF ram_reg_1524__5_ ( .D(n8430), .CP(wclk), .Q(ram[4189]) );
  DFF ram_reg_1524__4_ ( .D(n8429), .CP(wclk), .Q(ram[4188]) );
  DFF ram_reg_1524__3_ ( .D(n8428), .CP(wclk), .Q(ram[4187]) );
  DFF ram_reg_1524__2_ ( .D(n8427), .CP(wclk), .Q(ram[4186]) );
  DFF ram_reg_1524__1_ ( .D(n8426), .CP(wclk), .Q(ram[4185]) );
  DFF ram_reg_1524__0_ ( .D(n8425), .CP(wclk), .Q(ram[4184]) );
  DFF ram_reg_1528__7_ ( .D(n8400), .CP(wclk), .Q(ram[4159]) );
  DFF ram_reg_1528__6_ ( .D(n8399), .CP(wclk), .Q(ram[4158]) );
  DFF ram_reg_1528__5_ ( .D(n8398), .CP(wclk), .Q(ram[4157]) );
  DFF ram_reg_1528__4_ ( .D(n8397), .CP(wclk), .Q(ram[4156]) );
  DFF ram_reg_1528__3_ ( .D(n8396), .CP(wclk), .Q(ram[4155]) );
  DFF ram_reg_1528__2_ ( .D(n8395), .CP(wclk), .Q(ram[4154]) );
  DFF ram_reg_1528__1_ ( .D(n8394), .CP(wclk), .Q(ram[4153]) );
  DFF ram_reg_1528__0_ ( .D(n8393), .CP(wclk), .Q(ram[4152]) );
  DFF ram_reg_1532__7_ ( .D(n8368), .CP(wclk), .Q(ram[4127]) );
  DFF ram_reg_1532__6_ ( .D(n8367), .CP(wclk), .Q(ram[4126]) );
  DFF ram_reg_1532__5_ ( .D(n8366), .CP(wclk), .Q(ram[4125]) );
  DFF ram_reg_1532__4_ ( .D(n8365), .CP(wclk), .Q(ram[4124]) );
  DFF ram_reg_1532__3_ ( .D(n8364), .CP(wclk), .Q(ram[4123]) );
  DFF ram_reg_1532__2_ ( .D(n8363), .CP(wclk), .Q(ram[4122]) );
  DFF ram_reg_1532__1_ ( .D(n8362), .CP(wclk), .Q(ram[4121]) );
  DFF ram_reg_1532__0_ ( .D(n8361), .CP(wclk), .Q(ram[4120]) );
  DFF ram_reg_1544__7_ ( .D(n8272), .CP(wclk), .Q(ram[4031]) );
  DFF ram_reg_1544__6_ ( .D(n8271), .CP(wclk), .Q(ram[4030]) );
  DFF ram_reg_1544__5_ ( .D(n8270), .CP(wclk), .Q(ram[4029]) );
  DFF ram_reg_1544__4_ ( .D(n8269), .CP(wclk), .Q(ram[4028]) );
  DFF ram_reg_1544__3_ ( .D(n8268), .CP(wclk), .Q(ram[4027]) );
  DFF ram_reg_1544__2_ ( .D(n8267), .CP(wclk), .Q(ram[4026]) );
  DFF ram_reg_1544__1_ ( .D(n8266), .CP(wclk), .Q(ram[4025]) );
  DFF ram_reg_1544__0_ ( .D(n8265), .CP(wclk), .Q(ram[4024]) );
  DFF ram_reg_1576__7_ ( .D(n8016), .CP(wclk), .Q(ram[3775]) );
  DFF ram_reg_1576__6_ ( .D(n8015), .CP(wclk), .Q(ram[3774]) );
  DFF ram_reg_1576__5_ ( .D(n8014), .CP(wclk), .Q(ram[3773]) );
  DFF ram_reg_1576__4_ ( .D(n8013), .CP(wclk), .Q(ram[3772]) );
  DFF ram_reg_1576__3_ ( .D(n8012), .CP(wclk), .Q(ram[3771]) );
  DFF ram_reg_1576__2_ ( .D(n8011), .CP(wclk), .Q(ram[3770]) );
  DFF ram_reg_1576__1_ ( .D(n8010), .CP(wclk), .Q(ram[3769]) );
  DFF ram_reg_1576__0_ ( .D(n8009), .CP(wclk), .Q(ram[3768]) );
  DFF ram_reg_1580__7_ ( .D(n7984), .CP(wclk), .Q(ram[3743]) );
  DFF ram_reg_1580__6_ ( .D(n7983), .CP(wclk), .Q(ram[3742]) );
  DFF ram_reg_1580__5_ ( .D(n7982), .CP(wclk), .Q(ram[3741]) );
  DFF ram_reg_1580__4_ ( .D(n7981), .CP(wclk), .Q(ram[3740]) );
  DFF ram_reg_1580__3_ ( .D(n7980), .CP(wclk), .Q(ram[3739]) );
  DFF ram_reg_1580__2_ ( .D(n7979), .CP(wclk), .Q(ram[3738]) );
  DFF ram_reg_1580__1_ ( .D(n7978), .CP(wclk), .Q(ram[3737]) );
  DFF ram_reg_1580__0_ ( .D(n7977), .CP(wclk), .Q(ram[3736]) );
  DFF ram_reg_1592__7_ ( .D(n7888), .CP(wclk), .Q(ram[3647]) );
  DFF ram_reg_1592__6_ ( .D(n7887), .CP(wclk), .Q(ram[3646]) );
  DFF ram_reg_1592__5_ ( .D(n7886), .CP(wclk), .Q(ram[3645]) );
  DFF ram_reg_1592__4_ ( .D(n7885), .CP(wclk), .Q(ram[3644]) );
  DFF ram_reg_1592__3_ ( .D(n7884), .CP(wclk), .Q(ram[3643]) );
  DFF ram_reg_1592__2_ ( .D(n7883), .CP(wclk), .Q(ram[3642]) );
  DFF ram_reg_1592__1_ ( .D(n7882), .CP(wclk), .Q(ram[3641]) );
  DFF ram_reg_1592__0_ ( .D(n7881), .CP(wclk), .Q(ram[3640]) );
  DFF ram_reg_1596__7_ ( .D(n7856), .CP(wclk), .Q(ram[3615]) );
  DFF ram_reg_1596__6_ ( .D(n7855), .CP(wclk), .Q(ram[3614]) );
  DFF ram_reg_1596__5_ ( .D(n7854), .CP(wclk), .Q(ram[3613]) );
  DFF ram_reg_1596__4_ ( .D(n7853), .CP(wclk), .Q(ram[3612]) );
  DFF ram_reg_1596__3_ ( .D(n7852), .CP(wclk), .Q(ram[3611]) );
  DFF ram_reg_1596__2_ ( .D(n7851), .CP(wclk), .Q(ram[3610]) );
  DFF ram_reg_1596__1_ ( .D(n7850), .CP(wclk), .Q(ram[3609]) );
  DFF ram_reg_1596__0_ ( .D(n7849), .CP(wclk), .Q(ram[3608]) );
  DFF ram_reg_1664__7_ ( .D(n7312), .CP(wclk), .Q(ram[3071]) );
  DFF ram_reg_1664__6_ ( .D(n7311), .CP(wclk), .Q(ram[3070]) );
  DFF ram_reg_1664__5_ ( .D(n7310), .CP(wclk), .Q(ram[3069]) );
  DFF ram_reg_1664__4_ ( .D(n7309), .CP(wclk), .Q(ram[3068]) );
  DFF ram_reg_1664__3_ ( .D(n7308), .CP(wclk), .Q(ram[3067]) );
  DFF ram_reg_1664__2_ ( .D(n7307), .CP(wclk), .Q(ram[3066]) );
  DFF ram_reg_1664__1_ ( .D(n7306), .CP(wclk), .Q(ram[3065]) );
  DFF ram_reg_1664__0_ ( .D(n7305), .CP(wclk), .Q(ram[3064]) );
  DFF ram_reg_1672__7_ ( .D(n7248), .CP(wclk), .Q(ram[3007]) );
  DFF ram_reg_1672__6_ ( .D(n7247), .CP(wclk), .Q(ram[3006]) );
  DFF ram_reg_1672__5_ ( .D(n7246), .CP(wclk), .Q(ram[3005]) );
  DFF ram_reg_1672__4_ ( .D(n7245), .CP(wclk), .Q(ram[3004]) );
  DFF ram_reg_1672__3_ ( .D(n7244), .CP(wclk), .Q(ram[3003]) );
  DFF ram_reg_1672__2_ ( .D(n7243), .CP(wclk), .Q(ram[3002]) );
  DFF ram_reg_1672__1_ ( .D(n7242), .CP(wclk), .Q(ram[3001]) );
  DFF ram_reg_1672__0_ ( .D(n7241), .CP(wclk), .Q(ram[3000]) );
  DFF ram_reg_1676__7_ ( .D(n7216), .CP(wclk), .Q(ram[2975]) );
  DFF ram_reg_1676__6_ ( .D(n7215), .CP(wclk), .Q(ram[2974]) );
  DFF ram_reg_1676__5_ ( .D(n7214), .CP(wclk), .Q(ram[2973]) );
  DFF ram_reg_1676__4_ ( .D(n7213), .CP(wclk), .Q(ram[2972]) );
  DFF ram_reg_1676__3_ ( .D(n7212), .CP(wclk), .Q(ram[2971]) );
  DFF ram_reg_1676__2_ ( .D(n7211), .CP(wclk), .Q(ram[2970]) );
  DFF ram_reg_1676__1_ ( .D(n7210), .CP(wclk), .Q(ram[2969]) );
  DFF ram_reg_1676__0_ ( .D(n7209), .CP(wclk), .Q(ram[2968]) );
  DFF ram_reg_1688__7_ ( .D(n7120), .CP(wclk), .Q(ram[2879]) );
  DFF ram_reg_1688__6_ ( .D(n7119), .CP(wclk), .Q(ram[2878]) );
  DFF ram_reg_1688__5_ ( .D(n7118), .CP(wclk), .Q(ram[2877]) );
  DFF ram_reg_1688__4_ ( .D(n7117), .CP(wclk), .Q(ram[2876]) );
  DFF ram_reg_1688__3_ ( .D(n7116), .CP(wclk), .Q(ram[2875]) );
  DFF ram_reg_1688__2_ ( .D(n7115), .CP(wclk), .Q(ram[2874]) );
  DFF ram_reg_1688__1_ ( .D(n7114), .CP(wclk), .Q(ram[2873]) );
  DFF ram_reg_1688__0_ ( .D(n7113), .CP(wclk), .Q(ram[2872]) );
  DFF ram_reg_1692__7_ ( .D(n7088), .CP(wclk), .Q(ram[2847]) );
  DFF ram_reg_1692__6_ ( .D(n7087), .CP(wclk), .Q(ram[2846]) );
  DFF ram_reg_1692__5_ ( .D(n7086), .CP(wclk), .Q(ram[2845]) );
  DFF ram_reg_1692__4_ ( .D(n7085), .CP(wclk), .Q(ram[2844]) );
  DFF ram_reg_1692__3_ ( .D(n7084), .CP(wclk), .Q(ram[2843]) );
  DFF ram_reg_1692__2_ ( .D(n7083), .CP(wclk), .Q(ram[2842]) );
  DFF ram_reg_1692__1_ ( .D(n7082), .CP(wclk), .Q(ram[2841]) );
  DFF ram_reg_1692__0_ ( .D(n7081), .CP(wclk), .Q(ram[2840]) );
  DFF ram_reg_1696__7_ ( .D(n7056), .CP(wclk), .Q(ram[2815]) );
  DFF ram_reg_1696__6_ ( .D(n7055), .CP(wclk), .Q(ram[2814]) );
  DFF ram_reg_1696__5_ ( .D(n7054), .CP(wclk), .Q(ram[2813]) );
  DFF ram_reg_1696__4_ ( .D(n7053), .CP(wclk), .Q(ram[2812]) );
  DFF ram_reg_1696__3_ ( .D(n7052), .CP(wclk), .Q(ram[2811]) );
  DFF ram_reg_1696__2_ ( .D(n7051), .CP(wclk), .Q(ram[2810]) );
  DFF ram_reg_1696__1_ ( .D(n7050), .CP(wclk), .Q(ram[2809]) );
  DFF ram_reg_1696__0_ ( .D(n7049), .CP(wclk), .Q(ram[2808]) );
  DFF ram_reg_1704__7_ ( .D(n6992), .CP(wclk), .Q(ram[2751]) );
  DFF ram_reg_1704__6_ ( .D(n6991), .CP(wclk), .Q(ram[2750]) );
  DFF ram_reg_1704__5_ ( .D(n6990), .CP(wclk), .Q(ram[2749]) );
  DFF ram_reg_1704__4_ ( .D(n6989), .CP(wclk), .Q(ram[2748]) );
  DFF ram_reg_1704__3_ ( .D(n6988), .CP(wclk), .Q(ram[2747]) );
  DFF ram_reg_1704__2_ ( .D(n6987), .CP(wclk), .Q(ram[2746]) );
  DFF ram_reg_1704__1_ ( .D(n6986), .CP(wclk), .Q(ram[2745]) );
  DFF ram_reg_1704__0_ ( .D(n6985), .CP(wclk), .Q(ram[2744]) );
  DFF ram_reg_1708__7_ ( .D(n6960), .CP(wclk), .Q(ram[2719]) );
  DFF ram_reg_1708__6_ ( .D(n6959), .CP(wclk), .Q(ram[2718]) );
  DFF ram_reg_1708__5_ ( .D(n6958), .CP(wclk), .Q(ram[2717]) );
  DFF ram_reg_1708__4_ ( .D(n6957), .CP(wclk), .Q(ram[2716]) );
  DFF ram_reg_1708__3_ ( .D(n6956), .CP(wclk), .Q(ram[2715]) );
  DFF ram_reg_1708__2_ ( .D(n6955), .CP(wclk), .Q(ram[2714]) );
  DFF ram_reg_1708__1_ ( .D(n6954), .CP(wclk), .Q(ram[2713]) );
  DFF ram_reg_1708__0_ ( .D(n6953), .CP(wclk), .Q(ram[2712]) );
  DFF ram_reg_1712__7_ ( .D(n6928), .CP(wclk), .Q(ram[2687]) );
  DFF ram_reg_1712__6_ ( .D(n6927), .CP(wclk), .Q(ram[2686]) );
  DFF ram_reg_1712__5_ ( .D(n6926), .CP(wclk), .Q(ram[2685]) );
  DFF ram_reg_1712__4_ ( .D(n6925), .CP(wclk), .Q(ram[2684]) );
  DFF ram_reg_1712__3_ ( .D(n6924), .CP(wclk), .Q(ram[2683]) );
  DFF ram_reg_1712__2_ ( .D(n6923), .CP(wclk), .Q(ram[2682]) );
  DFF ram_reg_1712__1_ ( .D(n6922), .CP(wclk), .Q(ram[2681]) );
  DFF ram_reg_1712__0_ ( .D(n6921), .CP(wclk), .Q(ram[2680]) );
  DFF ram_reg_1720__7_ ( .D(n6864), .CP(wclk), .Q(ram[2623]) );
  DFF ram_reg_1720__6_ ( .D(n6863), .CP(wclk), .Q(ram[2622]) );
  DFF ram_reg_1720__5_ ( .D(n6862), .CP(wclk), .Q(ram[2621]) );
  DFF ram_reg_1720__4_ ( .D(n6861), .CP(wclk), .Q(ram[2620]) );
  DFF ram_reg_1720__3_ ( .D(n6860), .CP(wclk), .Q(ram[2619]) );
  DFF ram_reg_1720__2_ ( .D(n6859), .CP(wclk), .Q(ram[2618]) );
  DFF ram_reg_1720__1_ ( .D(n6858), .CP(wclk), .Q(ram[2617]) );
  DFF ram_reg_1720__0_ ( .D(n6857), .CP(wclk), .Q(ram[2616]) );
  DFF ram_reg_1724__7_ ( .D(n6832), .CP(wclk), .Q(ram[2591]) );
  DFF ram_reg_1724__6_ ( .D(n6831), .CP(wclk), .Q(ram[2590]) );
  DFF ram_reg_1724__5_ ( .D(n6830), .CP(wclk), .Q(ram[2589]) );
  DFF ram_reg_1724__4_ ( .D(n6829), .CP(wclk), .Q(ram[2588]) );
  DFF ram_reg_1724__3_ ( .D(n6828), .CP(wclk), .Q(ram[2587]) );
  DFF ram_reg_1724__2_ ( .D(n6827), .CP(wclk), .Q(ram[2586]) );
  DFF ram_reg_1724__1_ ( .D(n6826), .CP(wclk), .Q(ram[2585]) );
  DFF ram_reg_1724__0_ ( .D(n6825), .CP(wclk), .Q(ram[2584]) );
  DFF ram_reg_1736__7_ ( .D(n6736), .CP(wclk), .Q(ram[2495]) );
  DFF ram_reg_1736__6_ ( .D(n6735), .CP(wclk), .Q(ram[2494]) );
  DFF ram_reg_1736__5_ ( .D(n6734), .CP(wclk), .Q(ram[2493]) );
  DFF ram_reg_1736__4_ ( .D(n6733), .CP(wclk), .Q(ram[2492]) );
  DFF ram_reg_1736__3_ ( .D(n6732), .CP(wclk), .Q(ram[2491]) );
  DFF ram_reg_1736__2_ ( .D(n6731), .CP(wclk), .Q(ram[2490]) );
  DFF ram_reg_1736__1_ ( .D(n6730), .CP(wclk), .Q(ram[2489]) );
  DFF ram_reg_1736__0_ ( .D(n6729), .CP(wclk), .Q(ram[2488]) );
  DFF ram_reg_1740__7_ ( .D(n6704), .CP(wclk), .Q(ram[2463]) );
  DFF ram_reg_1740__6_ ( .D(n6703), .CP(wclk), .Q(ram[2462]) );
  DFF ram_reg_1740__5_ ( .D(n6702), .CP(wclk), .Q(ram[2461]) );
  DFF ram_reg_1740__4_ ( .D(n6701), .CP(wclk), .Q(ram[2460]) );
  DFF ram_reg_1740__3_ ( .D(n6700), .CP(wclk), .Q(ram[2459]) );
  DFF ram_reg_1740__2_ ( .D(n6699), .CP(wclk), .Q(ram[2458]) );
  DFF ram_reg_1740__1_ ( .D(n6698), .CP(wclk), .Q(ram[2457]) );
  DFF ram_reg_1740__0_ ( .D(n6697), .CP(wclk), .Q(ram[2456]) );
  DFF ram_reg_1752__7_ ( .D(n6608), .CP(wclk), .Q(ram[2367]) );
  DFF ram_reg_1752__6_ ( .D(n6607), .CP(wclk), .Q(ram[2366]) );
  DFF ram_reg_1752__5_ ( .D(n6606), .CP(wclk), .Q(ram[2365]) );
  DFF ram_reg_1752__4_ ( .D(n6605), .CP(wclk), .Q(ram[2364]) );
  DFF ram_reg_1752__3_ ( .D(n6604), .CP(wclk), .Q(ram[2363]) );
  DFF ram_reg_1752__2_ ( .D(n6603), .CP(wclk), .Q(ram[2362]) );
  DFF ram_reg_1752__1_ ( .D(n6602), .CP(wclk), .Q(ram[2361]) );
  DFF ram_reg_1752__0_ ( .D(n6601), .CP(wclk), .Q(ram[2360]) );
  DFF ram_reg_1760__7_ ( .D(n6544), .CP(wclk), .Q(ram[2303]) );
  DFF ram_reg_1760__6_ ( .D(n6543), .CP(wclk), .Q(ram[2302]) );
  DFF ram_reg_1760__5_ ( .D(n6542), .CP(wclk), .Q(ram[2301]) );
  DFF ram_reg_1760__4_ ( .D(n6541), .CP(wclk), .Q(ram[2300]) );
  DFF ram_reg_1760__3_ ( .D(n6540), .CP(wclk), .Q(ram[2299]) );
  DFF ram_reg_1760__2_ ( .D(n6539), .CP(wclk), .Q(ram[2298]) );
  DFF ram_reg_1760__1_ ( .D(n6538), .CP(wclk), .Q(ram[2297]) );
  DFF ram_reg_1760__0_ ( .D(n6537), .CP(wclk), .Q(ram[2296]) );
  DFF ram_reg_1768__7_ ( .D(n6480), .CP(wclk), .Q(ram[2239]) );
  DFF ram_reg_1768__6_ ( .D(n6479), .CP(wclk), .Q(ram[2238]) );
  DFF ram_reg_1768__5_ ( .D(n6478), .CP(wclk), .Q(ram[2237]) );
  DFF ram_reg_1768__4_ ( .D(n6477), .CP(wclk), .Q(ram[2236]) );
  DFF ram_reg_1768__3_ ( .D(n6476), .CP(wclk), .Q(ram[2235]) );
  DFF ram_reg_1768__2_ ( .D(n6475), .CP(wclk), .Q(ram[2234]) );
  DFF ram_reg_1768__1_ ( .D(n6474), .CP(wclk), .Q(ram[2233]) );
  DFF ram_reg_1768__0_ ( .D(n6473), .CP(wclk), .Q(ram[2232]) );
  DFF ram_reg_1772__7_ ( .D(n6448), .CP(wclk), .Q(ram[2207]) );
  DFF ram_reg_1772__6_ ( .D(n6447), .CP(wclk), .Q(ram[2206]) );
  DFF ram_reg_1772__5_ ( .D(n6446), .CP(wclk), .Q(ram[2205]) );
  DFF ram_reg_1772__4_ ( .D(n6445), .CP(wclk), .Q(ram[2204]) );
  DFF ram_reg_1772__3_ ( .D(n6444), .CP(wclk), .Q(ram[2203]) );
  DFF ram_reg_1772__2_ ( .D(n6443), .CP(wclk), .Q(ram[2202]) );
  DFF ram_reg_1772__1_ ( .D(n6442), .CP(wclk), .Q(ram[2201]) );
  DFF ram_reg_1772__0_ ( .D(n6441), .CP(wclk), .Q(ram[2200]) );
  DFF ram_reg_1776__7_ ( .D(n6416), .CP(wclk), .Q(ram[2175]) );
  DFF ram_reg_1776__6_ ( .D(n6415), .CP(wclk), .Q(ram[2174]) );
  DFF ram_reg_1776__5_ ( .D(n6414), .CP(wclk), .Q(ram[2173]) );
  DFF ram_reg_1776__4_ ( .D(n6413), .CP(wclk), .Q(ram[2172]) );
  DFF ram_reg_1776__3_ ( .D(n6412), .CP(wclk), .Q(ram[2171]) );
  DFF ram_reg_1776__2_ ( .D(n6411), .CP(wclk), .Q(ram[2170]) );
  DFF ram_reg_1776__1_ ( .D(n6410), .CP(wclk), .Q(ram[2169]) );
  DFF ram_reg_1776__0_ ( .D(n6409), .CP(wclk), .Q(ram[2168]) );
  DFF ram_reg_1784__7_ ( .D(n6352), .CP(wclk), .Q(ram[2111]) );
  DFF ram_reg_1784__6_ ( .D(n6351), .CP(wclk), .Q(ram[2110]) );
  DFF ram_reg_1784__5_ ( .D(n6350), .CP(wclk), .Q(ram[2109]) );
  DFF ram_reg_1784__4_ ( .D(n6349), .CP(wclk), .Q(ram[2108]) );
  DFF ram_reg_1784__3_ ( .D(n6348), .CP(wclk), .Q(ram[2107]) );
  DFF ram_reg_1784__2_ ( .D(n6347), .CP(wclk), .Q(ram[2106]) );
  DFF ram_reg_1784__1_ ( .D(n6346), .CP(wclk), .Q(ram[2105]) );
  DFF ram_reg_1784__0_ ( .D(n6345), .CP(wclk), .Q(ram[2104]) );
  DFF ram_reg_1788__7_ ( .D(n6320), .CP(wclk), .Q(ram[2079]) );
  DFF ram_reg_1788__6_ ( .D(n6319), .CP(wclk), .Q(ram[2078]) );
  DFF ram_reg_1788__5_ ( .D(n6318), .CP(wclk), .Q(ram[2077]) );
  DFF ram_reg_1788__4_ ( .D(n6317), .CP(wclk), .Q(ram[2076]) );
  DFF ram_reg_1788__3_ ( .D(n6316), .CP(wclk), .Q(ram[2075]) );
  DFF ram_reg_1788__2_ ( .D(n6315), .CP(wclk), .Q(ram[2074]) );
  DFF ram_reg_1788__1_ ( .D(n6314), .CP(wclk), .Q(ram[2073]) );
  DFF ram_reg_1788__0_ ( .D(n6313), .CP(wclk), .Q(ram[2072]) );
  DFF ram_reg_1800__7_ ( .D(n6224), .CP(wclk), .Q(ram[1983]) );
  DFF ram_reg_1800__6_ ( .D(n6223), .CP(wclk), .Q(ram[1982]) );
  DFF ram_reg_1800__5_ ( .D(n6222), .CP(wclk), .Q(ram[1981]) );
  DFF ram_reg_1800__4_ ( .D(n6221), .CP(wclk), .Q(ram[1980]) );
  DFF ram_reg_1800__3_ ( .D(n6220), .CP(wclk), .Q(ram[1979]) );
  DFF ram_reg_1800__2_ ( .D(n6219), .CP(wclk), .Q(ram[1978]) );
  DFF ram_reg_1800__1_ ( .D(n6218), .CP(wclk), .Q(ram[1977]) );
  DFF ram_reg_1800__0_ ( .D(n6217), .CP(wclk), .Q(ram[1976]) );
  DFF ram_reg_1832__7_ ( .D(n5968), .CP(wclk), .Q(ram[1727]) );
  DFF ram_reg_1832__6_ ( .D(n5967), .CP(wclk), .Q(ram[1726]) );
  DFF ram_reg_1832__5_ ( .D(n5966), .CP(wclk), .Q(ram[1725]) );
  DFF ram_reg_1832__4_ ( .D(n5965), .CP(wclk), .Q(ram[1724]) );
  DFF ram_reg_1832__3_ ( .D(n5964), .CP(wclk), .Q(ram[1723]) );
  DFF ram_reg_1832__2_ ( .D(n5963), .CP(wclk), .Q(ram[1722]) );
  DFF ram_reg_1832__1_ ( .D(n5962), .CP(wclk), .Q(ram[1721]) );
  DFF ram_reg_1832__0_ ( .D(n5961), .CP(wclk), .Q(ram[1720]) );
  DFF ram_reg_1836__7_ ( .D(n5936), .CP(wclk), .Q(ram[1695]) );
  DFF ram_reg_1836__6_ ( .D(n5935), .CP(wclk), .Q(ram[1694]) );
  DFF ram_reg_1836__5_ ( .D(n5934), .CP(wclk), .Q(ram[1693]) );
  DFF ram_reg_1836__4_ ( .D(n5933), .CP(wclk), .Q(ram[1692]) );
  DFF ram_reg_1836__3_ ( .D(n5932), .CP(wclk), .Q(ram[1691]) );
  DFF ram_reg_1836__2_ ( .D(n5931), .CP(wclk), .Q(ram[1690]) );
  DFF ram_reg_1836__1_ ( .D(n5930), .CP(wclk), .Q(ram[1689]) );
  DFF ram_reg_1836__0_ ( .D(n5929), .CP(wclk), .Q(ram[1688]) );
  DFF ram_reg_1848__7_ ( .D(n5840), .CP(wclk), .Q(ram[1599]) );
  DFF ram_reg_1848__6_ ( .D(n5839), .CP(wclk), .Q(ram[1598]) );
  DFF ram_reg_1848__5_ ( .D(n5838), .CP(wclk), .Q(ram[1597]) );
  DFF ram_reg_1848__4_ ( .D(n5837), .CP(wclk), .Q(ram[1596]) );
  DFF ram_reg_1848__3_ ( .D(n5836), .CP(wclk), .Q(ram[1595]) );
  DFF ram_reg_1848__2_ ( .D(n5835), .CP(wclk), .Q(ram[1594]) );
  DFF ram_reg_1848__1_ ( .D(n5834), .CP(wclk), .Q(ram[1593]) );
  DFF ram_reg_1848__0_ ( .D(n5833), .CP(wclk), .Q(ram[1592]) );
  DFF ram_reg_1852__7_ ( .D(n5808), .CP(wclk), .Q(ram[1567]) );
  DFF ram_reg_1852__6_ ( .D(n5807), .CP(wclk), .Q(ram[1566]) );
  DFF ram_reg_1852__5_ ( .D(n5806), .CP(wclk), .Q(ram[1565]) );
  DFF ram_reg_1852__4_ ( .D(n5805), .CP(wclk), .Q(ram[1564]) );
  DFF ram_reg_1852__3_ ( .D(n5804), .CP(wclk), .Q(ram[1563]) );
  DFF ram_reg_1852__2_ ( .D(n5803), .CP(wclk), .Q(ram[1562]) );
  DFF ram_reg_1852__1_ ( .D(n5802), .CP(wclk), .Q(ram[1561]) );
  DFF ram_reg_1852__0_ ( .D(n5801), .CP(wclk), .Q(ram[1560]) );
  DFF ram_reg_1920__7_ ( .D(n5264), .CP(wclk), .Q(ram[1023]) );
  DFF ram_reg_1920__6_ ( .D(n5263), .CP(wclk), .Q(ram[1022]) );
  DFF ram_reg_1920__5_ ( .D(n5262), .CP(wclk), .Q(ram[1021]) );
  DFF ram_reg_1920__4_ ( .D(n5261), .CP(wclk), .Q(ram[1020]) );
  DFF ram_reg_1920__3_ ( .D(n5260), .CP(wclk), .Q(ram[1019]) );
  DFF ram_reg_1920__2_ ( .D(n5259), .CP(wclk), .Q(ram[1018]) );
  DFF ram_reg_1920__1_ ( .D(n5258), .CP(wclk), .Q(ram[1017]) );
  DFF ram_reg_1920__0_ ( .D(n5257), .CP(wclk), .Q(ram[1016]) );
  DFF ram_reg_1928__7_ ( .D(n5200), .CP(wclk), .Q(ram[959]) );
  DFF ram_reg_1928__6_ ( .D(n5199), .CP(wclk), .Q(ram[958]) );
  DFF ram_reg_1928__5_ ( .D(n5198), .CP(wclk), .Q(ram[957]) );
  DFF ram_reg_1928__4_ ( .D(n5197), .CP(wclk), .Q(ram[956]) );
  DFF ram_reg_1928__3_ ( .D(n5196), .CP(wclk), .Q(ram[955]) );
  DFF ram_reg_1928__2_ ( .D(n5195), .CP(wclk), .Q(ram[954]) );
  DFF ram_reg_1928__1_ ( .D(n5194), .CP(wclk), .Q(ram[953]) );
  DFF ram_reg_1928__0_ ( .D(n5193), .CP(wclk), .Q(ram[952]) );
  DFF ram_reg_1932__7_ ( .D(n5168), .CP(wclk), .Q(ram[927]) );
  DFF ram_reg_1932__6_ ( .D(n5167), .CP(wclk), .Q(ram[926]) );
  DFF ram_reg_1932__5_ ( .D(n5166), .CP(wclk), .Q(ram[925]) );
  DFF ram_reg_1932__4_ ( .D(n5165), .CP(wclk), .Q(ram[924]) );
  DFF ram_reg_1932__3_ ( .D(n5164), .CP(wclk), .Q(ram[923]) );
  DFF ram_reg_1932__2_ ( .D(n5163), .CP(wclk), .Q(ram[922]) );
  DFF ram_reg_1932__1_ ( .D(n5162), .CP(wclk), .Q(ram[921]) );
  DFF ram_reg_1932__0_ ( .D(n5161), .CP(wclk), .Q(ram[920]) );
  DFF ram_reg_1944__7_ ( .D(n5072), .CP(wclk), .Q(ram[831]) );
  DFF ram_reg_1944__6_ ( .D(n5071), .CP(wclk), .Q(ram[830]) );
  DFF ram_reg_1944__5_ ( .D(n5070), .CP(wclk), .Q(ram[829]) );
  DFF ram_reg_1944__4_ ( .D(n5069), .CP(wclk), .Q(ram[828]) );
  DFF ram_reg_1944__3_ ( .D(n5068), .CP(wclk), .Q(ram[827]) );
  DFF ram_reg_1944__2_ ( .D(n5067), .CP(wclk), .Q(ram[826]) );
  DFF ram_reg_1944__1_ ( .D(n5066), .CP(wclk), .Q(ram[825]) );
  DFF ram_reg_1944__0_ ( .D(n5065), .CP(wclk), .Q(ram[824]) );
  DFF ram_reg_1948__7_ ( .D(n5040), .CP(wclk), .Q(ram[799]) );
  DFF ram_reg_1948__6_ ( .D(n5039), .CP(wclk), .Q(ram[798]) );
  DFF ram_reg_1948__5_ ( .D(n5038), .CP(wclk), .Q(ram[797]) );
  DFF ram_reg_1948__4_ ( .D(n5037), .CP(wclk), .Q(ram[796]) );
  DFF ram_reg_1948__3_ ( .D(n5036), .CP(wclk), .Q(ram[795]) );
  DFF ram_reg_1948__2_ ( .D(n5035), .CP(wclk), .Q(ram[794]) );
  DFF ram_reg_1948__1_ ( .D(n5034), .CP(wclk), .Q(ram[793]) );
  DFF ram_reg_1948__0_ ( .D(n5033), .CP(wclk), .Q(ram[792]) );
  DFF ram_reg_1952__7_ ( .D(n5008), .CP(wclk), .Q(ram[767]) );
  DFF ram_reg_1952__6_ ( .D(n5007), .CP(wclk), .Q(ram[766]) );
  DFF ram_reg_1952__5_ ( .D(n5006), .CP(wclk), .Q(ram[765]) );
  DFF ram_reg_1952__4_ ( .D(n5005), .CP(wclk), .Q(ram[764]) );
  DFF ram_reg_1952__3_ ( .D(n5004), .CP(wclk), .Q(ram[763]) );
  DFF ram_reg_1952__2_ ( .D(n5003), .CP(wclk), .Q(ram[762]) );
  DFF ram_reg_1952__1_ ( .D(n5002), .CP(wclk), .Q(ram[761]) );
  DFF ram_reg_1952__0_ ( .D(n5001), .CP(wclk), .Q(ram[760]) );
  DFF ram_reg_1960__7_ ( .D(n4944), .CP(wclk), .Q(ram[703]) );
  DFF ram_reg_1960__6_ ( .D(n4943), .CP(wclk), .Q(ram[702]) );
  DFF ram_reg_1960__5_ ( .D(n4942), .CP(wclk), .Q(ram[701]) );
  DFF ram_reg_1960__4_ ( .D(n4941), .CP(wclk), .Q(ram[700]) );
  DFF ram_reg_1960__3_ ( .D(n4940), .CP(wclk), .Q(ram[699]) );
  DFF ram_reg_1960__2_ ( .D(n4939), .CP(wclk), .Q(ram[698]) );
  DFF ram_reg_1960__1_ ( .D(n4938), .CP(wclk), .Q(ram[697]) );
  DFF ram_reg_1960__0_ ( .D(n4937), .CP(wclk), .Q(ram[696]) );
  DFF ram_reg_1964__7_ ( .D(n4912), .CP(wclk), .Q(ram[671]) );
  DFF ram_reg_1964__6_ ( .D(n4911), .CP(wclk), .Q(ram[670]) );
  DFF ram_reg_1964__5_ ( .D(n4910), .CP(wclk), .Q(ram[669]) );
  DFF ram_reg_1964__4_ ( .D(n4909), .CP(wclk), .Q(ram[668]) );
  DFF ram_reg_1964__3_ ( .D(n4908), .CP(wclk), .Q(ram[667]) );
  DFF ram_reg_1964__2_ ( .D(n4907), .CP(wclk), .Q(ram[666]) );
  DFF ram_reg_1964__1_ ( .D(n4906), .CP(wclk), .Q(ram[665]) );
  DFF ram_reg_1964__0_ ( .D(n4905), .CP(wclk), .Q(ram[664]) );
  DFF ram_reg_1968__7_ ( .D(n4880), .CP(wclk), .Q(ram[639]) );
  DFF ram_reg_1968__6_ ( .D(n4879), .CP(wclk), .Q(ram[638]) );
  DFF ram_reg_1968__5_ ( .D(n4878), .CP(wclk), .Q(ram[637]) );
  DFF ram_reg_1968__4_ ( .D(n4877), .CP(wclk), .Q(ram[636]) );
  DFF ram_reg_1968__3_ ( .D(n4876), .CP(wclk), .Q(ram[635]) );
  DFF ram_reg_1968__2_ ( .D(n4875), .CP(wclk), .Q(ram[634]) );
  DFF ram_reg_1968__1_ ( .D(n4874), .CP(wclk), .Q(ram[633]) );
  DFF ram_reg_1968__0_ ( .D(n4873), .CP(wclk), .Q(ram[632]) );
  DFF ram_reg_1976__7_ ( .D(n4816), .CP(wclk), .Q(ram[575]) );
  DFF ram_reg_1976__6_ ( .D(n4815), .CP(wclk), .Q(ram[574]) );
  DFF ram_reg_1976__5_ ( .D(n4814), .CP(wclk), .Q(ram[573]) );
  DFF ram_reg_1976__4_ ( .D(n4813), .CP(wclk), .Q(ram[572]) );
  DFF ram_reg_1976__3_ ( .D(n4812), .CP(wclk), .Q(ram[571]) );
  DFF ram_reg_1976__2_ ( .D(n4811), .CP(wclk), .Q(ram[570]) );
  DFF ram_reg_1976__1_ ( .D(n4810), .CP(wclk), .Q(ram[569]) );
  DFF ram_reg_1976__0_ ( .D(n4809), .CP(wclk), .Q(ram[568]) );
  DFF ram_reg_1980__7_ ( .D(n4784), .CP(wclk), .Q(ram[543]) );
  DFF ram_reg_1980__6_ ( .D(n4783), .CP(wclk), .Q(ram[542]) );
  DFF ram_reg_1980__5_ ( .D(n4782), .CP(wclk), .Q(ram[541]) );
  DFF ram_reg_1980__4_ ( .D(n4781), .CP(wclk), .Q(ram[540]) );
  DFF ram_reg_1980__3_ ( .D(n4780), .CP(wclk), .Q(ram[539]) );
  DFF ram_reg_1980__2_ ( .D(n4779), .CP(wclk), .Q(ram[538]) );
  DFF ram_reg_1980__1_ ( .D(n4778), .CP(wclk), .Q(ram[537]) );
  DFF ram_reg_1980__0_ ( .D(n4777), .CP(wclk), .Q(ram[536]) );
  DFF ram_reg_1992__7_ ( .D(n4688), .CP(wclk), .Q(ram[447]) );
  DFF ram_reg_1992__6_ ( .D(n4687), .CP(wclk), .Q(ram[446]) );
  DFF ram_reg_1992__5_ ( .D(n4686), .CP(wclk), .Q(ram[445]) );
  DFF ram_reg_1992__4_ ( .D(n4685), .CP(wclk), .Q(ram[444]) );
  DFF ram_reg_1992__3_ ( .D(n4684), .CP(wclk), .Q(ram[443]) );
  DFF ram_reg_1992__2_ ( .D(n4683), .CP(wclk), .Q(ram[442]) );
  DFF ram_reg_1992__1_ ( .D(n4682), .CP(wclk), .Q(ram[441]) );
  DFF ram_reg_1992__0_ ( .D(n4681), .CP(wclk), .Q(ram[440]) );
  DFF ram_reg_1996__7_ ( .D(n4656), .CP(wclk), .Q(ram[415]) );
  DFF ram_reg_1996__6_ ( .D(n4655), .CP(wclk), .Q(ram[414]) );
  DFF ram_reg_1996__5_ ( .D(n4654), .CP(wclk), .Q(ram[413]) );
  DFF ram_reg_1996__4_ ( .D(n4653), .CP(wclk), .Q(ram[412]) );
  DFF ram_reg_1996__3_ ( .D(n4652), .CP(wclk), .Q(ram[411]) );
  DFF ram_reg_1996__2_ ( .D(n4651), .CP(wclk), .Q(ram[410]) );
  DFF ram_reg_1996__1_ ( .D(n4650), .CP(wclk), .Q(ram[409]) );
  DFF ram_reg_1996__0_ ( .D(n4649), .CP(wclk), .Q(ram[408]) );
  DFF ram_reg_2008__7_ ( .D(n4560), .CP(wclk), .Q(ram[319]) );
  DFF ram_reg_2008__6_ ( .D(n4559), .CP(wclk), .Q(ram[318]) );
  DFF ram_reg_2008__5_ ( .D(n4558), .CP(wclk), .Q(ram[317]) );
  DFF ram_reg_2008__4_ ( .D(n4557), .CP(wclk), .Q(ram[316]) );
  DFF ram_reg_2008__3_ ( .D(n4556), .CP(wclk), .Q(ram[315]) );
  DFF ram_reg_2008__2_ ( .D(n4555), .CP(wclk), .Q(ram[314]) );
  DFF ram_reg_2008__1_ ( .D(n4554), .CP(wclk), .Q(ram[313]) );
  DFF ram_reg_2008__0_ ( .D(n4553), .CP(wclk), .Q(ram[312]) );
  DFF ram_reg_2012__7_ ( .D(n4528), .CP(wclk), .Q(ram[287]) );
  DFF ram_reg_2012__6_ ( .D(n4527), .CP(wclk), .Q(ram[286]) );
  DFF ram_reg_2012__5_ ( .D(n4526), .CP(wclk), .Q(ram[285]) );
  DFF ram_reg_2012__4_ ( .D(n4525), .CP(wclk), .Q(ram[284]) );
  DFF ram_reg_2012__3_ ( .D(n4524), .CP(wclk), .Q(ram[283]) );
  DFF ram_reg_2012__2_ ( .D(n4523), .CP(wclk), .Q(ram[282]) );
  DFF ram_reg_2012__1_ ( .D(n4522), .CP(wclk), .Q(ram[281]) );
  DFF ram_reg_2012__0_ ( .D(n4521), .CP(wclk), .Q(ram[280]) );
  DFF ram_reg_2016__7_ ( .D(n4496), .CP(wclk), .Q(ram[255]) );
  DFF ram_reg_2016__6_ ( .D(n4495), .CP(wclk), .Q(ram[254]) );
  DFF ram_reg_2016__5_ ( .D(n4494), .CP(wclk), .Q(ram[253]) );
  DFF ram_reg_2016__4_ ( .D(n4493), .CP(wclk), .Q(ram[252]) );
  DFF ram_reg_2016__3_ ( .D(n4492), .CP(wclk), .Q(ram[251]) );
  DFF ram_reg_2016__2_ ( .D(n4491), .CP(wclk), .Q(ram[250]) );
  DFF ram_reg_2016__1_ ( .D(n4490), .CP(wclk), .Q(ram[249]) );
  DFF ram_reg_2016__0_ ( .D(n4489), .CP(wclk), .Q(ram[248]) );
  DFF ram_reg_2024__7_ ( .D(n4432), .CP(wclk), .Q(ram[191]) );
  DFF ram_reg_2024__6_ ( .D(n4431), .CP(wclk), .Q(ram[190]) );
  DFF ram_reg_2024__5_ ( .D(n4430), .CP(wclk), .Q(ram[189]) );
  DFF ram_reg_2024__4_ ( .D(n4429), .CP(wclk), .Q(ram[188]) );
  DFF ram_reg_2024__3_ ( .D(n4428), .CP(wclk), .Q(ram[187]) );
  DFF ram_reg_2024__2_ ( .D(n4427), .CP(wclk), .Q(ram[186]) );
  DFF ram_reg_2024__1_ ( .D(n4426), .CP(wclk), .Q(ram[185]) );
  DFF ram_reg_2024__0_ ( .D(n4425), .CP(wclk), .Q(ram[184]) );
  DFF ram_reg_2028__7_ ( .D(n4400), .CP(wclk), .Q(ram[159]) );
  DFF ram_reg_2028__6_ ( .D(n4399), .CP(wclk), .Q(ram[158]) );
  DFF ram_reg_2028__5_ ( .D(n4398), .CP(wclk), .Q(ram[157]) );
  DFF ram_reg_2028__4_ ( .D(n4397), .CP(wclk), .Q(ram[156]) );
  DFF ram_reg_2028__3_ ( .D(n4396), .CP(wclk), .Q(ram[155]) );
  DFF ram_reg_2028__2_ ( .D(n4395), .CP(wclk), .Q(ram[154]) );
  DFF ram_reg_2028__1_ ( .D(n4394), .CP(wclk), .Q(ram[153]) );
  DFF ram_reg_2028__0_ ( .D(n4393), .CP(wclk), .Q(ram[152]) );
  DFF ram_reg_2032__7_ ( .D(n4368), .CP(wclk), .Q(ram[127]) );
  DFF ram_reg_2032__6_ ( .D(n4367), .CP(wclk), .Q(ram[126]) );
  DFF ram_reg_2032__5_ ( .D(n4366), .CP(wclk), .Q(ram[125]) );
  DFF ram_reg_2032__4_ ( .D(n4365), .CP(wclk), .Q(ram[124]) );
  DFF ram_reg_2032__3_ ( .D(n4364), .CP(wclk), .Q(ram[123]) );
  DFF ram_reg_2032__2_ ( .D(n4363), .CP(wclk), .Q(ram[122]) );
  DFF ram_reg_2032__1_ ( .D(n4362), .CP(wclk), .Q(ram[121]) );
  DFF ram_reg_2032__0_ ( .D(n4361), .CP(wclk), .Q(ram[120]) );
  DFF ram_reg_2040__7_ ( .D(n4304), .CP(wclk), .Q(ram[63]) );
  DFF ram_reg_2040__6_ ( .D(n4303), .CP(wclk), .Q(ram[62]) );
  DFF ram_reg_2040__5_ ( .D(n4302), .CP(wclk), .Q(ram[61]) );
  DFF ram_reg_2040__4_ ( .D(n4301), .CP(wclk), .Q(ram[60]) );
  DFF ram_reg_2040__3_ ( .D(n4300), .CP(wclk), .Q(ram[59]) );
  DFF ram_reg_2040__2_ ( .D(n4299), .CP(wclk), .Q(ram[58]) );
  DFF ram_reg_2040__1_ ( .D(n4298), .CP(wclk), .Q(ram[57]) );
  DFF ram_reg_2040__0_ ( .D(n4297), .CP(wclk), .Q(ram[56]) );
  DFF ram_reg_2044__7_ ( .D(n4272), .CP(wclk), .Q(ram[31]) );
  DFF ram_reg_2044__6_ ( .D(n4271), .CP(wclk), .Q(ram[30]) );
  DFF ram_reg_2044__5_ ( .D(n4270), .CP(wclk), .Q(ram[29]) );
  DFF ram_reg_2044__4_ ( .D(n4269), .CP(wclk), .Q(ram[28]) );
  DFF ram_reg_2044__3_ ( .D(n4268), .CP(wclk), .Q(ram[27]) );
  DFF ram_reg_2044__2_ ( .D(n4267), .CP(wclk), .Q(ram[26]) );
  DFF ram_reg_2044__1_ ( .D(n4266), .CP(wclk), .Q(ram[25]) );
  DFF ram_reg_2044__0_ ( .D(n4265), .CP(wclk), .Q(ram[24]) );
  DFF ram_reg_138__7_ ( .D(n19520), .CP(wclk), .Q(ram[15279]) );
  DFF ram_reg_138__6_ ( .D(n19519), .CP(wclk), .Q(ram[15278]) );
  DFF ram_reg_138__5_ ( .D(n19518), .CP(wclk), .Q(ram[15277]) );
  DFF ram_reg_138__4_ ( .D(n19517), .CP(wclk), .Q(ram[15276]) );
  DFF ram_reg_138__3_ ( .D(n19516), .CP(wclk), .Q(ram[15275]) );
  DFF ram_reg_138__2_ ( .D(n19515), .CP(wclk), .Q(ram[15274]) );
  DFF ram_reg_138__1_ ( .D(n19514), .CP(wclk), .Q(ram[15273]) );
  DFF ram_reg_138__0_ ( .D(n19513), .CP(wclk), .Q(ram[15272]) );
  DFF ram_reg_170__7_ ( .D(n19264), .CP(wclk), .Q(ram[15023]) );
  DFF ram_reg_170__6_ ( .D(n19263), .CP(wclk), .Q(ram[15022]) );
  DFF ram_reg_170__5_ ( .D(n19262), .CP(wclk), .Q(ram[15021]) );
  DFF ram_reg_170__4_ ( .D(n19261), .CP(wclk), .Q(ram[15020]) );
  DFF ram_reg_170__3_ ( .D(n19260), .CP(wclk), .Q(ram[15019]) );
  DFF ram_reg_170__2_ ( .D(n19259), .CP(wclk), .Q(ram[15018]) );
  DFF ram_reg_170__1_ ( .D(n19258), .CP(wclk), .Q(ram[15017]) );
  DFF ram_reg_170__0_ ( .D(n19257), .CP(wclk), .Q(ram[15016]) );
  DFF ram_reg_174__7_ ( .D(n19232), .CP(wclk), .Q(ram[14991]) );
  DFF ram_reg_174__6_ ( .D(n19231), .CP(wclk), .Q(ram[14990]) );
  DFF ram_reg_174__5_ ( .D(n19230), .CP(wclk), .Q(ram[14989]) );
  DFF ram_reg_174__4_ ( .D(n19229), .CP(wclk), .Q(ram[14988]) );
  DFF ram_reg_174__3_ ( .D(n19228), .CP(wclk), .Q(ram[14987]) );
  DFF ram_reg_174__2_ ( .D(n19227), .CP(wclk), .Q(ram[14986]) );
  DFF ram_reg_174__1_ ( .D(n19226), .CP(wclk), .Q(ram[14985]) );
  DFF ram_reg_174__0_ ( .D(n19225), .CP(wclk), .Q(ram[14984]) );
  DFF ram_reg_186__7_ ( .D(n19136), .CP(wclk), .Q(ram[14895]) );
  DFF ram_reg_186__6_ ( .D(n19135), .CP(wclk), .Q(ram[14894]) );
  DFF ram_reg_186__5_ ( .D(n19134), .CP(wclk), .Q(ram[14893]) );
  DFF ram_reg_186__4_ ( .D(n19133), .CP(wclk), .Q(ram[14892]) );
  DFF ram_reg_186__3_ ( .D(n19132), .CP(wclk), .Q(ram[14891]) );
  DFF ram_reg_186__2_ ( .D(n19131), .CP(wclk), .Q(ram[14890]) );
  DFF ram_reg_186__1_ ( .D(n19130), .CP(wclk), .Q(ram[14889]) );
  DFF ram_reg_186__0_ ( .D(n19129), .CP(wclk), .Q(ram[14888]) );
  DFF ram_reg_190__7_ ( .D(n19104), .CP(wclk), .Q(ram[14863]) );
  DFF ram_reg_190__6_ ( .D(n19103), .CP(wclk), .Q(ram[14862]) );
  DFF ram_reg_190__5_ ( .D(n19102), .CP(wclk), .Q(ram[14861]) );
  DFF ram_reg_190__4_ ( .D(n19101), .CP(wclk), .Q(ram[14860]) );
  DFF ram_reg_190__3_ ( .D(n19100), .CP(wclk), .Q(ram[14859]) );
  DFF ram_reg_190__2_ ( .D(n19099), .CP(wclk), .Q(ram[14858]) );
  DFF ram_reg_190__1_ ( .D(n19098), .CP(wclk), .Q(ram[14857]) );
  DFF ram_reg_190__0_ ( .D(n19097), .CP(wclk), .Q(ram[14856]) );
  DFF ram_reg_234__7_ ( .D(n18752), .CP(wclk), .Q(ram[14511]) );
  DFF ram_reg_234__6_ ( .D(n18751), .CP(wclk), .Q(ram[14510]) );
  DFF ram_reg_234__5_ ( .D(n18750), .CP(wclk), .Q(ram[14509]) );
  DFF ram_reg_234__4_ ( .D(n18749), .CP(wclk), .Q(ram[14508]) );
  DFF ram_reg_234__3_ ( .D(n18748), .CP(wclk), .Q(ram[14507]) );
  DFF ram_reg_234__2_ ( .D(n18747), .CP(wclk), .Q(ram[14506]) );
  DFF ram_reg_234__1_ ( .D(n18746), .CP(wclk), .Q(ram[14505]) );
  DFF ram_reg_234__0_ ( .D(n18745), .CP(wclk), .Q(ram[14504]) );
  DFF ram_reg_250__7_ ( .D(n18624), .CP(wclk), .Q(ram[14383]) );
  DFF ram_reg_250__6_ ( .D(n18623), .CP(wclk), .Q(ram[14382]) );
  DFF ram_reg_250__5_ ( .D(n18622), .CP(wclk), .Q(ram[14381]) );
  DFF ram_reg_250__4_ ( .D(n18621), .CP(wclk), .Q(ram[14380]) );
  DFF ram_reg_250__3_ ( .D(n18620), .CP(wclk), .Q(ram[14379]) );
  DFF ram_reg_250__2_ ( .D(n18619), .CP(wclk), .Q(ram[14378]) );
  DFF ram_reg_250__1_ ( .D(n18618), .CP(wclk), .Q(ram[14377]) );
  DFF ram_reg_250__0_ ( .D(n18617), .CP(wclk), .Q(ram[14376]) );
  DFF ram_reg_254__7_ ( .D(n18592), .CP(wclk), .Q(ram[14351]) );
  DFF ram_reg_254__6_ ( .D(n18591), .CP(wclk), .Q(ram[14350]) );
  DFF ram_reg_254__5_ ( .D(n18590), .CP(wclk), .Q(ram[14349]) );
  DFF ram_reg_254__4_ ( .D(n18589), .CP(wclk), .Q(ram[14348]) );
  DFF ram_reg_254__3_ ( .D(n18588), .CP(wclk), .Q(ram[14347]) );
  DFF ram_reg_254__2_ ( .D(n18587), .CP(wclk), .Q(ram[14346]) );
  DFF ram_reg_254__1_ ( .D(n18586), .CP(wclk), .Q(ram[14345]) );
  DFF ram_reg_254__0_ ( .D(n18585), .CP(wclk), .Q(ram[14344]) );
  DFF ram_reg_314__7_ ( .D(n18112), .CP(wclk), .Q(ram[13871]) );
  DFF ram_reg_314__6_ ( .D(n18111), .CP(wclk), .Q(ram[13870]) );
  DFF ram_reg_314__5_ ( .D(n18110), .CP(wclk), .Q(ram[13869]) );
  DFF ram_reg_314__4_ ( .D(n18109), .CP(wclk), .Q(ram[13868]) );
  DFF ram_reg_314__3_ ( .D(n18108), .CP(wclk), .Q(ram[13867]) );
  DFF ram_reg_314__2_ ( .D(n18107), .CP(wclk), .Q(ram[13866]) );
  DFF ram_reg_314__1_ ( .D(n18106), .CP(wclk), .Q(ram[13865]) );
  DFF ram_reg_314__0_ ( .D(n18105), .CP(wclk), .Q(ram[13864]) );
  DFF ram_reg_394__7_ ( .D(n17472), .CP(wclk), .Q(ram[13231]) );
  DFF ram_reg_394__6_ ( .D(n17471), .CP(wclk), .Q(ram[13230]) );
  DFF ram_reg_394__5_ ( .D(n17470), .CP(wclk), .Q(ram[13229]) );
  DFF ram_reg_394__4_ ( .D(n17469), .CP(wclk), .Q(ram[13228]) );
  DFF ram_reg_394__3_ ( .D(n17468), .CP(wclk), .Q(ram[13227]) );
  DFF ram_reg_394__2_ ( .D(n17467), .CP(wclk), .Q(ram[13226]) );
  DFF ram_reg_394__1_ ( .D(n17466), .CP(wclk), .Q(ram[13225]) );
  DFF ram_reg_394__0_ ( .D(n17465), .CP(wclk), .Q(ram[13224]) );
  DFF ram_reg_398__7_ ( .D(n17440), .CP(wclk), .Q(ram[13199]) );
  DFF ram_reg_398__6_ ( .D(n17439), .CP(wclk), .Q(ram[13198]) );
  DFF ram_reg_398__5_ ( .D(n17438), .CP(wclk), .Q(ram[13197]) );
  DFF ram_reg_398__4_ ( .D(n17437), .CP(wclk), .Q(ram[13196]) );
  DFF ram_reg_398__3_ ( .D(n17436), .CP(wclk), .Q(ram[13195]) );
  DFF ram_reg_398__2_ ( .D(n17435), .CP(wclk), .Q(ram[13194]) );
  DFF ram_reg_398__1_ ( .D(n17434), .CP(wclk), .Q(ram[13193]) );
  DFF ram_reg_398__0_ ( .D(n17433), .CP(wclk), .Q(ram[13192]) );
  DFF ram_reg_426__7_ ( .D(n17216), .CP(wclk), .Q(ram[12975]) );
  DFF ram_reg_426__6_ ( .D(n17215), .CP(wclk), .Q(ram[12974]) );
  DFF ram_reg_426__5_ ( .D(n17214), .CP(wclk), .Q(ram[12973]) );
  DFF ram_reg_426__4_ ( .D(n17213), .CP(wclk), .Q(ram[12972]) );
  DFF ram_reg_426__3_ ( .D(n17212), .CP(wclk), .Q(ram[12971]) );
  DFF ram_reg_426__2_ ( .D(n17211), .CP(wclk), .Q(ram[12970]) );
  DFF ram_reg_426__1_ ( .D(n17210), .CP(wclk), .Q(ram[12969]) );
  DFF ram_reg_426__0_ ( .D(n17209), .CP(wclk), .Q(ram[12968]) );
  DFF ram_reg_430__7_ ( .D(n17184), .CP(wclk), .Q(ram[12943]) );
  DFF ram_reg_430__6_ ( .D(n17183), .CP(wclk), .Q(ram[12942]) );
  DFF ram_reg_430__5_ ( .D(n17182), .CP(wclk), .Q(ram[12941]) );
  DFF ram_reg_430__4_ ( .D(n17181), .CP(wclk), .Q(ram[12940]) );
  DFF ram_reg_430__3_ ( .D(n17180), .CP(wclk), .Q(ram[12939]) );
  DFF ram_reg_430__2_ ( .D(n17179), .CP(wclk), .Q(ram[12938]) );
  DFF ram_reg_430__1_ ( .D(n17178), .CP(wclk), .Q(ram[12937]) );
  DFF ram_reg_430__0_ ( .D(n17177), .CP(wclk), .Q(ram[12936]) );
  DFF ram_reg_434__7_ ( .D(n17152), .CP(wclk), .Q(ram[12911]) );
  DFF ram_reg_434__6_ ( .D(n17151), .CP(wclk), .Q(ram[12910]) );
  DFF ram_reg_434__5_ ( .D(n17150), .CP(wclk), .Q(ram[12909]) );
  DFF ram_reg_434__4_ ( .D(n17149), .CP(wclk), .Q(ram[12908]) );
  DFF ram_reg_434__3_ ( .D(n17148), .CP(wclk), .Q(ram[12907]) );
  DFF ram_reg_434__2_ ( .D(n17147), .CP(wclk), .Q(ram[12906]) );
  DFF ram_reg_434__1_ ( .D(n17146), .CP(wclk), .Q(ram[12905]) );
  DFF ram_reg_434__0_ ( .D(n17145), .CP(wclk), .Q(ram[12904]) );
  DFF ram_reg_442__7_ ( .D(n17088), .CP(wclk), .Q(ram[12847]) );
  DFF ram_reg_442__6_ ( .D(n17087), .CP(wclk), .Q(ram[12846]) );
  DFF ram_reg_442__5_ ( .D(n17086), .CP(wclk), .Q(ram[12845]) );
  DFF ram_reg_442__4_ ( .D(n17085), .CP(wclk), .Q(ram[12844]) );
  DFF ram_reg_442__3_ ( .D(n17084), .CP(wclk), .Q(ram[12843]) );
  DFF ram_reg_442__2_ ( .D(n17083), .CP(wclk), .Q(ram[12842]) );
  DFF ram_reg_442__1_ ( .D(n17082), .CP(wclk), .Q(ram[12841]) );
  DFF ram_reg_442__0_ ( .D(n17081), .CP(wclk), .Q(ram[12840]) );
  DFF ram_reg_446__7_ ( .D(n17056), .CP(wclk), .Q(ram[12815]) );
  DFF ram_reg_446__6_ ( .D(n17055), .CP(wclk), .Q(ram[12814]) );
  DFF ram_reg_446__5_ ( .D(n17054), .CP(wclk), .Q(ram[12813]) );
  DFF ram_reg_446__4_ ( .D(n17053), .CP(wclk), .Q(ram[12812]) );
  DFF ram_reg_446__3_ ( .D(n17052), .CP(wclk), .Q(ram[12811]) );
  DFF ram_reg_446__2_ ( .D(n17051), .CP(wclk), .Q(ram[12810]) );
  DFF ram_reg_446__1_ ( .D(n17050), .CP(wclk), .Q(ram[12809]) );
  DFF ram_reg_446__0_ ( .D(n17049), .CP(wclk), .Q(ram[12808]) );
  DFF ram_reg_458__7_ ( .D(n16960), .CP(wclk), .Q(ram[12719]) );
  DFF ram_reg_458__6_ ( .D(n16959), .CP(wclk), .Q(ram[12718]) );
  DFF ram_reg_458__5_ ( .D(n16958), .CP(wclk), .Q(ram[12717]) );
  DFF ram_reg_458__4_ ( .D(n16957), .CP(wclk), .Q(ram[12716]) );
  DFF ram_reg_458__3_ ( .D(n16956), .CP(wclk), .Q(ram[12715]) );
  DFF ram_reg_458__2_ ( .D(n16955), .CP(wclk), .Q(ram[12714]) );
  DFF ram_reg_458__1_ ( .D(n16954), .CP(wclk), .Q(ram[12713]) );
  DFF ram_reg_458__0_ ( .D(n16953), .CP(wclk), .Q(ram[12712]) );
  DFF ram_reg_490__7_ ( .D(n16704), .CP(wclk), .Q(ram[12463]) );
  DFF ram_reg_490__6_ ( .D(n16703), .CP(wclk), .Q(ram[12462]) );
  DFF ram_reg_490__5_ ( .D(n16702), .CP(wclk), .Q(ram[12461]) );
  DFF ram_reg_490__4_ ( .D(n16701), .CP(wclk), .Q(ram[12460]) );
  DFF ram_reg_490__3_ ( .D(n16700), .CP(wclk), .Q(ram[12459]) );
  DFF ram_reg_490__2_ ( .D(n16699), .CP(wclk), .Q(ram[12458]) );
  DFF ram_reg_490__1_ ( .D(n16698), .CP(wclk), .Q(ram[12457]) );
  DFF ram_reg_490__0_ ( .D(n16697), .CP(wclk), .Q(ram[12456]) );
  DFF ram_reg_494__7_ ( .D(n16672), .CP(wclk), .Q(ram[12431]) );
  DFF ram_reg_494__6_ ( .D(n16671), .CP(wclk), .Q(ram[12430]) );
  DFF ram_reg_494__5_ ( .D(n16670), .CP(wclk), .Q(ram[12429]) );
  DFF ram_reg_494__4_ ( .D(n16669), .CP(wclk), .Q(ram[12428]) );
  DFF ram_reg_494__3_ ( .D(n16668), .CP(wclk), .Q(ram[12427]) );
  DFF ram_reg_494__2_ ( .D(n16667), .CP(wclk), .Q(ram[12426]) );
  DFF ram_reg_494__1_ ( .D(n16666), .CP(wclk), .Q(ram[12425]) );
  DFF ram_reg_494__0_ ( .D(n16665), .CP(wclk), .Q(ram[12424]) );
  DFF ram_reg_506__7_ ( .D(n16576), .CP(wclk), .Q(ram[12335]) );
  DFF ram_reg_506__6_ ( .D(n16575), .CP(wclk), .Q(ram[12334]) );
  DFF ram_reg_506__5_ ( .D(n16574), .CP(wclk), .Q(ram[12333]) );
  DFF ram_reg_506__4_ ( .D(n16573), .CP(wclk), .Q(ram[12332]) );
  DFF ram_reg_506__3_ ( .D(n16572), .CP(wclk), .Q(ram[12331]) );
  DFF ram_reg_506__2_ ( .D(n16571), .CP(wclk), .Q(ram[12330]) );
  DFF ram_reg_506__1_ ( .D(n16570), .CP(wclk), .Q(ram[12329]) );
  DFF ram_reg_506__0_ ( .D(n16569), .CP(wclk), .Q(ram[12328]) );
  DFF ram_reg_510__7_ ( .D(n16544), .CP(wclk), .Q(ram[12303]) );
  DFF ram_reg_510__6_ ( .D(n16543), .CP(wclk), .Q(ram[12302]) );
  DFF ram_reg_510__5_ ( .D(n16542), .CP(wclk), .Q(ram[12301]) );
  DFF ram_reg_510__4_ ( .D(n16541), .CP(wclk), .Q(ram[12300]) );
  DFF ram_reg_510__3_ ( .D(n16540), .CP(wclk), .Q(ram[12299]) );
  DFF ram_reg_510__2_ ( .D(n16539), .CP(wclk), .Q(ram[12298]) );
  DFF ram_reg_510__1_ ( .D(n16538), .CP(wclk), .Q(ram[12297]) );
  DFF ram_reg_510__0_ ( .D(n16537), .CP(wclk), .Q(ram[12296]) );
  DFF ram_reg_522__7_ ( .D(n16448), .CP(wclk), .Q(ram[12207]) );
  DFF ram_reg_522__6_ ( .D(n16447), .CP(wclk), .Q(ram[12206]) );
  DFF ram_reg_522__5_ ( .D(n16446), .CP(wclk), .Q(ram[12205]) );
  DFF ram_reg_522__4_ ( .D(n16445), .CP(wclk), .Q(ram[12204]) );
  DFF ram_reg_522__3_ ( .D(n16444), .CP(wclk), .Q(ram[12203]) );
  DFF ram_reg_522__2_ ( .D(n16443), .CP(wclk), .Q(ram[12202]) );
  DFF ram_reg_522__1_ ( .D(n16442), .CP(wclk), .Q(ram[12201]) );
  DFF ram_reg_522__0_ ( .D(n16441), .CP(wclk), .Q(ram[12200]) );
  DFF ram_reg_554__7_ ( .D(n16192), .CP(wclk), .Q(ram[11951]) );
  DFF ram_reg_554__6_ ( .D(n16191), .CP(wclk), .Q(ram[11950]) );
  DFF ram_reg_554__5_ ( .D(n16190), .CP(wclk), .Q(ram[11949]) );
  DFF ram_reg_554__4_ ( .D(n16189), .CP(wclk), .Q(ram[11948]) );
  DFF ram_reg_554__3_ ( .D(n16188), .CP(wclk), .Q(ram[11947]) );
  DFF ram_reg_554__2_ ( .D(n16187), .CP(wclk), .Q(ram[11946]) );
  DFF ram_reg_554__1_ ( .D(n16186), .CP(wclk), .Q(ram[11945]) );
  DFF ram_reg_554__0_ ( .D(n16185), .CP(wclk), .Q(ram[11944]) );
  DFF ram_reg_558__7_ ( .D(n16160), .CP(wclk), .Q(ram[11919]) );
  DFF ram_reg_558__6_ ( .D(n16159), .CP(wclk), .Q(ram[11918]) );
  DFF ram_reg_558__5_ ( .D(n16158), .CP(wclk), .Q(ram[11917]) );
  DFF ram_reg_558__4_ ( .D(n16157), .CP(wclk), .Q(ram[11916]) );
  DFF ram_reg_558__3_ ( .D(n16156), .CP(wclk), .Q(ram[11915]) );
  DFF ram_reg_558__2_ ( .D(n16155), .CP(wclk), .Q(ram[11914]) );
  DFF ram_reg_558__1_ ( .D(n16154), .CP(wclk), .Q(ram[11913]) );
  DFF ram_reg_558__0_ ( .D(n16153), .CP(wclk), .Q(ram[11912]) );
  DFF ram_reg_570__7_ ( .D(n16064), .CP(wclk), .Q(ram[11823]) );
  DFF ram_reg_570__6_ ( .D(n16063), .CP(wclk), .Q(ram[11822]) );
  DFF ram_reg_570__5_ ( .D(n16062), .CP(wclk), .Q(ram[11821]) );
  DFF ram_reg_570__4_ ( .D(n16061), .CP(wclk), .Q(ram[11820]) );
  DFF ram_reg_570__3_ ( .D(n16060), .CP(wclk), .Q(ram[11819]) );
  DFF ram_reg_570__2_ ( .D(n16059), .CP(wclk), .Q(ram[11818]) );
  DFF ram_reg_570__1_ ( .D(n16058), .CP(wclk), .Q(ram[11817]) );
  DFF ram_reg_570__0_ ( .D(n16057), .CP(wclk), .Q(ram[11816]) );
  DFF ram_reg_574__7_ ( .D(n16032), .CP(wclk), .Q(ram[11791]) );
  DFF ram_reg_574__6_ ( .D(n16031), .CP(wclk), .Q(ram[11790]) );
  DFF ram_reg_574__5_ ( .D(n16030), .CP(wclk), .Q(ram[11789]) );
  DFF ram_reg_574__4_ ( .D(n16029), .CP(wclk), .Q(ram[11788]) );
  DFF ram_reg_574__3_ ( .D(n16028), .CP(wclk), .Q(ram[11787]) );
  DFF ram_reg_574__2_ ( .D(n16027), .CP(wclk), .Q(ram[11786]) );
  DFF ram_reg_574__1_ ( .D(n16026), .CP(wclk), .Q(ram[11785]) );
  DFF ram_reg_574__0_ ( .D(n16025), .CP(wclk), .Q(ram[11784]) );
  DFF ram_reg_642__7_ ( .D(n15488), .CP(wclk), .Q(ram[11247]) );
  DFF ram_reg_642__6_ ( .D(n15487), .CP(wclk), .Q(ram[11246]) );
  DFF ram_reg_642__5_ ( .D(n15486), .CP(wclk), .Q(ram[11245]) );
  DFF ram_reg_642__4_ ( .D(n15485), .CP(wclk), .Q(ram[11244]) );
  DFF ram_reg_642__3_ ( .D(n15484), .CP(wclk), .Q(ram[11243]) );
  DFF ram_reg_642__2_ ( .D(n15483), .CP(wclk), .Q(ram[11242]) );
  DFF ram_reg_642__1_ ( .D(n15482), .CP(wclk), .Q(ram[11241]) );
  DFF ram_reg_642__0_ ( .D(n15481), .CP(wclk), .Q(ram[11240]) );
  DFF ram_reg_650__7_ ( .D(n15424), .CP(wclk), .Q(ram[11183]) );
  DFF ram_reg_650__6_ ( .D(n15423), .CP(wclk), .Q(ram[11182]) );
  DFF ram_reg_650__5_ ( .D(n15422), .CP(wclk), .Q(ram[11181]) );
  DFF ram_reg_650__4_ ( .D(n15421), .CP(wclk), .Q(ram[11180]) );
  DFF ram_reg_650__3_ ( .D(n15420), .CP(wclk), .Q(ram[11179]) );
  DFF ram_reg_650__2_ ( .D(n15419), .CP(wclk), .Q(ram[11178]) );
  DFF ram_reg_650__1_ ( .D(n15418), .CP(wclk), .Q(ram[11177]) );
  DFF ram_reg_650__0_ ( .D(n15417), .CP(wclk), .Q(ram[11176]) );
  DFF ram_reg_654__7_ ( .D(n15392), .CP(wclk), .Q(ram[11151]) );
  DFF ram_reg_654__6_ ( .D(n15391), .CP(wclk), .Q(ram[11150]) );
  DFF ram_reg_654__5_ ( .D(n15390), .CP(wclk), .Q(ram[11149]) );
  DFF ram_reg_654__4_ ( .D(n15389), .CP(wclk), .Q(ram[11148]) );
  DFF ram_reg_654__3_ ( .D(n15388), .CP(wclk), .Q(ram[11147]) );
  DFF ram_reg_654__2_ ( .D(n15387), .CP(wclk), .Q(ram[11146]) );
  DFF ram_reg_654__1_ ( .D(n15386), .CP(wclk), .Q(ram[11145]) );
  DFF ram_reg_654__0_ ( .D(n15385), .CP(wclk), .Q(ram[11144]) );
  DFF ram_reg_666__7_ ( .D(n15296), .CP(wclk), .Q(ram[11055]) );
  DFF ram_reg_666__6_ ( .D(n15295), .CP(wclk), .Q(ram[11054]) );
  DFF ram_reg_666__5_ ( .D(n15294), .CP(wclk), .Q(ram[11053]) );
  DFF ram_reg_666__4_ ( .D(n15293), .CP(wclk), .Q(ram[11052]) );
  DFF ram_reg_666__3_ ( .D(n15292), .CP(wclk), .Q(ram[11051]) );
  DFF ram_reg_666__2_ ( .D(n15291), .CP(wclk), .Q(ram[11050]) );
  DFF ram_reg_666__1_ ( .D(n15290), .CP(wclk), .Q(ram[11049]) );
  DFF ram_reg_666__0_ ( .D(n15289), .CP(wclk), .Q(ram[11048]) );
  DFF ram_reg_670__7_ ( .D(n15264), .CP(wclk), .Q(ram[11023]) );
  DFF ram_reg_670__6_ ( .D(n15263), .CP(wclk), .Q(ram[11022]) );
  DFF ram_reg_670__5_ ( .D(n15262), .CP(wclk), .Q(ram[11021]) );
  DFF ram_reg_670__4_ ( .D(n15261), .CP(wclk), .Q(ram[11020]) );
  DFF ram_reg_670__3_ ( .D(n15260), .CP(wclk), .Q(ram[11019]) );
  DFF ram_reg_670__2_ ( .D(n15259), .CP(wclk), .Q(ram[11018]) );
  DFF ram_reg_670__1_ ( .D(n15258), .CP(wclk), .Q(ram[11017]) );
  DFF ram_reg_670__0_ ( .D(n15257), .CP(wclk), .Q(ram[11016]) );
  DFF ram_reg_674__7_ ( .D(n15232), .CP(wclk), .Q(ram[10991]) );
  DFF ram_reg_674__6_ ( .D(n15231), .CP(wclk), .Q(ram[10990]) );
  DFF ram_reg_674__5_ ( .D(n15230), .CP(wclk), .Q(ram[10989]) );
  DFF ram_reg_674__4_ ( .D(n15229), .CP(wclk), .Q(ram[10988]) );
  DFF ram_reg_674__3_ ( .D(n15228), .CP(wclk), .Q(ram[10987]) );
  DFF ram_reg_674__2_ ( .D(n15227), .CP(wclk), .Q(ram[10986]) );
  DFF ram_reg_674__1_ ( .D(n15226), .CP(wclk), .Q(ram[10985]) );
  DFF ram_reg_674__0_ ( .D(n15225), .CP(wclk), .Q(ram[10984]) );
  DFF ram_reg_682__7_ ( .D(n15168), .CP(wclk), .Q(ram[10927]) );
  DFF ram_reg_682__6_ ( .D(n15167), .CP(wclk), .Q(ram[10926]) );
  DFF ram_reg_682__5_ ( .D(n15166), .CP(wclk), .Q(ram[10925]) );
  DFF ram_reg_682__4_ ( .D(n15165), .CP(wclk), .Q(ram[10924]) );
  DFF ram_reg_682__3_ ( .D(n15164), .CP(wclk), .Q(ram[10923]) );
  DFF ram_reg_682__2_ ( .D(n15163), .CP(wclk), .Q(ram[10922]) );
  DFF ram_reg_682__1_ ( .D(n15162), .CP(wclk), .Q(ram[10921]) );
  DFF ram_reg_682__0_ ( .D(n15161), .CP(wclk), .Q(ram[10920]) );
  DFF ram_reg_686__7_ ( .D(n15136), .CP(wclk), .Q(ram[10895]) );
  DFF ram_reg_686__6_ ( .D(n15135), .CP(wclk), .Q(ram[10894]) );
  DFF ram_reg_686__5_ ( .D(n15134), .CP(wclk), .Q(ram[10893]) );
  DFF ram_reg_686__4_ ( .D(n15133), .CP(wclk), .Q(ram[10892]) );
  DFF ram_reg_686__3_ ( .D(n15132), .CP(wclk), .Q(ram[10891]) );
  DFF ram_reg_686__2_ ( .D(n15131), .CP(wclk), .Q(ram[10890]) );
  DFF ram_reg_686__1_ ( .D(n15130), .CP(wclk), .Q(ram[10889]) );
  DFF ram_reg_686__0_ ( .D(n15129), .CP(wclk), .Q(ram[10888]) );
  DFF ram_reg_690__7_ ( .D(n15104), .CP(wclk), .Q(ram[10863]) );
  DFF ram_reg_690__6_ ( .D(n15103), .CP(wclk), .Q(ram[10862]) );
  DFF ram_reg_690__5_ ( .D(n15102), .CP(wclk), .Q(ram[10861]) );
  DFF ram_reg_690__4_ ( .D(n15101), .CP(wclk), .Q(ram[10860]) );
  DFF ram_reg_690__3_ ( .D(n15100), .CP(wclk), .Q(ram[10859]) );
  DFF ram_reg_690__2_ ( .D(n15099), .CP(wclk), .Q(ram[10858]) );
  DFF ram_reg_690__1_ ( .D(n15098), .CP(wclk), .Q(ram[10857]) );
  DFF ram_reg_690__0_ ( .D(n15097), .CP(wclk), .Q(ram[10856]) );
  DFF ram_reg_698__7_ ( .D(n15040), .CP(wclk), .Q(ram[10799]) );
  DFF ram_reg_698__6_ ( .D(n15039), .CP(wclk), .Q(ram[10798]) );
  DFF ram_reg_698__5_ ( .D(n15038), .CP(wclk), .Q(ram[10797]) );
  DFF ram_reg_698__4_ ( .D(n15037), .CP(wclk), .Q(ram[10796]) );
  DFF ram_reg_698__3_ ( .D(n15036), .CP(wclk), .Q(ram[10795]) );
  DFF ram_reg_698__2_ ( .D(n15035), .CP(wclk), .Q(ram[10794]) );
  DFF ram_reg_698__1_ ( .D(n15034), .CP(wclk), .Q(ram[10793]) );
  DFF ram_reg_698__0_ ( .D(n15033), .CP(wclk), .Q(ram[10792]) );
  DFF ram_reg_702__7_ ( .D(n15008), .CP(wclk), .Q(ram[10767]) );
  DFF ram_reg_702__6_ ( .D(n15007), .CP(wclk), .Q(ram[10766]) );
  DFF ram_reg_702__5_ ( .D(n15006), .CP(wclk), .Q(ram[10765]) );
  DFF ram_reg_702__4_ ( .D(n15005), .CP(wclk), .Q(ram[10764]) );
  DFF ram_reg_702__3_ ( .D(n15004), .CP(wclk), .Q(ram[10763]) );
  DFF ram_reg_702__2_ ( .D(n15003), .CP(wclk), .Q(ram[10762]) );
  DFF ram_reg_702__1_ ( .D(n15002), .CP(wclk), .Q(ram[10761]) );
  DFF ram_reg_702__0_ ( .D(n15001), .CP(wclk), .Q(ram[10760]) );
  DFF ram_reg_714__7_ ( .D(n14912), .CP(wclk), .Q(ram[10671]) );
  DFF ram_reg_714__6_ ( .D(n14911), .CP(wclk), .Q(ram[10670]) );
  DFF ram_reg_714__5_ ( .D(n14910), .CP(wclk), .Q(ram[10669]) );
  DFF ram_reg_714__4_ ( .D(n14909), .CP(wclk), .Q(ram[10668]) );
  DFF ram_reg_714__3_ ( .D(n14908), .CP(wclk), .Q(ram[10667]) );
  DFF ram_reg_714__2_ ( .D(n14907), .CP(wclk), .Q(ram[10666]) );
  DFF ram_reg_714__1_ ( .D(n14906), .CP(wclk), .Q(ram[10665]) );
  DFF ram_reg_714__0_ ( .D(n14905), .CP(wclk), .Q(ram[10664]) );
  DFF ram_reg_718__7_ ( .D(n14880), .CP(wclk), .Q(ram[10639]) );
  DFF ram_reg_718__6_ ( .D(n14879), .CP(wclk), .Q(ram[10638]) );
  DFF ram_reg_718__5_ ( .D(n14878), .CP(wclk), .Q(ram[10637]) );
  DFF ram_reg_718__4_ ( .D(n14877), .CP(wclk), .Q(ram[10636]) );
  DFF ram_reg_718__3_ ( .D(n14876), .CP(wclk), .Q(ram[10635]) );
  DFF ram_reg_718__2_ ( .D(n14875), .CP(wclk), .Q(ram[10634]) );
  DFF ram_reg_718__1_ ( .D(n14874), .CP(wclk), .Q(ram[10633]) );
  DFF ram_reg_718__0_ ( .D(n14873), .CP(wclk), .Q(ram[10632]) );
  DFF ram_reg_730__7_ ( .D(n14784), .CP(wclk), .Q(ram[10543]) );
  DFF ram_reg_730__6_ ( .D(n14783), .CP(wclk), .Q(ram[10542]) );
  DFF ram_reg_730__5_ ( .D(n14782), .CP(wclk), .Q(ram[10541]) );
  DFF ram_reg_730__4_ ( .D(n14781), .CP(wclk), .Q(ram[10540]) );
  DFF ram_reg_730__3_ ( .D(n14780), .CP(wclk), .Q(ram[10539]) );
  DFF ram_reg_730__2_ ( .D(n14779), .CP(wclk), .Q(ram[10538]) );
  DFF ram_reg_730__1_ ( .D(n14778), .CP(wclk), .Q(ram[10537]) );
  DFF ram_reg_730__0_ ( .D(n14777), .CP(wclk), .Q(ram[10536]) );
  DFF ram_reg_738__7_ ( .D(n14720), .CP(wclk), .Q(ram[10479]) );
  DFF ram_reg_738__6_ ( .D(n14719), .CP(wclk), .Q(ram[10478]) );
  DFF ram_reg_738__5_ ( .D(n14718), .CP(wclk), .Q(ram[10477]) );
  DFF ram_reg_738__4_ ( .D(n14717), .CP(wclk), .Q(ram[10476]) );
  DFF ram_reg_738__3_ ( .D(n14716), .CP(wclk), .Q(ram[10475]) );
  DFF ram_reg_738__2_ ( .D(n14715), .CP(wclk), .Q(ram[10474]) );
  DFF ram_reg_738__1_ ( .D(n14714), .CP(wclk), .Q(ram[10473]) );
  DFF ram_reg_738__0_ ( .D(n14713), .CP(wclk), .Q(ram[10472]) );
  DFF ram_reg_746__7_ ( .D(n14656), .CP(wclk), .Q(ram[10415]) );
  DFF ram_reg_746__6_ ( .D(n14655), .CP(wclk), .Q(ram[10414]) );
  DFF ram_reg_746__5_ ( .D(n14654), .CP(wclk), .Q(ram[10413]) );
  DFF ram_reg_746__4_ ( .D(n14653), .CP(wclk), .Q(ram[10412]) );
  DFF ram_reg_746__3_ ( .D(n14652), .CP(wclk), .Q(ram[10411]) );
  DFF ram_reg_746__2_ ( .D(n14651), .CP(wclk), .Q(ram[10410]) );
  DFF ram_reg_746__1_ ( .D(n14650), .CP(wclk), .Q(ram[10409]) );
  DFF ram_reg_746__0_ ( .D(n14649), .CP(wclk), .Q(ram[10408]) );
  DFF ram_reg_750__7_ ( .D(n14624), .CP(wclk), .Q(ram[10383]) );
  DFF ram_reg_750__6_ ( .D(n14623), .CP(wclk), .Q(ram[10382]) );
  DFF ram_reg_750__5_ ( .D(n14622), .CP(wclk), .Q(ram[10381]) );
  DFF ram_reg_750__4_ ( .D(n14621), .CP(wclk), .Q(ram[10380]) );
  DFF ram_reg_750__3_ ( .D(n14620), .CP(wclk), .Q(ram[10379]) );
  DFF ram_reg_750__2_ ( .D(n14619), .CP(wclk), .Q(ram[10378]) );
  DFF ram_reg_750__1_ ( .D(n14618), .CP(wclk), .Q(ram[10377]) );
  DFF ram_reg_750__0_ ( .D(n14617), .CP(wclk), .Q(ram[10376]) );
  DFF ram_reg_754__7_ ( .D(n14592), .CP(wclk), .Q(ram[10351]) );
  DFF ram_reg_754__6_ ( .D(n14591), .CP(wclk), .Q(ram[10350]) );
  DFF ram_reg_754__5_ ( .D(n14590), .CP(wclk), .Q(ram[10349]) );
  DFF ram_reg_754__4_ ( .D(n14589), .CP(wclk), .Q(ram[10348]) );
  DFF ram_reg_754__3_ ( .D(n14588), .CP(wclk), .Q(ram[10347]) );
  DFF ram_reg_754__2_ ( .D(n14587), .CP(wclk), .Q(ram[10346]) );
  DFF ram_reg_754__1_ ( .D(n14586), .CP(wclk), .Q(ram[10345]) );
  DFF ram_reg_754__0_ ( .D(n14585), .CP(wclk), .Q(ram[10344]) );
  DFF ram_reg_762__7_ ( .D(n14528), .CP(wclk), .Q(ram[10287]) );
  DFF ram_reg_762__6_ ( .D(n14527), .CP(wclk), .Q(ram[10286]) );
  DFF ram_reg_762__5_ ( .D(n14526), .CP(wclk), .Q(ram[10285]) );
  DFF ram_reg_762__4_ ( .D(n14525), .CP(wclk), .Q(ram[10284]) );
  DFF ram_reg_762__3_ ( .D(n14524), .CP(wclk), .Q(ram[10283]) );
  DFF ram_reg_762__2_ ( .D(n14523), .CP(wclk), .Q(ram[10282]) );
  DFF ram_reg_762__1_ ( .D(n14522), .CP(wclk), .Q(ram[10281]) );
  DFF ram_reg_762__0_ ( .D(n14521), .CP(wclk), .Q(ram[10280]) );
  DFF ram_reg_766__7_ ( .D(n14496), .CP(wclk), .Q(ram[10255]) );
  DFF ram_reg_766__6_ ( .D(n14495), .CP(wclk), .Q(ram[10254]) );
  DFF ram_reg_766__5_ ( .D(n14494), .CP(wclk), .Q(ram[10253]) );
  DFF ram_reg_766__4_ ( .D(n14493), .CP(wclk), .Q(ram[10252]) );
  DFF ram_reg_766__3_ ( .D(n14492), .CP(wclk), .Q(ram[10251]) );
  DFF ram_reg_766__2_ ( .D(n14491), .CP(wclk), .Q(ram[10250]) );
  DFF ram_reg_766__1_ ( .D(n14490), .CP(wclk), .Q(ram[10249]) );
  DFF ram_reg_766__0_ ( .D(n14489), .CP(wclk), .Q(ram[10248]) );
  DFF ram_reg_778__7_ ( .D(n14400), .CP(wclk), .Q(ram[10159]) );
  DFF ram_reg_778__6_ ( .D(n14399), .CP(wclk), .Q(ram[10158]) );
  DFF ram_reg_778__5_ ( .D(n14398), .CP(wclk), .Q(ram[10157]) );
  DFF ram_reg_778__4_ ( .D(n14397), .CP(wclk), .Q(ram[10156]) );
  DFF ram_reg_778__3_ ( .D(n14396), .CP(wclk), .Q(ram[10155]) );
  DFF ram_reg_778__2_ ( .D(n14395), .CP(wclk), .Q(ram[10154]) );
  DFF ram_reg_778__1_ ( .D(n14394), .CP(wclk), .Q(ram[10153]) );
  DFF ram_reg_778__0_ ( .D(n14393), .CP(wclk), .Q(ram[10152]) );
  DFF ram_reg_810__7_ ( .D(n14144), .CP(wclk), .Q(ram[9903]) );
  DFF ram_reg_810__6_ ( .D(n14143), .CP(wclk), .Q(ram[9902]) );
  DFF ram_reg_810__5_ ( .D(n14142), .CP(wclk), .Q(ram[9901]) );
  DFF ram_reg_810__4_ ( .D(n14141), .CP(wclk), .Q(ram[9900]) );
  DFF ram_reg_810__3_ ( .D(n14140), .CP(wclk), .Q(ram[9899]) );
  DFF ram_reg_810__2_ ( .D(n14139), .CP(wclk), .Q(ram[9898]) );
  DFF ram_reg_810__1_ ( .D(n14138), .CP(wclk), .Q(ram[9897]) );
  DFF ram_reg_810__0_ ( .D(n14137), .CP(wclk), .Q(ram[9896]) );
  DFF ram_reg_814__7_ ( .D(n14112), .CP(wclk), .Q(ram[9871]) );
  DFF ram_reg_814__6_ ( .D(n14111), .CP(wclk), .Q(ram[9870]) );
  DFF ram_reg_814__5_ ( .D(n14110), .CP(wclk), .Q(ram[9869]) );
  DFF ram_reg_814__4_ ( .D(n14109), .CP(wclk), .Q(ram[9868]) );
  DFF ram_reg_814__3_ ( .D(n14108), .CP(wclk), .Q(ram[9867]) );
  DFF ram_reg_814__2_ ( .D(n14107), .CP(wclk), .Q(ram[9866]) );
  DFF ram_reg_814__1_ ( .D(n14106), .CP(wclk), .Q(ram[9865]) );
  DFF ram_reg_814__0_ ( .D(n14105), .CP(wclk), .Q(ram[9864]) );
  DFF ram_reg_826__7_ ( .D(n14016), .CP(wclk), .Q(ram[9775]) );
  DFF ram_reg_826__6_ ( .D(n14015), .CP(wclk), .Q(ram[9774]) );
  DFF ram_reg_826__5_ ( .D(n14014), .CP(wclk), .Q(ram[9773]) );
  DFF ram_reg_826__4_ ( .D(n14013), .CP(wclk), .Q(ram[9772]) );
  DFF ram_reg_826__3_ ( .D(n14012), .CP(wclk), .Q(ram[9771]) );
  DFF ram_reg_826__2_ ( .D(n14011), .CP(wclk), .Q(ram[9770]) );
  DFF ram_reg_826__1_ ( .D(n14010), .CP(wclk), .Q(ram[9769]) );
  DFF ram_reg_826__0_ ( .D(n14009), .CP(wclk), .Q(ram[9768]) );
  DFF ram_reg_830__7_ ( .D(n13984), .CP(wclk), .Q(ram[9743]) );
  DFF ram_reg_830__6_ ( .D(n13983), .CP(wclk), .Q(ram[9742]) );
  DFF ram_reg_830__5_ ( .D(n13982), .CP(wclk), .Q(ram[9741]) );
  DFF ram_reg_830__4_ ( .D(n13981), .CP(wclk), .Q(ram[9740]) );
  DFF ram_reg_830__3_ ( .D(n13980), .CP(wclk), .Q(ram[9739]) );
  DFF ram_reg_830__2_ ( .D(n13979), .CP(wclk), .Q(ram[9738]) );
  DFF ram_reg_830__1_ ( .D(n13978), .CP(wclk), .Q(ram[9737]) );
  DFF ram_reg_830__0_ ( .D(n13977), .CP(wclk), .Q(ram[9736]) );
  DFF ram_reg_898__7_ ( .D(n13440), .CP(wclk), .Q(ram[9199]) );
  DFF ram_reg_898__6_ ( .D(n13439), .CP(wclk), .Q(ram[9198]) );
  DFF ram_reg_898__5_ ( .D(n13438), .CP(wclk), .Q(ram[9197]) );
  DFF ram_reg_898__4_ ( .D(n13437), .CP(wclk), .Q(ram[9196]) );
  DFF ram_reg_898__3_ ( .D(n13436), .CP(wclk), .Q(ram[9195]) );
  DFF ram_reg_898__2_ ( .D(n13435), .CP(wclk), .Q(ram[9194]) );
  DFF ram_reg_898__1_ ( .D(n13434), .CP(wclk), .Q(ram[9193]) );
  DFF ram_reg_898__0_ ( .D(n13433), .CP(wclk), .Q(ram[9192]) );
  DFF ram_reg_906__7_ ( .D(n13376), .CP(wclk), .Q(ram[9135]) );
  DFF ram_reg_906__6_ ( .D(n13375), .CP(wclk), .Q(ram[9134]) );
  DFF ram_reg_906__5_ ( .D(n13374), .CP(wclk), .Q(ram[9133]) );
  DFF ram_reg_906__4_ ( .D(n13373), .CP(wclk), .Q(ram[9132]) );
  DFF ram_reg_906__3_ ( .D(n13372), .CP(wclk), .Q(ram[9131]) );
  DFF ram_reg_906__2_ ( .D(n13371), .CP(wclk), .Q(ram[9130]) );
  DFF ram_reg_906__1_ ( .D(n13370), .CP(wclk), .Q(ram[9129]) );
  DFF ram_reg_906__0_ ( .D(n13369), .CP(wclk), .Q(ram[9128]) );
  DFF ram_reg_910__7_ ( .D(n13344), .CP(wclk), .Q(ram[9103]) );
  DFF ram_reg_910__6_ ( .D(n13343), .CP(wclk), .Q(ram[9102]) );
  DFF ram_reg_910__5_ ( .D(n13342), .CP(wclk), .Q(ram[9101]) );
  DFF ram_reg_910__4_ ( .D(n13341), .CP(wclk), .Q(ram[9100]) );
  DFF ram_reg_910__3_ ( .D(n13340), .CP(wclk), .Q(ram[9099]) );
  DFF ram_reg_910__2_ ( .D(n13339), .CP(wclk), .Q(ram[9098]) );
  DFF ram_reg_910__1_ ( .D(n13338), .CP(wclk), .Q(ram[9097]) );
  DFF ram_reg_910__0_ ( .D(n13337), .CP(wclk), .Q(ram[9096]) );
  DFF ram_reg_922__7_ ( .D(n13248), .CP(wclk), .Q(ram[9007]) );
  DFF ram_reg_922__6_ ( .D(n13247), .CP(wclk), .Q(ram[9006]) );
  DFF ram_reg_922__5_ ( .D(n13246), .CP(wclk), .Q(ram[9005]) );
  DFF ram_reg_922__4_ ( .D(n13245), .CP(wclk), .Q(ram[9004]) );
  DFF ram_reg_922__3_ ( .D(n13244), .CP(wclk), .Q(ram[9003]) );
  DFF ram_reg_922__2_ ( .D(n13243), .CP(wclk), .Q(ram[9002]) );
  DFF ram_reg_922__1_ ( .D(n13242), .CP(wclk), .Q(ram[9001]) );
  DFF ram_reg_922__0_ ( .D(n13241), .CP(wclk), .Q(ram[9000]) );
  DFF ram_reg_926__7_ ( .D(n13216), .CP(wclk), .Q(ram[8975]) );
  DFF ram_reg_926__6_ ( .D(n13215), .CP(wclk), .Q(ram[8974]) );
  DFF ram_reg_926__5_ ( .D(n13214), .CP(wclk), .Q(ram[8973]) );
  DFF ram_reg_926__4_ ( .D(n13213), .CP(wclk), .Q(ram[8972]) );
  DFF ram_reg_926__3_ ( .D(n13212), .CP(wclk), .Q(ram[8971]) );
  DFF ram_reg_926__2_ ( .D(n13211), .CP(wclk), .Q(ram[8970]) );
  DFF ram_reg_926__1_ ( .D(n13210), .CP(wclk), .Q(ram[8969]) );
  DFF ram_reg_926__0_ ( .D(n13209), .CP(wclk), .Q(ram[8968]) );
  DFF ram_reg_930__7_ ( .D(n13184), .CP(wclk), .Q(ram[8943]) );
  DFF ram_reg_930__6_ ( .D(n13183), .CP(wclk), .Q(ram[8942]) );
  DFF ram_reg_930__5_ ( .D(n13182), .CP(wclk), .Q(ram[8941]) );
  DFF ram_reg_930__4_ ( .D(n13181), .CP(wclk), .Q(ram[8940]) );
  DFF ram_reg_930__3_ ( .D(n13180), .CP(wclk), .Q(ram[8939]) );
  DFF ram_reg_930__2_ ( .D(n13179), .CP(wclk), .Q(ram[8938]) );
  DFF ram_reg_930__1_ ( .D(n13178), .CP(wclk), .Q(ram[8937]) );
  DFF ram_reg_930__0_ ( .D(n13177), .CP(wclk), .Q(ram[8936]) );
  DFF ram_reg_938__7_ ( .D(n13120), .CP(wclk), .Q(ram[8879]) );
  DFF ram_reg_938__6_ ( .D(n13119), .CP(wclk), .Q(ram[8878]) );
  DFF ram_reg_938__5_ ( .D(n13118), .CP(wclk), .Q(ram[8877]) );
  DFF ram_reg_938__4_ ( .D(n13117), .CP(wclk), .Q(ram[8876]) );
  DFF ram_reg_938__3_ ( .D(n13116), .CP(wclk), .Q(ram[8875]) );
  DFF ram_reg_938__2_ ( .D(n13115), .CP(wclk), .Q(ram[8874]) );
  DFF ram_reg_938__1_ ( .D(n13114), .CP(wclk), .Q(ram[8873]) );
  DFF ram_reg_938__0_ ( .D(n13113), .CP(wclk), .Q(ram[8872]) );
  DFF ram_reg_942__7_ ( .D(n13088), .CP(wclk), .Q(ram[8847]) );
  DFF ram_reg_942__6_ ( .D(n13087), .CP(wclk), .Q(ram[8846]) );
  DFF ram_reg_942__5_ ( .D(n13086), .CP(wclk), .Q(ram[8845]) );
  DFF ram_reg_942__4_ ( .D(n13085), .CP(wclk), .Q(ram[8844]) );
  DFF ram_reg_942__3_ ( .D(n13084), .CP(wclk), .Q(ram[8843]) );
  DFF ram_reg_942__2_ ( .D(n13083), .CP(wclk), .Q(ram[8842]) );
  DFF ram_reg_942__1_ ( .D(n13082), .CP(wclk), .Q(ram[8841]) );
  DFF ram_reg_942__0_ ( .D(n13081), .CP(wclk), .Q(ram[8840]) );
  DFF ram_reg_946__7_ ( .D(n13056), .CP(wclk), .Q(ram[8815]) );
  DFF ram_reg_946__6_ ( .D(n13055), .CP(wclk), .Q(ram[8814]) );
  DFF ram_reg_946__5_ ( .D(n13054), .CP(wclk), .Q(ram[8813]) );
  DFF ram_reg_946__4_ ( .D(n13053), .CP(wclk), .Q(ram[8812]) );
  DFF ram_reg_946__3_ ( .D(n13052), .CP(wclk), .Q(ram[8811]) );
  DFF ram_reg_946__2_ ( .D(n13051), .CP(wclk), .Q(ram[8810]) );
  DFF ram_reg_946__1_ ( .D(n13050), .CP(wclk), .Q(ram[8809]) );
  DFF ram_reg_946__0_ ( .D(n13049), .CP(wclk), .Q(ram[8808]) );
  DFF ram_reg_954__7_ ( .D(n12992), .CP(wclk), .Q(ram[8751]) );
  DFF ram_reg_954__6_ ( .D(n12991), .CP(wclk), .Q(ram[8750]) );
  DFF ram_reg_954__5_ ( .D(n12990), .CP(wclk), .Q(ram[8749]) );
  DFF ram_reg_954__4_ ( .D(n12989), .CP(wclk), .Q(ram[8748]) );
  DFF ram_reg_954__3_ ( .D(n12988), .CP(wclk), .Q(ram[8747]) );
  DFF ram_reg_954__2_ ( .D(n12987), .CP(wclk), .Q(ram[8746]) );
  DFF ram_reg_954__1_ ( .D(n12986), .CP(wclk), .Q(ram[8745]) );
  DFF ram_reg_954__0_ ( .D(n12985), .CP(wclk), .Q(ram[8744]) );
  DFF ram_reg_958__7_ ( .D(n12960), .CP(wclk), .Q(ram[8719]) );
  DFF ram_reg_958__6_ ( .D(n12959), .CP(wclk), .Q(ram[8718]) );
  DFF ram_reg_958__5_ ( .D(n12958), .CP(wclk), .Q(ram[8717]) );
  DFF ram_reg_958__4_ ( .D(n12957), .CP(wclk), .Q(ram[8716]) );
  DFF ram_reg_958__3_ ( .D(n12956), .CP(wclk), .Q(ram[8715]) );
  DFF ram_reg_958__2_ ( .D(n12955), .CP(wclk), .Q(ram[8714]) );
  DFF ram_reg_958__1_ ( .D(n12954), .CP(wclk), .Q(ram[8713]) );
  DFF ram_reg_958__0_ ( .D(n12953), .CP(wclk), .Q(ram[8712]) );
  DFF ram_reg_970__7_ ( .D(n12864), .CP(wclk), .Q(ram[8623]) );
  DFF ram_reg_970__6_ ( .D(n12863), .CP(wclk), .Q(ram[8622]) );
  DFF ram_reg_970__5_ ( .D(n12862), .CP(wclk), .Q(ram[8621]) );
  DFF ram_reg_970__4_ ( .D(n12861), .CP(wclk), .Q(ram[8620]) );
  DFF ram_reg_970__3_ ( .D(n12860), .CP(wclk), .Q(ram[8619]) );
  DFF ram_reg_970__2_ ( .D(n12859), .CP(wclk), .Q(ram[8618]) );
  DFF ram_reg_970__1_ ( .D(n12858), .CP(wclk), .Q(ram[8617]) );
  DFF ram_reg_970__0_ ( .D(n12857), .CP(wclk), .Q(ram[8616]) );
  DFF ram_reg_974__7_ ( .D(n12832), .CP(wclk), .Q(ram[8591]) );
  DFF ram_reg_974__6_ ( .D(n12831), .CP(wclk), .Q(ram[8590]) );
  DFF ram_reg_974__5_ ( .D(n12830), .CP(wclk), .Q(ram[8589]) );
  DFF ram_reg_974__4_ ( .D(n12829), .CP(wclk), .Q(ram[8588]) );
  DFF ram_reg_974__3_ ( .D(n12828), .CP(wclk), .Q(ram[8587]) );
  DFF ram_reg_974__2_ ( .D(n12827), .CP(wclk), .Q(ram[8586]) );
  DFF ram_reg_974__1_ ( .D(n12826), .CP(wclk), .Q(ram[8585]) );
  DFF ram_reg_974__0_ ( .D(n12825), .CP(wclk), .Q(ram[8584]) );
  DFF ram_reg_986__7_ ( .D(n12736), .CP(wclk), .Q(ram[8495]) );
  DFF ram_reg_986__6_ ( .D(n12735), .CP(wclk), .Q(ram[8494]) );
  DFF ram_reg_986__5_ ( .D(n12734), .CP(wclk), .Q(ram[8493]) );
  DFF ram_reg_986__4_ ( .D(n12733), .CP(wclk), .Q(ram[8492]) );
  DFF ram_reg_986__3_ ( .D(n12732), .CP(wclk), .Q(ram[8491]) );
  DFF ram_reg_986__2_ ( .D(n12731), .CP(wclk), .Q(ram[8490]) );
  DFF ram_reg_986__1_ ( .D(n12730), .CP(wclk), .Q(ram[8489]) );
  DFF ram_reg_986__0_ ( .D(n12729), .CP(wclk), .Q(ram[8488]) );
  DFF ram_reg_990__7_ ( .D(n12704), .CP(wclk), .Q(ram[8463]) );
  DFF ram_reg_990__6_ ( .D(n12703), .CP(wclk), .Q(ram[8462]) );
  DFF ram_reg_990__5_ ( .D(n12702), .CP(wclk), .Q(ram[8461]) );
  DFF ram_reg_990__4_ ( .D(n12701), .CP(wclk), .Q(ram[8460]) );
  DFF ram_reg_990__3_ ( .D(n12700), .CP(wclk), .Q(ram[8459]) );
  DFF ram_reg_990__2_ ( .D(n12699), .CP(wclk), .Q(ram[8458]) );
  DFF ram_reg_990__1_ ( .D(n12698), .CP(wclk), .Q(ram[8457]) );
  DFF ram_reg_990__0_ ( .D(n12697), .CP(wclk), .Q(ram[8456]) );
  DFF ram_reg_994__7_ ( .D(n12672), .CP(wclk), .Q(ram[8431]) );
  DFF ram_reg_994__6_ ( .D(n12671), .CP(wclk), .Q(ram[8430]) );
  DFF ram_reg_994__5_ ( .D(n12670), .CP(wclk), .Q(ram[8429]) );
  DFF ram_reg_994__4_ ( .D(n12669), .CP(wclk), .Q(ram[8428]) );
  DFF ram_reg_994__3_ ( .D(n12668), .CP(wclk), .Q(ram[8427]) );
  DFF ram_reg_994__2_ ( .D(n12667), .CP(wclk), .Q(ram[8426]) );
  DFF ram_reg_994__1_ ( .D(n12666), .CP(wclk), .Q(ram[8425]) );
  DFF ram_reg_994__0_ ( .D(n12665), .CP(wclk), .Q(ram[8424]) );
  DFF ram_reg_1002__7_ ( .D(n12608), .CP(wclk), .Q(ram[8367]) );
  DFF ram_reg_1002__6_ ( .D(n12607), .CP(wclk), .Q(ram[8366]) );
  DFF ram_reg_1002__5_ ( .D(n12606), .CP(wclk), .Q(ram[8365]) );
  DFF ram_reg_1002__4_ ( .D(n12605), .CP(wclk), .Q(ram[8364]) );
  DFF ram_reg_1002__3_ ( .D(n12604), .CP(wclk), .Q(ram[8363]) );
  DFF ram_reg_1002__2_ ( .D(n12603), .CP(wclk), .Q(ram[8362]) );
  DFF ram_reg_1002__1_ ( .D(n12602), .CP(wclk), .Q(ram[8361]) );
  DFF ram_reg_1002__0_ ( .D(n12601), .CP(wclk), .Q(ram[8360]) );
  DFF ram_reg_1006__7_ ( .D(n12576), .CP(wclk), .Q(ram[8335]) );
  DFF ram_reg_1006__6_ ( .D(n12575), .CP(wclk), .Q(ram[8334]) );
  DFF ram_reg_1006__5_ ( .D(n12574), .CP(wclk), .Q(ram[8333]) );
  DFF ram_reg_1006__4_ ( .D(n12573), .CP(wclk), .Q(ram[8332]) );
  DFF ram_reg_1006__3_ ( .D(n12572), .CP(wclk), .Q(ram[8331]) );
  DFF ram_reg_1006__2_ ( .D(n12571), .CP(wclk), .Q(ram[8330]) );
  DFF ram_reg_1006__1_ ( .D(n12570), .CP(wclk), .Q(ram[8329]) );
  DFF ram_reg_1006__0_ ( .D(n12569), .CP(wclk), .Q(ram[8328]) );
  DFF ram_reg_1010__7_ ( .D(n12544), .CP(wclk), .Q(ram[8303]) );
  DFF ram_reg_1010__6_ ( .D(n12543), .CP(wclk), .Q(ram[8302]) );
  DFF ram_reg_1010__5_ ( .D(n12542), .CP(wclk), .Q(ram[8301]) );
  DFF ram_reg_1010__4_ ( .D(n12541), .CP(wclk), .Q(ram[8300]) );
  DFF ram_reg_1010__3_ ( .D(n12540), .CP(wclk), .Q(ram[8299]) );
  DFF ram_reg_1010__2_ ( .D(n12539), .CP(wclk), .Q(ram[8298]) );
  DFF ram_reg_1010__1_ ( .D(n12538), .CP(wclk), .Q(ram[8297]) );
  DFF ram_reg_1010__0_ ( .D(n12537), .CP(wclk), .Q(ram[8296]) );
  DFF ram_reg_1018__7_ ( .D(n12480), .CP(wclk), .Q(ram[8239]) );
  DFF ram_reg_1018__6_ ( .D(n12479), .CP(wclk), .Q(ram[8238]) );
  DFF ram_reg_1018__5_ ( .D(n12478), .CP(wclk), .Q(ram[8237]) );
  DFF ram_reg_1018__4_ ( .D(n12477), .CP(wclk), .Q(ram[8236]) );
  DFF ram_reg_1018__3_ ( .D(n12476), .CP(wclk), .Q(ram[8235]) );
  DFF ram_reg_1018__2_ ( .D(n12475), .CP(wclk), .Q(ram[8234]) );
  DFF ram_reg_1018__1_ ( .D(n12474), .CP(wclk), .Q(ram[8233]) );
  DFF ram_reg_1018__0_ ( .D(n12473), .CP(wclk), .Q(ram[8232]) );
  DFF ram_reg_1022__7_ ( .D(n12448), .CP(wclk), .Q(ram[8207]) );
  DFF ram_reg_1022__6_ ( .D(n12447), .CP(wclk), .Q(ram[8206]) );
  DFF ram_reg_1022__5_ ( .D(n12446), .CP(wclk), .Q(ram[8205]) );
  DFF ram_reg_1022__4_ ( .D(n12445), .CP(wclk), .Q(ram[8204]) );
  DFF ram_reg_1022__3_ ( .D(n12444), .CP(wclk), .Q(ram[8203]) );
  DFF ram_reg_1022__2_ ( .D(n12443), .CP(wclk), .Q(ram[8202]) );
  DFF ram_reg_1022__1_ ( .D(n12442), .CP(wclk), .Q(ram[8201]) );
  DFF ram_reg_1022__0_ ( .D(n12441), .CP(wclk), .Q(ram[8200]) );
  DFF ram_reg_1066__7_ ( .D(n12096), .CP(wclk), .Q(ram[7855]) );
  DFF ram_reg_1066__6_ ( .D(n12095), .CP(wclk), .Q(ram[7854]) );
  DFF ram_reg_1066__5_ ( .D(n12094), .CP(wclk), .Q(ram[7853]) );
  DFF ram_reg_1066__4_ ( .D(n12093), .CP(wclk), .Q(ram[7852]) );
  DFF ram_reg_1066__3_ ( .D(n12092), .CP(wclk), .Q(ram[7851]) );
  DFF ram_reg_1066__2_ ( .D(n12091), .CP(wclk), .Q(ram[7850]) );
  DFF ram_reg_1066__1_ ( .D(n12090), .CP(wclk), .Q(ram[7849]) );
  DFF ram_reg_1066__0_ ( .D(n12089), .CP(wclk), .Q(ram[7848]) );
  DFF ram_reg_1082__7_ ( .D(n11968), .CP(wclk), .Q(ram[7727]) );
  DFF ram_reg_1082__6_ ( .D(n11967), .CP(wclk), .Q(ram[7726]) );
  DFF ram_reg_1082__5_ ( .D(n11966), .CP(wclk), .Q(ram[7725]) );
  DFF ram_reg_1082__4_ ( .D(n11965), .CP(wclk), .Q(ram[7724]) );
  DFF ram_reg_1082__3_ ( .D(n11964), .CP(wclk), .Q(ram[7723]) );
  DFF ram_reg_1082__2_ ( .D(n11963), .CP(wclk), .Q(ram[7722]) );
  DFF ram_reg_1082__1_ ( .D(n11962), .CP(wclk), .Q(ram[7721]) );
  DFF ram_reg_1082__0_ ( .D(n11961), .CP(wclk), .Q(ram[7720]) );
  DFF ram_reg_1162__7_ ( .D(n11328), .CP(wclk), .Q(ram[7087]) );
  DFF ram_reg_1162__6_ ( .D(n11327), .CP(wclk), .Q(ram[7086]) );
  DFF ram_reg_1162__5_ ( .D(n11326), .CP(wclk), .Q(ram[7085]) );
  DFF ram_reg_1162__4_ ( .D(n11325), .CP(wclk), .Q(ram[7084]) );
  DFF ram_reg_1162__3_ ( .D(n11324), .CP(wclk), .Q(ram[7083]) );
  DFF ram_reg_1162__2_ ( .D(n11323), .CP(wclk), .Q(ram[7082]) );
  DFF ram_reg_1162__1_ ( .D(n11322), .CP(wclk), .Q(ram[7081]) );
  DFF ram_reg_1162__0_ ( .D(n11321), .CP(wclk), .Q(ram[7080]) );
  DFF ram_reg_1166__7_ ( .D(n11296), .CP(wclk), .Q(ram[7055]) );
  DFF ram_reg_1166__6_ ( .D(n11295), .CP(wclk), .Q(ram[7054]) );
  DFF ram_reg_1166__5_ ( .D(n11294), .CP(wclk), .Q(ram[7053]) );
  DFF ram_reg_1166__4_ ( .D(n11293), .CP(wclk), .Q(ram[7052]) );
  DFF ram_reg_1166__3_ ( .D(n11292), .CP(wclk), .Q(ram[7051]) );
  DFF ram_reg_1166__2_ ( .D(n11291), .CP(wclk), .Q(ram[7050]) );
  DFF ram_reg_1166__1_ ( .D(n11290), .CP(wclk), .Q(ram[7049]) );
  DFF ram_reg_1166__0_ ( .D(n11289), .CP(wclk), .Q(ram[7048]) );
  DFF ram_reg_1178__7_ ( .D(n11200), .CP(wclk), .Q(ram[6959]) );
  DFF ram_reg_1178__6_ ( .D(n11199), .CP(wclk), .Q(ram[6958]) );
  DFF ram_reg_1178__5_ ( .D(n11198), .CP(wclk), .Q(ram[6957]) );
  DFF ram_reg_1178__4_ ( .D(n11197), .CP(wclk), .Q(ram[6956]) );
  DFF ram_reg_1178__3_ ( .D(n11196), .CP(wclk), .Q(ram[6955]) );
  DFF ram_reg_1178__2_ ( .D(n11195), .CP(wclk), .Q(ram[6954]) );
  DFF ram_reg_1178__1_ ( .D(n11194), .CP(wclk), .Q(ram[6953]) );
  DFF ram_reg_1178__0_ ( .D(n11193), .CP(wclk), .Q(ram[6952]) );
  DFF ram_reg_1182__7_ ( .D(n11168), .CP(wclk), .Q(ram[6927]) );
  DFF ram_reg_1182__6_ ( .D(n11167), .CP(wclk), .Q(ram[6926]) );
  DFF ram_reg_1182__5_ ( .D(n11166), .CP(wclk), .Q(ram[6925]) );
  DFF ram_reg_1182__4_ ( .D(n11165), .CP(wclk), .Q(ram[6924]) );
  DFF ram_reg_1182__3_ ( .D(n11164), .CP(wclk), .Q(ram[6923]) );
  DFF ram_reg_1182__2_ ( .D(n11163), .CP(wclk), .Q(ram[6922]) );
  DFF ram_reg_1182__1_ ( .D(n11162), .CP(wclk), .Q(ram[6921]) );
  DFF ram_reg_1182__0_ ( .D(n11161), .CP(wclk), .Q(ram[6920]) );
  DFF ram_reg_1186__7_ ( .D(n11136), .CP(wclk), .Q(ram[6895]) );
  DFF ram_reg_1186__6_ ( .D(n11135), .CP(wclk), .Q(ram[6894]) );
  DFF ram_reg_1186__5_ ( .D(n11134), .CP(wclk), .Q(ram[6893]) );
  DFF ram_reg_1186__4_ ( .D(n11133), .CP(wclk), .Q(ram[6892]) );
  DFF ram_reg_1186__3_ ( .D(n11132), .CP(wclk), .Q(ram[6891]) );
  DFF ram_reg_1186__2_ ( .D(n11131), .CP(wclk), .Q(ram[6890]) );
  DFF ram_reg_1186__1_ ( .D(n11130), .CP(wclk), .Q(ram[6889]) );
  DFF ram_reg_1186__0_ ( .D(n11129), .CP(wclk), .Q(ram[6888]) );
  DFF ram_reg_1194__7_ ( .D(n11072), .CP(wclk), .Q(ram[6831]) );
  DFF ram_reg_1194__6_ ( .D(n11071), .CP(wclk), .Q(ram[6830]) );
  DFF ram_reg_1194__5_ ( .D(n11070), .CP(wclk), .Q(ram[6829]) );
  DFF ram_reg_1194__4_ ( .D(n11069), .CP(wclk), .Q(ram[6828]) );
  DFF ram_reg_1194__3_ ( .D(n11068), .CP(wclk), .Q(ram[6827]) );
  DFF ram_reg_1194__2_ ( .D(n11067), .CP(wclk), .Q(ram[6826]) );
  DFF ram_reg_1194__1_ ( .D(n11066), .CP(wclk), .Q(ram[6825]) );
  DFF ram_reg_1194__0_ ( .D(n11065), .CP(wclk), .Q(ram[6824]) );
  DFF ram_reg_1198__7_ ( .D(n11040), .CP(wclk), .Q(ram[6799]) );
  DFF ram_reg_1198__6_ ( .D(n11039), .CP(wclk), .Q(ram[6798]) );
  DFF ram_reg_1198__5_ ( .D(n11038), .CP(wclk), .Q(ram[6797]) );
  DFF ram_reg_1198__4_ ( .D(n11037), .CP(wclk), .Q(ram[6796]) );
  DFF ram_reg_1198__3_ ( .D(n11036), .CP(wclk), .Q(ram[6795]) );
  DFF ram_reg_1198__2_ ( .D(n11035), .CP(wclk), .Q(ram[6794]) );
  DFF ram_reg_1198__1_ ( .D(n11034), .CP(wclk), .Q(ram[6793]) );
  DFF ram_reg_1198__0_ ( .D(n11033), .CP(wclk), .Q(ram[6792]) );
  DFF ram_reg_1202__7_ ( .D(n11008), .CP(wclk), .Q(ram[6767]) );
  DFF ram_reg_1202__6_ ( .D(n11007), .CP(wclk), .Q(ram[6766]) );
  DFF ram_reg_1202__5_ ( .D(n11006), .CP(wclk), .Q(ram[6765]) );
  DFF ram_reg_1202__4_ ( .D(n11005), .CP(wclk), .Q(ram[6764]) );
  DFF ram_reg_1202__3_ ( .D(n11004), .CP(wclk), .Q(ram[6763]) );
  DFF ram_reg_1202__2_ ( .D(n11003), .CP(wclk), .Q(ram[6762]) );
  DFF ram_reg_1202__1_ ( .D(n11002), .CP(wclk), .Q(ram[6761]) );
  DFF ram_reg_1202__0_ ( .D(n11001), .CP(wclk), .Q(ram[6760]) );
  DFF ram_reg_1210__7_ ( .D(n10944), .CP(wclk), .Q(ram[6703]) );
  DFF ram_reg_1210__6_ ( .D(n10943), .CP(wclk), .Q(ram[6702]) );
  DFF ram_reg_1210__5_ ( .D(n10942), .CP(wclk), .Q(ram[6701]) );
  DFF ram_reg_1210__4_ ( .D(n10941), .CP(wclk), .Q(ram[6700]) );
  DFF ram_reg_1210__3_ ( .D(n10940), .CP(wclk), .Q(ram[6699]) );
  DFF ram_reg_1210__2_ ( .D(n10939), .CP(wclk), .Q(ram[6698]) );
  DFF ram_reg_1210__1_ ( .D(n10938), .CP(wclk), .Q(ram[6697]) );
  DFF ram_reg_1210__0_ ( .D(n10937), .CP(wclk), .Q(ram[6696]) );
  DFF ram_reg_1214__7_ ( .D(n10912), .CP(wclk), .Q(ram[6671]) );
  DFF ram_reg_1214__6_ ( .D(n10911), .CP(wclk), .Q(ram[6670]) );
  DFF ram_reg_1214__5_ ( .D(n10910), .CP(wclk), .Q(ram[6669]) );
  DFF ram_reg_1214__4_ ( .D(n10909), .CP(wclk), .Q(ram[6668]) );
  DFF ram_reg_1214__3_ ( .D(n10908), .CP(wclk), .Q(ram[6667]) );
  DFF ram_reg_1214__2_ ( .D(n10907), .CP(wclk), .Q(ram[6666]) );
  DFF ram_reg_1214__1_ ( .D(n10906), .CP(wclk), .Q(ram[6665]) );
  DFF ram_reg_1214__0_ ( .D(n10905), .CP(wclk), .Q(ram[6664]) );
  DFF ram_reg_1226__7_ ( .D(n10816), .CP(wclk), .Q(ram[6575]) );
  DFF ram_reg_1226__6_ ( .D(n10815), .CP(wclk), .Q(ram[6574]) );
  DFF ram_reg_1226__5_ ( .D(n10814), .CP(wclk), .Q(ram[6573]) );
  DFF ram_reg_1226__4_ ( .D(n10813), .CP(wclk), .Q(ram[6572]) );
  DFF ram_reg_1226__3_ ( .D(n10812), .CP(wclk), .Q(ram[6571]) );
  DFF ram_reg_1226__2_ ( .D(n10811), .CP(wclk), .Q(ram[6570]) );
  DFF ram_reg_1226__1_ ( .D(n10810), .CP(wclk), .Q(ram[6569]) );
  DFF ram_reg_1226__0_ ( .D(n10809), .CP(wclk), .Q(ram[6568]) );
  DFF ram_reg_1242__7_ ( .D(n10688), .CP(wclk), .Q(ram[6447]) );
  DFF ram_reg_1242__6_ ( .D(n10687), .CP(wclk), .Q(ram[6446]) );
  DFF ram_reg_1242__5_ ( .D(n10686), .CP(wclk), .Q(ram[6445]) );
  DFF ram_reg_1242__4_ ( .D(n10685), .CP(wclk), .Q(ram[6444]) );
  DFF ram_reg_1242__3_ ( .D(n10684), .CP(wclk), .Q(ram[6443]) );
  DFF ram_reg_1242__2_ ( .D(n10683), .CP(wclk), .Q(ram[6442]) );
  DFF ram_reg_1242__1_ ( .D(n10682), .CP(wclk), .Q(ram[6441]) );
  DFF ram_reg_1242__0_ ( .D(n10681), .CP(wclk), .Q(ram[6440]) );
  DFF ram_reg_1258__7_ ( .D(n10560), .CP(wclk), .Q(ram[6319]) );
  DFF ram_reg_1258__6_ ( .D(n10559), .CP(wclk), .Q(ram[6318]) );
  DFF ram_reg_1258__5_ ( .D(n10558), .CP(wclk), .Q(ram[6317]) );
  DFF ram_reg_1258__4_ ( .D(n10557), .CP(wclk), .Q(ram[6316]) );
  DFF ram_reg_1258__3_ ( .D(n10556), .CP(wclk), .Q(ram[6315]) );
  DFF ram_reg_1258__2_ ( .D(n10555), .CP(wclk), .Q(ram[6314]) );
  DFF ram_reg_1258__1_ ( .D(n10554), .CP(wclk), .Q(ram[6313]) );
  DFF ram_reg_1258__0_ ( .D(n10553), .CP(wclk), .Q(ram[6312]) );
  DFF ram_reg_1262__7_ ( .D(n10528), .CP(wclk), .Q(ram[6287]) );
  DFF ram_reg_1262__6_ ( .D(n10527), .CP(wclk), .Q(ram[6286]) );
  DFF ram_reg_1262__5_ ( .D(n10526), .CP(wclk), .Q(ram[6285]) );
  DFF ram_reg_1262__4_ ( .D(n10525), .CP(wclk), .Q(ram[6284]) );
  DFF ram_reg_1262__3_ ( .D(n10524), .CP(wclk), .Q(ram[6283]) );
  DFF ram_reg_1262__2_ ( .D(n10523), .CP(wclk), .Q(ram[6282]) );
  DFF ram_reg_1262__1_ ( .D(n10522), .CP(wclk), .Q(ram[6281]) );
  DFF ram_reg_1262__0_ ( .D(n10521), .CP(wclk), .Q(ram[6280]) );
  DFF ram_reg_1274__7_ ( .D(n10432), .CP(wclk), .Q(ram[6191]) );
  DFF ram_reg_1274__6_ ( .D(n10431), .CP(wclk), .Q(ram[6190]) );
  DFF ram_reg_1274__5_ ( .D(n10430), .CP(wclk), .Q(ram[6189]) );
  DFF ram_reg_1274__4_ ( .D(n10429), .CP(wclk), .Q(ram[6188]) );
  DFF ram_reg_1274__3_ ( .D(n10428), .CP(wclk), .Q(ram[6187]) );
  DFF ram_reg_1274__2_ ( .D(n10427), .CP(wclk), .Q(ram[6186]) );
  DFF ram_reg_1274__1_ ( .D(n10426), .CP(wclk), .Q(ram[6185]) );
  DFF ram_reg_1274__0_ ( .D(n10425), .CP(wclk), .Q(ram[6184]) );
  DFF ram_reg_1278__7_ ( .D(n10400), .CP(wclk), .Q(ram[6159]) );
  DFF ram_reg_1278__6_ ( .D(n10399), .CP(wclk), .Q(ram[6158]) );
  DFF ram_reg_1278__5_ ( .D(n10398), .CP(wclk), .Q(ram[6157]) );
  DFF ram_reg_1278__4_ ( .D(n10397), .CP(wclk), .Q(ram[6156]) );
  DFF ram_reg_1278__3_ ( .D(n10396), .CP(wclk), .Q(ram[6155]) );
  DFF ram_reg_1278__2_ ( .D(n10395), .CP(wclk), .Q(ram[6154]) );
  DFF ram_reg_1278__1_ ( .D(n10394), .CP(wclk), .Q(ram[6153]) );
  DFF ram_reg_1278__0_ ( .D(n10393), .CP(wclk), .Q(ram[6152]) );
  DFF ram_reg_1290__7_ ( .D(n10304), .CP(wclk), .Q(ram[6063]) );
  DFF ram_reg_1290__6_ ( .D(n10303), .CP(wclk), .Q(ram[6062]) );
  DFF ram_reg_1290__5_ ( .D(n10302), .CP(wclk), .Q(ram[6061]) );
  DFF ram_reg_1290__4_ ( .D(n10301), .CP(wclk), .Q(ram[6060]) );
  DFF ram_reg_1290__3_ ( .D(n10300), .CP(wclk), .Q(ram[6059]) );
  DFF ram_reg_1290__2_ ( .D(n10299), .CP(wclk), .Q(ram[6058]) );
  DFF ram_reg_1290__1_ ( .D(n10298), .CP(wclk), .Q(ram[6057]) );
  DFF ram_reg_1290__0_ ( .D(n10297), .CP(wclk), .Q(ram[6056]) );
  DFF ram_reg_1294__7_ ( .D(n10272), .CP(wclk), .Q(ram[6031]) );
  DFF ram_reg_1294__6_ ( .D(n10271), .CP(wclk), .Q(ram[6030]) );
  DFF ram_reg_1294__5_ ( .D(n10270), .CP(wclk), .Q(ram[6029]) );
  DFF ram_reg_1294__4_ ( .D(n10269), .CP(wclk), .Q(ram[6028]) );
  DFF ram_reg_1294__3_ ( .D(n10268), .CP(wclk), .Q(ram[6027]) );
  DFF ram_reg_1294__2_ ( .D(n10267), .CP(wclk), .Q(ram[6026]) );
  DFF ram_reg_1294__1_ ( .D(n10266), .CP(wclk), .Q(ram[6025]) );
  DFF ram_reg_1294__0_ ( .D(n10265), .CP(wclk), .Q(ram[6024]) );
  DFF ram_reg_1306__7_ ( .D(n10176), .CP(wclk), .Q(ram[5935]) );
  DFF ram_reg_1306__6_ ( .D(n10175), .CP(wclk), .Q(ram[5934]) );
  DFF ram_reg_1306__5_ ( .D(n10174), .CP(wclk), .Q(ram[5933]) );
  DFF ram_reg_1306__4_ ( .D(n10173), .CP(wclk), .Q(ram[5932]) );
  DFF ram_reg_1306__3_ ( .D(n10172), .CP(wclk), .Q(ram[5931]) );
  DFF ram_reg_1306__2_ ( .D(n10171), .CP(wclk), .Q(ram[5930]) );
  DFF ram_reg_1306__1_ ( .D(n10170), .CP(wclk), .Q(ram[5929]) );
  DFF ram_reg_1306__0_ ( .D(n10169), .CP(wclk), .Q(ram[5928]) );
  DFF ram_reg_1322__7_ ( .D(n10048), .CP(wclk), .Q(ram[5807]) );
  DFF ram_reg_1322__6_ ( .D(n10047), .CP(wclk), .Q(ram[5806]) );
  DFF ram_reg_1322__5_ ( .D(n10046), .CP(wclk), .Q(ram[5805]) );
  DFF ram_reg_1322__4_ ( .D(n10045), .CP(wclk), .Q(ram[5804]) );
  DFF ram_reg_1322__3_ ( .D(n10044), .CP(wclk), .Q(ram[5803]) );
  DFF ram_reg_1322__2_ ( .D(n10043), .CP(wclk), .Q(ram[5802]) );
  DFF ram_reg_1322__1_ ( .D(n10042), .CP(wclk), .Q(ram[5801]) );
  DFF ram_reg_1322__0_ ( .D(n10041), .CP(wclk), .Q(ram[5800]) );
  DFF ram_reg_1326__7_ ( .D(n10016), .CP(wclk), .Q(ram[5775]) );
  DFF ram_reg_1326__6_ ( .D(n10015), .CP(wclk), .Q(ram[5774]) );
  DFF ram_reg_1326__5_ ( .D(n10014), .CP(wclk), .Q(ram[5773]) );
  DFF ram_reg_1326__4_ ( .D(n10013), .CP(wclk), .Q(ram[5772]) );
  DFF ram_reg_1326__3_ ( .D(n10012), .CP(wclk), .Q(ram[5771]) );
  DFF ram_reg_1326__2_ ( .D(n10011), .CP(wclk), .Q(ram[5770]) );
  DFF ram_reg_1326__1_ ( .D(n10010), .CP(wclk), .Q(ram[5769]) );
  DFF ram_reg_1326__0_ ( .D(n10009), .CP(wclk), .Q(ram[5768]) );
  DFF ram_reg_1338__7_ ( .D(n9920), .CP(wclk), .Q(ram[5679]) );
  DFF ram_reg_1338__6_ ( .D(n9919), .CP(wclk), .Q(ram[5678]) );
  DFF ram_reg_1338__5_ ( .D(n9918), .CP(wclk), .Q(ram[5677]) );
  DFF ram_reg_1338__4_ ( .D(n9917), .CP(wclk), .Q(ram[5676]) );
  DFF ram_reg_1338__3_ ( .D(n9916), .CP(wclk), .Q(ram[5675]) );
  DFF ram_reg_1338__2_ ( .D(n9915), .CP(wclk), .Q(ram[5674]) );
  DFF ram_reg_1338__1_ ( .D(n9914), .CP(wclk), .Q(ram[5673]) );
  DFF ram_reg_1338__0_ ( .D(n9913), .CP(wclk), .Q(ram[5672]) );
  DFF ram_reg_1342__7_ ( .D(n9888), .CP(wclk), .Q(ram[5647]) );
  DFF ram_reg_1342__6_ ( .D(n9887), .CP(wclk), .Q(ram[5646]) );
  DFF ram_reg_1342__5_ ( .D(n9886), .CP(wclk), .Q(ram[5645]) );
  DFF ram_reg_1342__4_ ( .D(n9885), .CP(wclk), .Q(ram[5644]) );
  DFF ram_reg_1342__3_ ( .D(n9884), .CP(wclk), .Q(ram[5643]) );
  DFF ram_reg_1342__2_ ( .D(n9883), .CP(wclk), .Q(ram[5642]) );
  DFF ram_reg_1342__1_ ( .D(n9882), .CP(wclk), .Q(ram[5641]) );
  DFF ram_reg_1342__0_ ( .D(n9881), .CP(wclk), .Q(ram[5640]) );
  DFF ram_reg_1386__7_ ( .D(n9536), .CP(wclk), .Q(ram[5295]) );
  DFF ram_reg_1386__6_ ( .D(n9535), .CP(wclk), .Q(ram[5294]) );
  DFF ram_reg_1386__5_ ( .D(n9534), .CP(wclk), .Q(ram[5293]) );
  DFF ram_reg_1386__4_ ( .D(n9533), .CP(wclk), .Q(ram[5292]) );
  DFF ram_reg_1386__3_ ( .D(n9532), .CP(wclk), .Q(ram[5291]) );
  DFF ram_reg_1386__2_ ( .D(n9531), .CP(wclk), .Q(ram[5290]) );
  DFF ram_reg_1386__1_ ( .D(n9530), .CP(wclk), .Q(ram[5289]) );
  DFF ram_reg_1386__0_ ( .D(n9529), .CP(wclk), .Q(ram[5288]) );
  DFF ram_reg_1402__7_ ( .D(n9408), .CP(wclk), .Q(ram[5167]) );
  DFF ram_reg_1402__6_ ( .D(n9407), .CP(wclk), .Q(ram[5166]) );
  DFF ram_reg_1402__5_ ( .D(n9406), .CP(wclk), .Q(ram[5165]) );
  DFF ram_reg_1402__4_ ( .D(n9405), .CP(wclk), .Q(ram[5164]) );
  DFF ram_reg_1402__3_ ( .D(n9404), .CP(wclk), .Q(ram[5163]) );
  DFF ram_reg_1402__2_ ( .D(n9403), .CP(wclk), .Q(ram[5162]) );
  DFF ram_reg_1402__1_ ( .D(n9402), .CP(wclk), .Q(ram[5161]) );
  DFF ram_reg_1402__0_ ( .D(n9401), .CP(wclk), .Q(ram[5160]) );
  DFF ram_reg_1410__7_ ( .D(n9344), .CP(wclk), .Q(ram[5103]) );
  DFF ram_reg_1410__6_ ( .D(n9343), .CP(wclk), .Q(ram[5102]) );
  DFF ram_reg_1410__5_ ( .D(n9342), .CP(wclk), .Q(ram[5101]) );
  DFF ram_reg_1410__4_ ( .D(n9341), .CP(wclk), .Q(ram[5100]) );
  DFF ram_reg_1410__3_ ( .D(n9340), .CP(wclk), .Q(ram[5099]) );
  DFF ram_reg_1410__2_ ( .D(n9339), .CP(wclk), .Q(ram[5098]) );
  DFF ram_reg_1410__1_ ( .D(n9338), .CP(wclk), .Q(ram[5097]) );
  DFF ram_reg_1410__0_ ( .D(n9337), .CP(wclk), .Q(ram[5096]) );
  DFF ram_reg_1418__7_ ( .D(n9280), .CP(wclk), .Q(ram[5039]) );
  DFF ram_reg_1418__6_ ( .D(n9279), .CP(wclk), .Q(ram[5038]) );
  DFF ram_reg_1418__5_ ( .D(n9278), .CP(wclk), .Q(ram[5037]) );
  DFF ram_reg_1418__4_ ( .D(n9277), .CP(wclk), .Q(ram[5036]) );
  DFF ram_reg_1418__3_ ( .D(n9276), .CP(wclk), .Q(ram[5035]) );
  DFF ram_reg_1418__2_ ( .D(n9275), .CP(wclk), .Q(ram[5034]) );
  DFF ram_reg_1418__1_ ( .D(n9274), .CP(wclk), .Q(ram[5033]) );
  DFF ram_reg_1418__0_ ( .D(n9273), .CP(wclk), .Q(ram[5032]) );
  DFF ram_reg_1422__7_ ( .D(n9248), .CP(wclk), .Q(ram[5007]) );
  DFF ram_reg_1422__6_ ( .D(n9247), .CP(wclk), .Q(ram[5006]) );
  DFF ram_reg_1422__5_ ( .D(n9246), .CP(wclk), .Q(ram[5005]) );
  DFF ram_reg_1422__4_ ( .D(n9245), .CP(wclk), .Q(ram[5004]) );
  DFF ram_reg_1422__3_ ( .D(n9244), .CP(wclk), .Q(ram[5003]) );
  DFF ram_reg_1422__2_ ( .D(n9243), .CP(wclk), .Q(ram[5002]) );
  DFF ram_reg_1422__1_ ( .D(n9242), .CP(wclk), .Q(ram[5001]) );
  DFF ram_reg_1422__0_ ( .D(n9241), .CP(wclk), .Q(ram[5000]) );
  DFF ram_reg_1426__7_ ( .D(n9216), .CP(wclk), .Q(ram[4975]) );
  DFF ram_reg_1426__6_ ( .D(n9215), .CP(wclk), .Q(ram[4974]) );
  DFF ram_reg_1426__5_ ( .D(n9214), .CP(wclk), .Q(ram[4973]) );
  DFF ram_reg_1426__4_ ( .D(n9213), .CP(wclk), .Q(ram[4972]) );
  DFF ram_reg_1426__3_ ( .D(n9212), .CP(wclk), .Q(ram[4971]) );
  DFF ram_reg_1426__2_ ( .D(n9211), .CP(wclk), .Q(ram[4970]) );
  DFF ram_reg_1426__1_ ( .D(n9210), .CP(wclk), .Q(ram[4969]) );
  DFF ram_reg_1426__0_ ( .D(n9209), .CP(wclk), .Q(ram[4968]) );
  DFF ram_reg_1434__7_ ( .D(n9152), .CP(wclk), .Q(ram[4911]) );
  DFF ram_reg_1434__6_ ( .D(n9151), .CP(wclk), .Q(ram[4910]) );
  DFF ram_reg_1434__5_ ( .D(n9150), .CP(wclk), .Q(ram[4909]) );
  DFF ram_reg_1434__4_ ( .D(n9149), .CP(wclk), .Q(ram[4908]) );
  DFF ram_reg_1434__3_ ( .D(n9148), .CP(wclk), .Q(ram[4907]) );
  DFF ram_reg_1434__2_ ( .D(n9147), .CP(wclk), .Q(ram[4906]) );
  DFF ram_reg_1434__1_ ( .D(n9146), .CP(wclk), .Q(ram[4905]) );
  DFF ram_reg_1434__0_ ( .D(n9145), .CP(wclk), .Q(ram[4904]) );
  DFF ram_reg_1438__7_ ( .D(n9120), .CP(wclk), .Q(ram[4879]) );
  DFF ram_reg_1438__6_ ( .D(n9119), .CP(wclk), .Q(ram[4878]) );
  DFF ram_reg_1438__5_ ( .D(n9118), .CP(wclk), .Q(ram[4877]) );
  DFF ram_reg_1438__4_ ( .D(n9117), .CP(wclk), .Q(ram[4876]) );
  DFF ram_reg_1438__3_ ( .D(n9116), .CP(wclk), .Q(ram[4875]) );
  DFF ram_reg_1438__2_ ( .D(n9115), .CP(wclk), .Q(ram[4874]) );
  DFF ram_reg_1438__1_ ( .D(n9114), .CP(wclk), .Q(ram[4873]) );
  DFF ram_reg_1438__0_ ( .D(n9113), .CP(wclk), .Q(ram[4872]) );
  DFF ram_reg_1442__7_ ( .D(n9088), .CP(wclk), .Q(ram[4847]) );
  DFF ram_reg_1442__6_ ( .D(n9087), .CP(wclk), .Q(ram[4846]) );
  DFF ram_reg_1442__5_ ( .D(n9086), .CP(wclk), .Q(ram[4845]) );
  DFF ram_reg_1442__4_ ( .D(n9085), .CP(wclk), .Q(ram[4844]) );
  DFF ram_reg_1442__3_ ( .D(n9084), .CP(wclk), .Q(ram[4843]) );
  DFF ram_reg_1442__2_ ( .D(n9083), .CP(wclk), .Q(ram[4842]) );
  DFF ram_reg_1442__1_ ( .D(n9082), .CP(wclk), .Q(ram[4841]) );
  DFF ram_reg_1442__0_ ( .D(n9081), .CP(wclk), .Q(ram[4840]) );
  DFF ram_reg_1446__7_ ( .D(n9056), .CP(wclk), .Q(ram[4815]) );
  DFF ram_reg_1446__6_ ( .D(n9055), .CP(wclk), .Q(ram[4814]) );
  DFF ram_reg_1446__5_ ( .D(n9054), .CP(wclk), .Q(ram[4813]) );
  DFF ram_reg_1446__4_ ( .D(n9053), .CP(wclk), .Q(ram[4812]) );
  DFF ram_reg_1446__3_ ( .D(n9052), .CP(wclk), .Q(ram[4811]) );
  DFF ram_reg_1446__2_ ( .D(n9051), .CP(wclk), .Q(ram[4810]) );
  DFF ram_reg_1446__1_ ( .D(n9050), .CP(wclk), .Q(ram[4809]) );
  DFF ram_reg_1446__0_ ( .D(n9049), .CP(wclk), .Q(ram[4808]) );
  DFF ram_reg_1450__7_ ( .D(n9024), .CP(wclk), .Q(ram[4783]) );
  DFF ram_reg_1450__6_ ( .D(n9023), .CP(wclk), .Q(ram[4782]) );
  DFF ram_reg_1450__5_ ( .D(n9022), .CP(wclk), .Q(ram[4781]) );
  DFF ram_reg_1450__4_ ( .D(n9021), .CP(wclk), .Q(ram[4780]) );
  DFF ram_reg_1450__3_ ( .D(n9020), .CP(wclk), .Q(ram[4779]) );
  DFF ram_reg_1450__2_ ( .D(n9019), .CP(wclk), .Q(ram[4778]) );
  DFF ram_reg_1450__1_ ( .D(n9018), .CP(wclk), .Q(ram[4777]) );
  DFF ram_reg_1450__0_ ( .D(n9017), .CP(wclk), .Q(ram[4776]) );
  DFF ram_reg_1454__7_ ( .D(n8992), .CP(wclk), .Q(ram[4751]) );
  DFF ram_reg_1454__6_ ( .D(n8991), .CP(wclk), .Q(ram[4750]) );
  DFF ram_reg_1454__5_ ( .D(n8990), .CP(wclk), .Q(ram[4749]) );
  DFF ram_reg_1454__4_ ( .D(n8989), .CP(wclk), .Q(ram[4748]) );
  DFF ram_reg_1454__3_ ( .D(n8988), .CP(wclk), .Q(ram[4747]) );
  DFF ram_reg_1454__2_ ( .D(n8987), .CP(wclk), .Q(ram[4746]) );
  DFF ram_reg_1454__1_ ( .D(n8986), .CP(wclk), .Q(ram[4745]) );
  DFF ram_reg_1454__0_ ( .D(n8985), .CP(wclk), .Q(ram[4744]) );
  DFF ram_reg_1458__7_ ( .D(n8960), .CP(wclk), .Q(ram[4719]) );
  DFF ram_reg_1458__6_ ( .D(n8959), .CP(wclk), .Q(ram[4718]) );
  DFF ram_reg_1458__5_ ( .D(n8958), .CP(wclk), .Q(ram[4717]) );
  DFF ram_reg_1458__4_ ( .D(n8957), .CP(wclk), .Q(ram[4716]) );
  DFF ram_reg_1458__3_ ( .D(n8956), .CP(wclk), .Q(ram[4715]) );
  DFF ram_reg_1458__2_ ( .D(n8955), .CP(wclk), .Q(ram[4714]) );
  DFF ram_reg_1458__1_ ( .D(n8954), .CP(wclk), .Q(ram[4713]) );
  DFF ram_reg_1458__0_ ( .D(n8953), .CP(wclk), .Q(ram[4712]) );
  DFF ram_reg_1462__7_ ( .D(n8928), .CP(wclk), .Q(ram[4687]) );
  DFF ram_reg_1462__6_ ( .D(n8927), .CP(wclk), .Q(ram[4686]) );
  DFF ram_reg_1462__5_ ( .D(n8926), .CP(wclk), .Q(ram[4685]) );
  DFF ram_reg_1462__4_ ( .D(n8925), .CP(wclk), .Q(ram[4684]) );
  DFF ram_reg_1462__3_ ( .D(n8924), .CP(wclk), .Q(ram[4683]) );
  DFF ram_reg_1462__2_ ( .D(n8923), .CP(wclk), .Q(ram[4682]) );
  DFF ram_reg_1462__1_ ( .D(n8922), .CP(wclk), .Q(ram[4681]) );
  DFF ram_reg_1462__0_ ( .D(n8921), .CP(wclk), .Q(ram[4680]) );
  DFF ram_reg_1466__7_ ( .D(n8896), .CP(wclk), .Q(ram[4655]) );
  DFF ram_reg_1466__6_ ( .D(n8895), .CP(wclk), .Q(ram[4654]) );
  DFF ram_reg_1466__5_ ( .D(n8894), .CP(wclk), .Q(ram[4653]) );
  DFF ram_reg_1466__4_ ( .D(n8893), .CP(wclk), .Q(ram[4652]) );
  DFF ram_reg_1466__3_ ( .D(n8892), .CP(wclk), .Q(ram[4651]) );
  DFF ram_reg_1466__2_ ( .D(n8891), .CP(wclk), .Q(ram[4650]) );
  DFF ram_reg_1466__1_ ( .D(n8890), .CP(wclk), .Q(ram[4649]) );
  DFF ram_reg_1466__0_ ( .D(n8889), .CP(wclk), .Q(ram[4648]) );
  DFF ram_reg_1470__7_ ( .D(n8864), .CP(wclk), .Q(ram[4623]) );
  DFF ram_reg_1470__6_ ( .D(n8863), .CP(wclk), .Q(ram[4622]) );
  DFF ram_reg_1470__5_ ( .D(n8862), .CP(wclk), .Q(ram[4621]) );
  DFF ram_reg_1470__4_ ( .D(n8861), .CP(wclk), .Q(ram[4620]) );
  DFF ram_reg_1470__3_ ( .D(n8860), .CP(wclk), .Q(ram[4619]) );
  DFF ram_reg_1470__2_ ( .D(n8859), .CP(wclk), .Q(ram[4618]) );
  DFF ram_reg_1470__1_ ( .D(n8858), .CP(wclk), .Q(ram[4617]) );
  DFF ram_reg_1470__0_ ( .D(n8857), .CP(wclk), .Q(ram[4616]) );
  DFF ram_reg_1474__7_ ( .D(n8832), .CP(wclk), .Q(ram[4591]) );
  DFF ram_reg_1474__6_ ( .D(n8831), .CP(wclk), .Q(ram[4590]) );
  DFF ram_reg_1474__5_ ( .D(n8830), .CP(wclk), .Q(ram[4589]) );
  DFF ram_reg_1474__4_ ( .D(n8829), .CP(wclk), .Q(ram[4588]) );
  DFF ram_reg_1474__3_ ( .D(n8828), .CP(wclk), .Q(ram[4587]) );
  DFF ram_reg_1474__2_ ( .D(n8827), .CP(wclk), .Q(ram[4586]) );
  DFF ram_reg_1474__1_ ( .D(n8826), .CP(wclk), .Q(ram[4585]) );
  DFF ram_reg_1474__0_ ( .D(n8825), .CP(wclk), .Q(ram[4584]) );
  DFF ram_reg_1482__7_ ( .D(n8768), .CP(wclk), .Q(ram[4527]) );
  DFF ram_reg_1482__6_ ( .D(n8767), .CP(wclk), .Q(ram[4526]) );
  DFF ram_reg_1482__5_ ( .D(n8766), .CP(wclk), .Q(ram[4525]) );
  DFF ram_reg_1482__4_ ( .D(n8765), .CP(wclk), .Q(ram[4524]) );
  DFF ram_reg_1482__3_ ( .D(n8764), .CP(wclk), .Q(ram[4523]) );
  DFF ram_reg_1482__2_ ( .D(n8763), .CP(wclk), .Q(ram[4522]) );
  DFF ram_reg_1482__1_ ( .D(n8762), .CP(wclk), .Q(ram[4521]) );
  DFF ram_reg_1482__0_ ( .D(n8761), .CP(wclk), .Q(ram[4520]) );
  DFF ram_reg_1486__7_ ( .D(n8736), .CP(wclk), .Q(ram[4495]) );
  DFF ram_reg_1486__6_ ( .D(n8735), .CP(wclk), .Q(ram[4494]) );
  DFF ram_reg_1486__5_ ( .D(n8734), .CP(wclk), .Q(ram[4493]) );
  DFF ram_reg_1486__4_ ( .D(n8733), .CP(wclk), .Q(ram[4492]) );
  DFF ram_reg_1486__3_ ( .D(n8732), .CP(wclk), .Q(ram[4491]) );
  DFF ram_reg_1486__2_ ( .D(n8731), .CP(wclk), .Q(ram[4490]) );
  DFF ram_reg_1486__1_ ( .D(n8730), .CP(wclk), .Q(ram[4489]) );
  DFF ram_reg_1486__0_ ( .D(n8729), .CP(wclk), .Q(ram[4488]) );
  DFF ram_reg_1498__7_ ( .D(n8640), .CP(wclk), .Q(ram[4399]) );
  DFF ram_reg_1498__6_ ( .D(n8639), .CP(wclk), .Q(ram[4398]) );
  DFF ram_reg_1498__5_ ( .D(n8638), .CP(wclk), .Q(ram[4397]) );
  DFF ram_reg_1498__4_ ( .D(n8637), .CP(wclk), .Q(ram[4396]) );
  DFF ram_reg_1498__3_ ( .D(n8636), .CP(wclk), .Q(ram[4395]) );
  DFF ram_reg_1498__2_ ( .D(n8635), .CP(wclk), .Q(ram[4394]) );
  DFF ram_reg_1498__1_ ( .D(n8634), .CP(wclk), .Q(ram[4393]) );
  DFF ram_reg_1498__0_ ( .D(n8633), .CP(wclk), .Q(ram[4392]) );
  DFF ram_reg_1502__7_ ( .D(n8608), .CP(wclk), .Q(ram[4367]) );
  DFF ram_reg_1502__6_ ( .D(n8607), .CP(wclk), .Q(ram[4366]) );
  DFF ram_reg_1502__5_ ( .D(n8606), .CP(wclk), .Q(ram[4365]) );
  DFF ram_reg_1502__4_ ( .D(n8605), .CP(wclk), .Q(ram[4364]) );
  DFF ram_reg_1502__3_ ( .D(n8604), .CP(wclk), .Q(ram[4363]) );
  DFF ram_reg_1502__2_ ( .D(n8603), .CP(wclk), .Q(ram[4362]) );
  DFF ram_reg_1502__1_ ( .D(n8602), .CP(wclk), .Q(ram[4361]) );
  DFF ram_reg_1502__0_ ( .D(n8601), .CP(wclk), .Q(ram[4360]) );
  DFF ram_reg_1506__7_ ( .D(n8576), .CP(wclk), .Q(ram[4335]) );
  DFF ram_reg_1506__6_ ( .D(n8575), .CP(wclk), .Q(ram[4334]) );
  DFF ram_reg_1506__5_ ( .D(n8574), .CP(wclk), .Q(ram[4333]) );
  DFF ram_reg_1506__4_ ( .D(n8573), .CP(wclk), .Q(ram[4332]) );
  DFF ram_reg_1506__3_ ( .D(n8572), .CP(wclk), .Q(ram[4331]) );
  DFF ram_reg_1506__2_ ( .D(n8571), .CP(wclk), .Q(ram[4330]) );
  DFF ram_reg_1506__1_ ( .D(n8570), .CP(wclk), .Q(ram[4329]) );
  DFF ram_reg_1506__0_ ( .D(n8569), .CP(wclk), .Q(ram[4328]) );
  DFF ram_reg_1514__7_ ( .D(n8512), .CP(wclk), .Q(ram[4271]) );
  DFF ram_reg_1514__6_ ( .D(n8511), .CP(wclk), .Q(ram[4270]) );
  DFF ram_reg_1514__5_ ( .D(n8510), .CP(wclk), .Q(ram[4269]) );
  DFF ram_reg_1514__4_ ( .D(n8509), .CP(wclk), .Q(ram[4268]) );
  DFF ram_reg_1514__3_ ( .D(n8508), .CP(wclk), .Q(ram[4267]) );
  DFF ram_reg_1514__2_ ( .D(n8507), .CP(wclk), .Q(ram[4266]) );
  DFF ram_reg_1514__1_ ( .D(n8506), .CP(wclk), .Q(ram[4265]) );
  DFF ram_reg_1514__0_ ( .D(n8505), .CP(wclk), .Q(ram[4264]) );
  DFF ram_reg_1518__7_ ( .D(n8480), .CP(wclk), .Q(ram[4239]) );
  DFF ram_reg_1518__6_ ( .D(n8479), .CP(wclk), .Q(ram[4238]) );
  DFF ram_reg_1518__5_ ( .D(n8478), .CP(wclk), .Q(ram[4237]) );
  DFF ram_reg_1518__4_ ( .D(n8477), .CP(wclk), .Q(ram[4236]) );
  DFF ram_reg_1518__3_ ( .D(n8476), .CP(wclk), .Q(ram[4235]) );
  DFF ram_reg_1518__2_ ( .D(n8475), .CP(wclk), .Q(ram[4234]) );
  DFF ram_reg_1518__1_ ( .D(n8474), .CP(wclk), .Q(ram[4233]) );
  DFF ram_reg_1518__0_ ( .D(n8473), .CP(wclk), .Q(ram[4232]) );
  DFF ram_reg_1522__7_ ( .D(n8448), .CP(wclk), .Q(ram[4207]) );
  DFF ram_reg_1522__6_ ( .D(n8447), .CP(wclk), .Q(ram[4206]) );
  DFF ram_reg_1522__5_ ( .D(n8446), .CP(wclk), .Q(ram[4205]) );
  DFF ram_reg_1522__4_ ( .D(n8445), .CP(wclk), .Q(ram[4204]) );
  DFF ram_reg_1522__3_ ( .D(n8444), .CP(wclk), .Q(ram[4203]) );
  DFF ram_reg_1522__2_ ( .D(n8443), .CP(wclk), .Q(ram[4202]) );
  DFF ram_reg_1522__1_ ( .D(n8442), .CP(wclk), .Q(ram[4201]) );
  DFF ram_reg_1522__0_ ( .D(n8441), .CP(wclk), .Q(ram[4200]) );
  DFF ram_reg_1530__7_ ( .D(n8384), .CP(wclk), .Q(ram[4143]) );
  DFF ram_reg_1530__6_ ( .D(n8383), .CP(wclk), .Q(ram[4142]) );
  DFF ram_reg_1530__5_ ( .D(n8382), .CP(wclk), .Q(ram[4141]) );
  DFF ram_reg_1530__4_ ( .D(n8381), .CP(wclk), .Q(ram[4140]) );
  DFF ram_reg_1530__3_ ( .D(n8380), .CP(wclk), .Q(ram[4139]) );
  DFF ram_reg_1530__2_ ( .D(n8379), .CP(wclk), .Q(ram[4138]) );
  DFF ram_reg_1530__1_ ( .D(n8378), .CP(wclk), .Q(ram[4137]) );
  DFF ram_reg_1530__0_ ( .D(n8377), .CP(wclk), .Q(ram[4136]) );
  DFF ram_reg_1534__7_ ( .D(n8352), .CP(wclk), .Q(ram[4111]) );
  DFF ram_reg_1534__6_ ( .D(n8351), .CP(wclk), .Q(ram[4110]) );
  DFF ram_reg_1534__5_ ( .D(n8350), .CP(wclk), .Q(ram[4109]) );
  DFF ram_reg_1534__4_ ( .D(n8349), .CP(wclk), .Q(ram[4108]) );
  DFF ram_reg_1534__3_ ( .D(n8348), .CP(wclk), .Q(ram[4107]) );
  DFF ram_reg_1534__2_ ( .D(n8347), .CP(wclk), .Q(ram[4106]) );
  DFF ram_reg_1534__1_ ( .D(n8346), .CP(wclk), .Q(ram[4105]) );
  DFF ram_reg_1534__0_ ( .D(n8345), .CP(wclk), .Q(ram[4104]) );
  DFF ram_reg_1578__7_ ( .D(n8000), .CP(wclk), .Q(ram[3759]) );
  DFF ram_reg_1578__6_ ( .D(n7999), .CP(wclk), .Q(ram[3758]) );
  DFF ram_reg_1578__5_ ( .D(n7998), .CP(wclk), .Q(ram[3757]) );
  DFF ram_reg_1578__4_ ( .D(n7997), .CP(wclk), .Q(ram[3756]) );
  DFF ram_reg_1578__3_ ( .D(n7996), .CP(wclk), .Q(ram[3755]) );
  DFF ram_reg_1578__2_ ( .D(n7995), .CP(wclk), .Q(ram[3754]) );
  DFF ram_reg_1578__1_ ( .D(n7994), .CP(wclk), .Q(ram[3753]) );
  DFF ram_reg_1578__0_ ( .D(n7993), .CP(wclk), .Q(ram[3752]) );
  DFF ram_reg_1594__7_ ( .D(n7872), .CP(wclk), .Q(ram[3631]) );
  DFF ram_reg_1594__6_ ( .D(n7871), .CP(wclk), .Q(ram[3630]) );
  DFF ram_reg_1594__5_ ( .D(n7870), .CP(wclk), .Q(ram[3629]) );
  DFF ram_reg_1594__4_ ( .D(n7869), .CP(wclk), .Q(ram[3628]) );
  DFF ram_reg_1594__3_ ( .D(n7868), .CP(wclk), .Q(ram[3627]) );
  DFF ram_reg_1594__2_ ( .D(n7867), .CP(wclk), .Q(ram[3626]) );
  DFF ram_reg_1594__1_ ( .D(n7866), .CP(wclk), .Q(ram[3625]) );
  DFF ram_reg_1594__0_ ( .D(n7865), .CP(wclk), .Q(ram[3624]) );
  DFF ram_reg_1674__7_ ( .D(n7232), .CP(wclk), .Q(ram[2991]) );
  DFF ram_reg_1674__6_ ( .D(n7231), .CP(wclk), .Q(ram[2990]) );
  DFF ram_reg_1674__5_ ( .D(n7230), .CP(wclk), .Q(ram[2989]) );
  DFF ram_reg_1674__4_ ( .D(n7229), .CP(wclk), .Q(ram[2988]) );
  DFF ram_reg_1674__3_ ( .D(n7228), .CP(wclk), .Q(ram[2987]) );
  DFF ram_reg_1674__2_ ( .D(n7227), .CP(wclk), .Q(ram[2986]) );
  DFF ram_reg_1674__1_ ( .D(n7226), .CP(wclk), .Q(ram[2985]) );
  DFF ram_reg_1674__0_ ( .D(n7225), .CP(wclk), .Q(ram[2984]) );
  DFF ram_reg_1678__7_ ( .D(n7200), .CP(wclk), .Q(ram[2959]) );
  DFF ram_reg_1678__6_ ( .D(n7199), .CP(wclk), .Q(ram[2958]) );
  DFF ram_reg_1678__5_ ( .D(n7198), .CP(wclk), .Q(ram[2957]) );
  DFF ram_reg_1678__4_ ( .D(n7197), .CP(wclk), .Q(ram[2956]) );
  DFF ram_reg_1678__3_ ( .D(n7196), .CP(wclk), .Q(ram[2955]) );
  DFF ram_reg_1678__2_ ( .D(n7195), .CP(wclk), .Q(ram[2954]) );
  DFF ram_reg_1678__1_ ( .D(n7194), .CP(wclk), .Q(ram[2953]) );
  DFF ram_reg_1678__0_ ( .D(n7193), .CP(wclk), .Q(ram[2952]) );
  DFF ram_reg_1690__7_ ( .D(n7104), .CP(wclk), .Q(ram[2863]) );
  DFF ram_reg_1690__6_ ( .D(n7103), .CP(wclk), .Q(ram[2862]) );
  DFF ram_reg_1690__5_ ( .D(n7102), .CP(wclk), .Q(ram[2861]) );
  DFF ram_reg_1690__4_ ( .D(n7101), .CP(wclk), .Q(ram[2860]) );
  DFF ram_reg_1690__3_ ( .D(n7100), .CP(wclk), .Q(ram[2859]) );
  DFF ram_reg_1690__2_ ( .D(n7099), .CP(wclk), .Q(ram[2858]) );
  DFF ram_reg_1690__1_ ( .D(n7098), .CP(wclk), .Q(ram[2857]) );
  DFF ram_reg_1690__0_ ( .D(n7097), .CP(wclk), .Q(ram[2856]) );
  DFF ram_reg_1698__7_ ( .D(n7040), .CP(wclk), .Q(ram[2799]) );
  DFF ram_reg_1698__6_ ( .D(n7039), .CP(wclk), .Q(ram[2798]) );
  DFF ram_reg_1698__5_ ( .D(n7038), .CP(wclk), .Q(ram[2797]) );
  DFF ram_reg_1698__4_ ( .D(n7037), .CP(wclk), .Q(ram[2796]) );
  DFF ram_reg_1698__3_ ( .D(n7036), .CP(wclk), .Q(ram[2795]) );
  DFF ram_reg_1698__2_ ( .D(n7035), .CP(wclk), .Q(ram[2794]) );
  DFF ram_reg_1698__1_ ( .D(n7034), .CP(wclk), .Q(ram[2793]) );
  DFF ram_reg_1698__0_ ( .D(n7033), .CP(wclk), .Q(ram[2792]) );
  DFF ram_reg_1706__7_ ( .D(n6976), .CP(wclk), .Q(ram[2735]) );
  DFF ram_reg_1706__6_ ( .D(n6975), .CP(wclk), .Q(ram[2734]) );
  DFF ram_reg_1706__5_ ( .D(n6974), .CP(wclk), .Q(ram[2733]) );
  DFF ram_reg_1706__4_ ( .D(n6973), .CP(wclk), .Q(ram[2732]) );
  DFF ram_reg_1706__3_ ( .D(n6972), .CP(wclk), .Q(ram[2731]) );
  DFF ram_reg_1706__2_ ( .D(n6971), .CP(wclk), .Q(ram[2730]) );
  DFF ram_reg_1706__1_ ( .D(n6970), .CP(wclk), .Q(ram[2729]) );
  DFF ram_reg_1706__0_ ( .D(n6969), .CP(wclk), .Q(ram[2728]) );
  DFF ram_reg_1710__7_ ( .D(n6944), .CP(wclk), .Q(ram[2703]) );
  DFF ram_reg_1710__6_ ( .D(n6943), .CP(wclk), .Q(ram[2702]) );
  DFF ram_reg_1710__5_ ( .D(n6942), .CP(wclk), .Q(ram[2701]) );
  DFF ram_reg_1710__4_ ( .D(n6941), .CP(wclk), .Q(ram[2700]) );
  DFF ram_reg_1710__3_ ( .D(n6940), .CP(wclk), .Q(ram[2699]) );
  DFF ram_reg_1710__2_ ( .D(n6939), .CP(wclk), .Q(ram[2698]) );
  DFF ram_reg_1710__1_ ( .D(n6938), .CP(wclk), .Q(ram[2697]) );
  DFF ram_reg_1710__0_ ( .D(n6937), .CP(wclk), .Q(ram[2696]) );
  DFF ram_reg_1714__7_ ( .D(n6912), .CP(wclk), .Q(ram[2671]) );
  DFF ram_reg_1714__6_ ( .D(n6911), .CP(wclk), .Q(ram[2670]) );
  DFF ram_reg_1714__5_ ( .D(n6910), .CP(wclk), .Q(ram[2669]) );
  DFF ram_reg_1714__4_ ( .D(n6909), .CP(wclk), .Q(ram[2668]) );
  DFF ram_reg_1714__3_ ( .D(n6908), .CP(wclk), .Q(ram[2667]) );
  DFF ram_reg_1714__2_ ( .D(n6907), .CP(wclk), .Q(ram[2666]) );
  DFF ram_reg_1714__1_ ( .D(n6906), .CP(wclk), .Q(ram[2665]) );
  DFF ram_reg_1714__0_ ( .D(n6905), .CP(wclk), .Q(ram[2664]) );
  DFF ram_reg_1722__7_ ( .D(n6848), .CP(wclk), .Q(ram[2607]) );
  DFF ram_reg_1722__6_ ( .D(n6847), .CP(wclk), .Q(ram[2606]) );
  DFF ram_reg_1722__5_ ( .D(n6846), .CP(wclk), .Q(ram[2605]) );
  DFF ram_reg_1722__4_ ( .D(n6845), .CP(wclk), .Q(ram[2604]) );
  DFF ram_reg_1722__3_ ( .D(n6844), .CP(wclk), .Q(ram[2603]) );
  DFF ram_reg_1722__2_ ( .D(n6843), .CP(wclk), .Q(ram[2602]) );
  DFF ram_reg_1722__1_ ( .D(n6842), .CP(wclk), .Q(ram[2601]) );
  DFF ram_reg_1722__0_ ( .D(n6841), .CP(wclk), .Q(ram[2600]) );
  DFF ram_reg_1726__7_ ( .D(n6816), .CP(wclk), .Q(ram[2575]) );
  DFF ram_reg_1726__6_ ( .D(n6815), .CP(wclk), .Q(ram[2574]) );
  DFF ram_reg_1726__5_ ( .D(n6814), .CP(wclk), .Q(ram[2573]) );
  DFF ram_reg_1726__4_ ( .D(n6813), .CP(wclk), .Q(ram[2572]) );
  DFF ram_reg_1726__3_ ( .D(n6812), .CP(wclk), .Q(ram[2571]) );
  DFF ram_reg_1726__2_ ( .D(n6811), .CP(wclk), .Q(ram[2570]) );
  DFF ram_reg_1726__1_ ( .D(n6810), .CP(wclk), .Q(ram[2569]) );
  DFF ram_reg_1726__0_ ( .D(n6809), .CP(wclk), .Q(ram[2568]) );
  DFF ram_reg_1738__7_ ( .D(n6720), .CP(wclk), .Q(ram[2479]) );
  DFF ram_reg_1738__6_ ( .D(n6719), .CP(wclk), .Q(ram[2478]) );
  DFF ram_reg_1738__5_ ( .D(n6718), .CP(wclk), .Q(ram[2477]) );
  DFF ram_reg_1738__4_ ( .D(n6717), .CP(wclk), .Q(ram[2476]) );
  DFF ram_reg_1738__3_ ( .D(n6716), .CP(wclk), .Q(ram[2475]) );
  DFF ram_reg_1738__2_ ( .D(n6715), .CP(wclk), .Q(ram[2474]) );
  DFF ram_reg_1738__1_ ( .D(n6714), .CP(wclk), .Q(ram[2473]) );
  DFF ram_reg_1738__0_ ( .D(n6713), .CP(wclk), .Q(ram[2472]) );
  DFF ram_reg_1770__7_ ( .D(n6464), .CP(wclk), .Q(ram[2223]) );
  DFF ram_reg_1770__6_ ( .D(n6463), .CP(wclk), .Q(ram[2222]) );
  DFF ram_reg_1770__5_ ( .D(n6462), .CP(wclk), .Q(ram[2221]) );
  DFF ram_reg_1770__4_ ( .D(n6461), .CP(wclk), .Q(ram[2220]) );
  DFF ram_reg_1770__3_ ( .D(n6460), .CP(wclk), .Q(ram[2219]) );
  DFF ram_reg_1770__2_ ( .D(n6459), .CP(wclk), .Q(ram[2218]) );
  DFF ram_reg_1770__1_ ( .D(n6458), .CP(wclk), .Q(ram[2217]) );
  DFF ram_reg_1770__0_ ( .D(n6457), .CP(wclk), .Q(ram[2216]) );
  DFF ram_reg_1774__7_ ( .D(n6432), .CP(wclk), .Q(ram[2191]) );
  DFF ram_reg_1774__6_ ( .D(n6431), .CP(wclk), .Q(ram[2190]) );
  DFF ram_reg_1774__5_ ( .D(n6430), .CP(wclk), .Q(ram[2189]) );
  DFF ram_reg_1774__4_ ( .D(n6429), .CP(wclk), .Q(ram[2188]) );
  DFF ram_reg_1774__3_ ( .D(n6428), .CP(wclk), .Q(ram[2187]) );
  DFF ram_reg_1774__2_ ( .D(n6427), .CP(wclk), .Q(ram[2186]) );
  DFF ram_reg_1774__1_ ( .D(n6426), .CP(wclk), .Q(ram[2185]) );
  DFF ram_reg_1774__0_ ( .D(n6425), .CP(wclk), .Q(ram[2184]) );
  DFF ram_reg_1786__7_ ( .D(n6336), .CP(wclk), .Q(ram[2095]) );
  DFF ram_reg_1786__6_ ( .D(n6335), .CP(wclk), .Q(ram[2094]) );
  DFF ram_reg_1786__5_ ( .D(n6334), .CP(wclk), .Q(ram[2093]) );
  DFF ram_reg_1786__4_ ( .D(n6333), .CP(wclk), .Q(ram[2092]) );
  DFF ram_reg_1786__3_ ( .D(n6332), .CP(wclk), .Q(ram[2091]) );
  DFF ram_reg_1786__2_ ( .D(n6331), .CP(wclk), .Q(ram[2090]) );
  DFF ram_reg_1786__1_ ( .D(n6330), .CP(wclk), .Q(ram[2089]) );
  DFF ram_reg_1786__0_ ( .D(n6329), .CP(wclk), .Q(ram[2088]) );
  DFF ram_reg_1790__7_ ( .D(n6304), .CP(wclk), .Q(ram[2063]) );
  DFF ram_reg_1790__6_ ( .D(n6303), .CP(wclk), .Q(ram[2062]) );
  DFF ram_reg_1790__5_ ( .D(n6302), .CP(wclk), .Q(ram[2061]) );
  DFF ram_reg_1790__4_ ( .D(n6301), .CP(wclk), .Q(ram[2060]) );
  DFF ram_reg_1790__3_ ( .D(n6300), .CP(wclk), .Q(ram[2059]) );
  DFF ram_reg_1790__2_ ( .D(n6299), .CP(wclk), .Q(ram[2058]) );
  DFF ram_reg_1790__1_ ( .D(n6298), .CP(wclk), .Q(ram[2057]) );
  DFF ram_reg_1790__0_ ( .D(n6297), .CP(wclk), .Q(ram[2056]) );
  DFF ram_reg_1834__7_ ( .D(n5952), .CP(wclk), .Q(ram[1711]) );
  DFF ram_reg_1834__6_ ( .D(n5951), .CP(wclk), .Q(ram[1710]) );
  DFF ram_reg_1834__5_ ( .D(n5950), .CP(wclk), .Q(ram[1709]) );
  DFF ram_reg_1834__4_ ( .D(n5949), .CP(wclk), .Q(ram[1708]) );
  DFF ram_reg_1834__3_ ( .D(n5948), .CP(wclk), .Q(ram[1707]) );
  DFF ram_reg_1834__2_ ( .D(n5947), .CP(wclk), .Q(ram[1706]) );
  DFF ram_reg_1834__1_ ( .D(n5946), .CP(wclk), .Q(ram[1705]) );
  DFF ram_reg_1834__0_ ( .D(n5945), .CP(wclk), .Q(ram[1704]) );
  DFF ram_reg_1850__7_ ( .D(n5824), .CP(wclk), .Q(ram[1583]) );
  DFF ram_reg_1850__6_ ( .D(n5823), .CP(wclk), .Q(ram[1582]) );
  DFF ram_reg_1850__5_ ( .D(n5822), .CP(wclk), .Q(ram[1581]) );
  DFF ram_reg_1850__4_ ( .D(n5821), .CP(wclk), .Q(ram[1580]) );
  DFF ram_reg_1850__3_ ( .D(n5820), .CP(wclk), .Q(ram[1579]) );
  DFF ram_reg_1850__2_ ( .D(n5819), .CP(wclk), .Q(ram[1578]) );
  DFF ram_reg_1850__1_ ( .D(n5818), .CP(wclk), .Q(ram[1577]) );
  DFF ram_reg_1850__0_ ( .D(n5817), .CP(wclk), .Q(ram[1576]) );
  DFF ram_reg_1854__7_ ( .D(n5792), .CP(wclk), .Q(ram[1551]) );
  DFF ram_reg_1854__6_ ( .D(n5791), .CP(wclk), .Q(ram[1550]) );
  DFF ram_reg_1854__5_ ( .D(n5790), .CP(wclk), .Q(ram[1549]) );
  DFF ram_reg_1854__4_ ( .D(n5789), .CP(wclk), .Q(ram[1548]) );
  DFF ram_reg_1854__3_ ( .D(n5788), .CP(wclk), .Q(ram[1547]) );
  DFF ram_reg_1854__2_ ( .D(n5787), .CP(wclk), .Q(ram[1546]) );
  DFF ram_reg_1854__1_ ( .D(n5786), .CP(wclk), .Q(ram[1545]) );
  DFF ram_reg_1854__0_ ( .D(n5785), .CP(wclk), .Q(ram[1544]) );
  DFF ram_reg_1930__7_ ( .D(n5184), .CP(wclk), .Q(ram[943]) );
  DFF ram_reg_1930__6_ ( .D(n5183), .CP(wclk), .Q(ram[942]) );
  DFF ram_reg_1930__5_ ( .D(n5182), .CP(wclk), .Q(ram[941]) );
  DFF ram_reg_1930__4_ ( .D(n5181), .CP(wclk), .Q(ram[940]) );
  DFF ram_reg_1930__3_ ( .D(n5180), .CP(wclk), .Q(ram[939]) );
  DFF ram_reg_1930__2_ ( .D(n5179), .CP(wclk), .Q(ram[938]) );
  DFF ram_reg_1930__1_ ( .D(n5178), .CP(wclk), .Q(ram[937]) );
  DFF ram_reg_1930__0_ ( .D(n5177), .CP(wclk), .Q(ram[936]) );
  DFF ram_reg_1934__7_ ( .D(n5152), .CP(wclk), .Q(ram[911]) );
  DFF ram_reg_1934__6_ ( .D(n5151), .CP(wclk), .Q(ram[910]) );
  DFF ram_reg_1934__5_ ( .D(n5150), .CP(wclk), .Q(ram[909]) );
  DFF ram_reg_1934__4_ ( .D(n5149), .CP(wclk), .Q(ram[908]) );
  DFF ram_reg_1934__3_ ( .D(n5148), .CP(wclk), .Q(ram[907]) );
  DFF ram_reg_1934__2_ ( .D(n5147), .CP(wclk), .Q(ram[906]) );
  DFF ram_reg_1934__1_ ( .D(n5146), .CP(wclk), .Q(ram[905]) );
  DFF ram_reg_1934__0_ ( .D(n5145), .CP(wclk), .Q(ram[904]) );
  DFF ram_reg_1946__7_ ( .D(n5056), .CP(wclk), .Q(ram[815]) );
  DFF ram_reg_1946__6_ ( .D(n5055), .CP(wclk), .Q(ram[814]) );
  DFF ram_reg_1946__5_ ( .D(n5054), .CP(wclk), .Q(ram[813]) );
  DFF ram_reg_1946__4_ ( .D(n5053), .CP(wclk), .Q(ram[812]) );
  DFF ram_reg_1946__3_ ( .D(n5052), .CP(wclk), .Q(ram[811]) );
  DFF ram_reg_1946__2_ ( .D(n5051), .CP(wclk), .Q(ram[810]) );
  DFF ram_reg_1946__1_ ( .D(n5050), .CP(wclk), .Q(ram[809]) );
  DFF ram_reg_1946__0_ ( .D(n5049), .CP(wclk), .Q(ram[808]) );
  DFF ram_reg_1950__7_ ( .D(n5024), .CP(wclk), .Q(ram[783]) );
  DFF ram_reg_1950__6_ ( .D(n5023), .CP(wclk), .Q(ram[782]) );
  DFF ram_reg_1950__5_ ( .D(n5022), .CP(wclk), .Q(ram[781]) );
  DFF ram_reg_1950__4_ ( .D(n5021), .CP(wclk), .Q(ram[780]) );
  DFF ram_reg_1950__3_ ( .D(n5020), .CP(wclk), .Q(ram[779]) );
  DFF ram_reg_1950__2_ ( .D(n5019), .CP(wclk), .Q(ram[778]) );
  DFF ram_reg_1950__1_ ( .D(n5018), .CP(wclk), .Q(ram[777]) );
  DFF ram_reg_1950__0_ ( .D(n5017), .CP(wclk), .Q(ram[776]) );
  DFF ram_reg_1954__7_ ( .D(n4992), .CP(wclk), .Q(ram[751]) );
  DFF ram_reg_1954__6_ ( .D(n4991), .CP(wclk), .Q(ram[750]) );
  DFF ram_reg_1954__5_ ( .D(n4990), .CP(wclk), .Q(ram[749]) );
  DFF ram_reg_1954__4_ ( .D(n4989), .CP(wclk), .Q(ram[748]) );
  DFF ram_reg_1954__3_ ( .D(n4988), .CP(wclk), .Q(ram[747]) );
  DFF ram_reg_1954__2_ ( .D(n4987), .CP(wclk), .Q(ram[746]) );
  DFF ram_reg_1954__1_ ( .D(n4986), .CP(wclk), .Q(ram[745]) );
  DFF ram_reg_1954__0_ ( .D(n4985), .CP(wclk), .Q(ram[744]) );
  DFF ram_reg_1962__7_ ( .D(n4928), .CP(wclk), .Q(ram[687]) );
  DFF ram_reg_1962__6_ ( .D(n4927), .CP(wclk), .Q(ram[686]) );
  DFF ram_reg_1962__5_ ( .D(n4926), .CP(wclk), .Q(ram[685]) );
  DFF ram_reg_1962__4_ ( .D(n4925), .CP(wclk), .Q(ram[684]) );
  DFF ram_reg_1962__3_ ( .D(n4924), .CP(wclk), .Q(ram[683]) );
  DFF ram_reg_1962__2_ ( .D(n4923), .CP(wclk), .Q(ram[682]) );
  DFF ram_reg_1962__1_ ( .D(n4922), .CP(wclk), .Q(ram[681]) );
  DFF ram_reg_1962__0_ ( .D(n4921), .CP(wclk), .Q(ram[680]) );
  DFF ram_reg_1966__7_ ( .D(n4896), .CP(wclk), .Q(ram[655]) );
  DFF ram_reg_1966__6_ ( .D(n4895), .CP(wclk), .Q(ram[654]) );
  DFF ram_reg_1966__5_ ( .D(n4894), .CP(wclk), .Q(ram[653]) );
  DFF ram_reg_1966__4_ ( .D(n4893), .CP(wclk), .Q(ram[652]) );
  DFF ram_reg_1966__3_ ( .D(n4892), .CP(wclk), .Q(ram[651]) );
  DFF ram_reg_1966__2_ ( .D(n4891), .CP(wclk), .Q(ram[650]) );
  DFF ram_reg_1966__1_ ( .D(n4890), .CP(wclk), .Q(ram[649]) );
  DFF ram_reg_1966__0_ ( .D(n4889), .CP(wclk), .Q(ram[648]) );
  DFF ram_reg_1970__7_ ( .D(n4864), .CP(wclk), .Q(ram[623]) );
  DFF ram_reg_1970__6_ ( .D(n4863), .CP(wclk), .Q(ram[622]) );
  DFF ram_reg_1970__5_ ( .D(n4862), .CP(wclk), .Q(ram[621]) );
  DFF ram_reg_1970__4_ ( .D(n4861), .CP(wclk), .Q(ram[620]) );
  DFF ram_reg_1970__3_ ( .D(n4860), .CP(wclk), .Q(ram[619]) );
  DFF ram_reg_1970__2_ ( .D(n4859), .CP(wclk), .Q(ram[618]) );
  DFF ram_reg_1970__1_ ( .D(n4858), .CP(wclk), .Q(ram[617]) );
  DFF ram_reg_1970__0_ ( .D(n4857), .CP(wclk), .Q(ram[616]) );
  DFF ram_reg_1978__7_ ( .D(n4800), .CP(wclk), .Q(ram[559]) );
  DFF ram_reg_1978__6_ ( .D(n4799), .CP(wclk), .Q(ram[558]) );
  DFF ram_reg_1978__5_ ( .D(n4798), .CP(wclk), .Q(ram[557]) );
  DFF ram_reg_1978__4_ ( .D(n4797), .CP(wclk), .Q(ram[556]) );
  DFF ram_reg_1978__3_ ( .D(n4796), .CP(wclk), .Q(ram[555]) );
  DFF ram_reg_1978__2_ ( .D(n4795), .CP(wclk), .Q(ram[554]) );
  DFF ram_reg_1978__1_ ( .D(n4794), .CP(wclk), .Q(ram[553]) );
  DFF ram_reg_1978__0_ ( .D(n4793), .CP(wclk), .Q(ram[552]) );
  DFF ram_reg_1982__7_ ( .D(n4768), .CP(wclk), .Q(ram[527]) );
  DFF ram_reg_1982__6_ ( .D(n4767), .CP(wclk), .Q(ram[526]) );
  DFF ram_reg_1982__5_ ( .D(n4766), .CP(wclk), .Q(ram[525]) );
  DFF ram_reg_1982__4_ ( .D(n4765), .CP(wclk), .Q(ram[524]) );
  DFF ram_reg_1982__3_ ( .D(n4764), .CP(wclk), .Q(ram[523]) );
  DFF ram_reg_1982__2_ ( .D(n4763), .CP(wclk), .Q(ram[522]) );
  DFF ram_reg_1982__1_ ( .D(n4762), .CP(wclk), .Q(ram[521]) );
  DFF ram_reg_1982__0_ ( .D(n4761), .CP(wclk), .Q(ram[520]) );
  DFF ram_reg_1994__7_ ( .D(n4672), .CP(wclk), .Q(ram[431]) );
  DFF ram_reg_1994__6_ ( .D(n4671), .CP(wclk), .Q(ram[430]) );
  DFF ram_reg_1994__5_ ( .D(n4670), .CP(wclk), .Q(ram[429]) );
  DFF ram_reg_1994__4_ ( .D(n4669), .CP(wclk), .Q(ram[428]) );
  DFF ram_reg_1994__3_ ( .D(n4668), .CP(wclk), .Q(ram[427]) );
  DFF ram_reg_1994__2_ ( .D(n4667), .CP(wclk), .Q(ram[426]) );
  DFF ram_reg_1994__1_ ( .D(n4666), .CP(wclk), .Q(ram[425]) );
  DFF ram_reg_1994__0_ ( .D(n4665), .CP(wclk), .Q(ram[424]) );
  DFF ram_reg_1998__7_ ( .D(n4640), .CP(wclk), .Q(ram[399]) );
  DFF ram_reg_1998__6_ ( .D(n4639), .CP(wclk), .Q(ram[398]) );
  DFF ram_reg_1998__5_ ( .D(n4638), .CP(wclk), .Q(ram[397]) );
  DFF ram_reg_1998__4_ ( .D(n4637), .CP(wclk), .Q(ram[396]) );
  DFF ram_reg_1998__3_ ( .D(n4636), .CP(wclk), .Q(ram[395]) );
  DFF ram_reg_1998__2_ ( .D(n4635), .CP(wclk), .Q(ram[394]) );
  DFF ram_reg_1998__1_ ( .D(n4634), .CP(wclk), .Q(ram[393]) );
  DFF ram_reg_1998__0_ ( .D(n4633), .CP(wclk), .Q(ram[392]) );
  DFF ram_reg_2010__7_ ( .D(n4544), .CP(wclk), .Q(ram[303]) );
  DFF ram_reg_2010__6_ ( .D(n4543), .CP(wclk), .Q(ram[302]) );
  DFF ram_reg_2010__5_ ( .D(n4542), .CP(wclk), .Q(ram[301]) );
  DFF ram_reg_2010__4_ ( .D(n4541), .CP(wclk), .Q(ram[300]) );
  DFF ram_reg_2010__3_ ( .D(n4540), .CP(wclk), .Q(ram[299]) );
  DFF ram_reg_2010__2_ ( .D(n4539), .CP(wclk), .Q(ram[298]) );
  DFF ram_reg_2010__1_ ( .D(n4538), .CP(wclk), .Q(ram[297]) );
  DFF ram_reg_2010__0_ ( .D(n4537), .CP(wclk), .Q(ram[296]) );
  DFF ram_reg_2026__7_ ( .D(n4416), .CP(wclk), .Q(ram[175]) );
  DFF ram_reg_2026__6_ ( .D(n4415), .CP(wclk), .Q(ram[174]) );
  DFF ram_reg_2026__5_ ( .D(n4414), .CP(wclk), .Q(ram[173]) );
  DFF ram_reg_2026__4_ ( .D(n4413), .CP(wclk), .Q(ram[172]) );
  DFF ram_reg_2026__3_ ( .D(n4412), .CP(wclk), .Q(ram[171]) );
  DFF ram_reg_2026__2_ ( .D(n4411), .CP(wclk), .Q(ram[170]) );
  DFF ram_reg_2026__1_ ( .D(n4410), .CP(wclk), .Q(ram[169]) );
  DFF ram_reg_2026__0_ ( .D(n4409), .CP(wclk), .Q(ram[168]) );
  DFF ram_reg_2030__7_ ( .D(n4384), .CP(wclk), .Q(ram[143]) );
  DFF ram_reg_2030__6_ ( .D(n4383), .CP(wclk), .Q(ram[142]) );
  DFF ram_reg_2030__5_ ( .D(n4382), .CP(wclk), .Q(ram[141]) );
  DFF ram_reg_2030__4_ ( .D(n4381), .CP(wclk), .Q(ram[140]) );
  DFF ram_reg_2030__3_ ( .D(n4380), .CP(wclk), .Q(ram[139]) );
  DFF ram_reg_2030__2_ ( .D(n4379), .CP(wclk), .Q(ram[138]) );
  DFF ram_reg_2030__1_ ( .D(n4378), .CP(wclk), .Q(ram[137]) );
  DFF ram_reg_2030__0_ ( .D(n4377), .CP(wclk), .Q(ram[136]) );
  DFF ram_reg_2034__7_ ( .D(n4352), .CP(wclk), .Q(ram[111]) );
  DFF ram_reg_2034__6_ ( .D(n4351), .CP(wclk), .Q(ram[110]) );
  DFF ram_reg_2034__5_ ( .D(n4350), .CP(wclk), .Q(ram[109]) );
  DFF ram_reg_2034__4_ ( .D(n4349), .CP(wclk), .Q(ram[108]) );
  DFF ram_reg_2034__3_ ( .D(n4348), .CP(wclk), .Q(ram[107]) );
  DFF ram_reg_2034__2_ ( .D(n4347), .CP(wclk), .Q(ram[106]) );
  DFF ram_reg_2034__1_ ( .D(n4346), .CP(wclk), .Q(ram[105]) );
  DFF ram_reg_2034__0_ ( .D(n4345), .CP(wclk), .Q(ram[104]) );
  DFF ram_reg_2042__7_ ( .D(n4288), .CP(wclk), .Q(ram[47]) );
  DFF ram_reg_2042__6_ ( .D(n4287), .CP(wclk), .Q(ram[46]) );
  DFF ram_reg_2042__5_ ( .D(n4286), .CP(wclk), .Q(ram[45]) );
  DFF ram_reg_2042__4_ ( .D(n4285), .CP(wclk), .Q(ram[44]) );
  DFF ram_reg_2042__3_ ( .D(n4284), .CP(wclk), .Q(ram[43]) );
  DFF ram_reg_2042__2_ ( .D(n4283), .CP(wclk), .Q(ram[42]) );
  DFF ram_reg_2042__1_ ( .D(n4282), .CP(wclk), .Q(ram[41]) );
  DFF ram_reg_2042__0_ ( .D(n4281), .CP(wclk), .Q(ram[40]) );
  DFF ram_reg_2046__7_ ( .D(n4256), .CP(wclk), .Q(ram[15]) );
  DFF ram_reg_2046__6_ ( .D(n4255), .CP(wclk), .Q(ram[14]) );
  DFF ram_reg_2046__5_ ( .D(n4254), .CP(wclk), .Q(ram[13]) );
  DFF ram_reg_2046__4_ ( .D(n4253), .CP(wclk), .Q(ram[12]) );
  DFF ram_reg_2046__3_ ( .D(n4252), .CP(wclk), .Q(ram[11]) );
  DFF ram_reg_2046__2_ ( .D(n4251), .CP(wclk), .Q(ram[10]) );
  DFF ram_reg_2046__1_ ( .D(n4250), .CP(wclk), .Q(ram[9]) );
  DFF ram_reg_2046__0_ ( .D(n4249), .CP(wclk), .Q(ram[8]) );
  DFF ram_reg_9__7_ ( .D(n20552), .CP(wclk), .Q(ram[16311]) );
  DFF ram_reg_9__6_ ( .D(n20551), .CP(wclk), .Q(ram[16310]) );
  DFF ram_reg_9__5_ ( .D(n20550), .CP(wclk), .Q(ram[16309]) );
  DFF ram_reg_9__4_ ( .D(n20549), .CP(wclk), .Q(ram[16308]) );
  DFF ram_reg_9__3_ ( .D(n20548), .CP(wclk), .Q(ram[16307]) );
  DFF ram_reg_9__2_ ( .D(n20547), .CP(wclk), .Q(ram[16306]) );
  DFF ram_reg_9__1_ ( .D(n20546), .CP(wclk), .Q(ram[16305]) );
  DFF ram_reg_9__0_ ( .D(n20545), .CP(wclk), .Q(ram[16304]) );
  DFF ram_reg_41__7_ ( .D(n20296), .CP(wclk), .Q(ram[16055]) );
  DFF ram_reg_41__6_ ( .D(n20295), .CP(wclk), .Q(ram[16054]) );
  DFF ram_reg_41__5_ ( .D(n20294), .CP(wclk), .Q(ram[16053]) );
  DFF ram_reg_41__4_ ( .D(n20293), .CP(wclk), .Q(ram[16052]) );
  DFF ram_reg_41__3_ ( .D(n20292), .CP(wclk), .Q(ram[16051]) );
  DFF ram_reg_41__2_ ( .D(n20291), .CP(wclk), .Q(ram[16050]) );
  DFF ram_reg_41__1_ ( .D(n20290), .CP(wclk), .Q(ram[16049]) );
  DFF ram_reg_41__0_ ( .D(n20289), .CP(wclk), .Q(ram[16048]) );
  DFF ram_reg_45__7_ ( .D(n20264), .CP(wclk), .Q(ram[16023]) );
  DFF ram_reg_45__6_ ( .D(n20263), .CP(wclk), .Q(ram[16022]) );
  DFF ram_reg_45__5_ ( .D(n20262), .CP(wclk), .Q(ram[16021]) );
  DFF ram_reg_45__4_ ( .D(n20261), .CP(wclk), .Q(ram[16020]) );
  DFF ram_reg_45__3_ ( .D(n20260), .CP(wclk), .Q(ram[16019]) );
  DFF ram_reg_45__2_ ( .D(n20259), .CP(wclk), .Q(ram[16018]) );
  DFF ram_reg_45__1_ ( .D(n20258), .CP(wclk), .Q(ram[16017]) );
  DFF ram_reg_45__0_ ( .D(n20257), .CP(wclk), .Q(ram[16016]) );
  DFF ram_reg_57__7_ ( .D(n20168), .CP(wclk), .Q(ram[15927]) );
  DFF ram_reg_57__6_ ( .D(n20167), .CP(wclk), .Q(ram[15926]) );
  DFF ram_reg_57__5_ ( .D(n20166), .CP(wclk), .Q(ram[15925]) );
  DFF ram_reg_57__4_ ( .D(n20165), .CP(wclk), .Q(ram[15924]) );
  DFF ram_reg_57__3_ ( .D(n20164), .CP(wclk), .Q(ram[15923]) );
  DFF ram_reg_57__2_ ( .D(n20163), .CP(wclk), .Q(ram[15922]) );
  DFF ram_reg_57__1_ ( .D(n20162), .CP(wclk), .Q(ram[15921]) );
  DFF ram_reg_57__0_ ( .D(n20161), .CP(wclk), .Q(ram[15920]) );
  DFF ram_reg_61__7_ ( .D(n20136), .CP(wclk), .Q(ram[15895]) );
  DFF ram_reg_61__6_ ( .D(n20135), .CP(wclk), .Q(ram[15894]) );
  DFF ram_reg_61__5_ ( .D(n20134), .CP(wclk), .Q(ram[15893]) );
  DFF ram_reg_61__4_ ( .D(n20133), .CP(wclk), .Q(ram[15892]) );
  DFF ram_reg_61__3_ ( .D(n20132), .CP(wclk), .Q(ram[15891]) );
  DFF ram_reg_61__2_ ( .D(n20131), .CP(wclk), .Q(ram[15890]) );
  DFF ram_reg_61__1_ ( .D(n20130), .CP(wclk), .Q(ram[15889]) );
  DFF ram_reg_61__0_ ( .D(n20129), .CP(wclk), .Q(ram[15888]) );
  DFF ram_reg_129__7_ ( .D(n19592), .CP(wclk), .Q(ram[15351]) );
  DFF ram_reg_129__6_ ( .D(n19591), .CP(wclk), .Q(ram[15350]) );
  DFF ram_reg_129__5_ ( .D(n19590), .CP(wclk), .Q(ram[15349]) );
  DFF ram_reg_129__4_ ( .D(n19589), .CP(wclk), .Q(ram[15348]) );
  DFF ram_reg_129__3_ ( .D(n19588), .CP(wclk), .Q(ram[15347]) );
  DFF ram_reg_129__2_ ( .D(n19587), .CP(wclk), .Q(ram[15346]) );
  DFF ram_reg_129__1_ ( .D(n19586), .CP(wclk), .Q(ram[15345]) );
  DFF ram_reg_129__0_ ( .D(n19585), .CP(wclk), .Q(ram[15344]) );
  DFF ram_reg_137__7_ ( .D(n19528), .CP(wclk), .Q(ram[15287]) );
  DFF ram_reg_137__6_ ( .D(n19527), .CP(wclk), .Q(ram[15286]) );
  DFF ram_reg_137__5_ ( .D(n19526), .CP(wclk), .Q(ram[15285]) );
  DFF ram_reg_137__4_ ( .D(n19525), .CP(wclk), .Q(ram[15284]) );
  DFF ram_reg_137__3_ ( .D(n19524), .CP(wclk), .Q(ram[15283]) );
  DFF ram_reg_137__2_ ( .D(n19523), .CP(wclk), .Q(ram[15282]) );
  DFF ram_reg_137__1_ ( .D(n19522), .CP(wclk), .Q(ram[15281]) );
  DFF ram_reg_137__0_ ( .D(n19521), .CP(wclk), .Q(ram[15280]) );
  DFF ram_reg_141__7_ ( .D(n19496), .CP(wclk), .Q(ram[15255]) );
  DFF ram_reg_141__6_ ( .D(n19495), .CP(wclk), .Q(ram[15254]) );
  DFF ram_reg_141__5_ ( .D(n19494), .CP(wclk), .Q(ram[15253]) );
  DFF ram_reg_141__4_ ( .D(n19493), .CP(wclk), .Q(ram[15252]) );
  DFF ram_reg_141__3_ ( .D(n19492), .CP(wclk), .Q(ram[15251]) );
  DFF ram_reg_141__2_ ( .D(n19491), .CP(wclk), .Q(ram[15250]) );
  DFF ram_reg_141__1_ ( .D(n19490), .CP(wclk), .Q(ram[15249]) );
  DFF ram_reg_141__0_ ( .D(n19489), .CP(wclk), .Q(ram[15248]) );
  DFF ram_reg_153__7_ ( .D(n19400), .CP(wclk), .Q(ram[15159]) );
  DFF ram_reg_153__6_ ( .D(n19399), .CP(wclk), .Q(ram[15158]) );
  DFF ram_reg_153__5_ ( .D(n19398), .CP(wclk), .Q(ram[15157]) );
  DFF ram_reg_153__4_ ( .D(n19397), .CP(wclk), .Q(ram[15156]) );
  DFF ram_reg_153__3_ ( .D(n19396), .CP(wclk), .Q(ram[15155]) );
  DFF ram_reg_153__2_ ( .D(n19395), .CP(wclk), .Q(ram[15154]) );
  DFF ram_reg_153__1_ ( .D(n19394), .CP(wclk), .Q(ram[15153]) );
  DFF ram_reg_153__0_ ( .D(n19393), .CP(wclk), .Q(ram[15152]) );
  DFF ram_reg_157__7_ ( .D(n19368), .CP(wclk), .Q(ram[15127]) );
  DFF ram_reg_157__6_ ( .D(n19367), .CP(wclk), .Q(ram[15126]) );
  DFF ram_reg_157__5_ ( .D(n19366), .CP(wclk), .Q(ram[15125]) );
  DFF ram_reg_157__4_ ( .D(n19365), .CP(wclk), .Q(ram[15124]) );
  DFF ram_reg_157__3_ ( .D(n19364), .CP(wclk), .Q(ram[15123]) );
  DFF ram_reg_157__2_ ( .D(n19363), .CP(wclk), .Q(ram[15122]) );
  DFF ram_reg_157__1_ ( .D(n19362), .CP(wclk), .Q(ram[15121]) );
  DFF ram_reg_157__0_ ( .D(n19361), .CP(wclk), .Q(ram[15120]) );
  DFF ram_reg_161__7_ ( .D(n19336), .CP(wclk), .Q(ram[15095]) );
  DFF ram_reg_161__6_ ( .D(n19335), .CP(wclk), .Q(ram[15094]) );
  DFF ram_reg_161__5_ ( .D(n19334), .CP(wclk), .Q(ram[15093]) );
  DFF ram_reg_161__4_ ( .D(n19333), .CP(wclk), .Q(ram[15092]) );
  DFF ram_reg_161__3_ ( .D(n19332), .CP(wclk), .Q(ram[15091]) );
  DFF ram_reg_161__2_ ( .D(n19331), .CP(wclk), .Q(ram[15090]) );
  DFF ram_reg_161__1_ ( .D(n19330), .CP(wclk), .Q(ram[15089]) );
  DFF ram_reg_161__0_ ( .D(n19329), .CP(wclk), .Q(ram[15088]) );
  DFF ram_reg_169__7_ ( .D(n19272), .CP(wclk), .Q(ram[15031]) );
  DFF ram_reg_169__6_ ( .D(n19271), .CP(wclk), .Q(ram[15030]) );
  DFF ram_reg_169__5_ ( .D(n19270), .CP(wclk), .Q(ram[15029]) );
  DFF ram_reg_169__4_ ( .D(n19269), .CP(wclk), .Q(ram[15028]) );
  DFF ram_reg_169__3_ ( .D(n19268), .CP(wclk), .Q(ram[15027]) );
  DFF ram_reg_169__2_ ( .D(n19267), .CP(wclk), .Q(ram[15026]) );
  DFF ram_reg_169__1_ ( .D(n19266), .CP(wclk), .Q(ram[15025]) );
  DFF ram_reg_169__0_ ( .D(n19265), .CP(wclk), .Q(ram[15024]) );
  DFF ram_reg_173__7_ ( .D(n19240), .CP(wclk), .Q(ram[14999]) );
  DFF ram_reg_173__6_ ( .D(n19239), .CP(wclk), .Q(ram[14998]) );
  DFF ram_reg_173__5_ ( .D(n19238), .CP(wclk), .Q(ram[14997]) );
  DFF ram_reg_173__4_ ( .D(n19237), .CP(wclk), .Q(ram[14996]) );
  DFF ram_reg_173__3_ ( .D(n19236), .CP(wclk), .Q(ram[14995]) );
  DFF ram_reg_173__2_ ( .D(n19235), .CP(wclk), .Q(ram[14994]) );
  DFF ram_reg_173__1_ ( .D(n19234), .CP(wclk), .Q(ram[14993]) );
  DFF ram_reg_173__0_ ( .D(n19233), .CP(wclk), .Q(ram[14992]) );
  DFF ram_reg_177__7_ ( .D(n19208), .CP(wclk), .Q(ram[14967]) );
  DFF ram_reg_177__6_ ( .D(n19207), .CP(wclk), .Q(ram[14966]) );
  DFF ram_reg_177__5_ ( .D(n19206), .CP(wclk), .Q(ram[14965]) );
  DFF ram_reg_177__4_ ( .D(n19205), .CP(wclk), .Q(ram[14964]) );
  DFF ram_reg_177__3_ ( .D(n19204), .CP(wclk), .Q(ram[14963]) );
  DFF ram_reg_177__2_ ( .D(n19203), .CP(wclk), .Q(ram[14962]) );
  DFF ram_reg_177__1_ ( .D(n19202), .CP(wclk), .Q(ram[14961]) );
  DFF ram_reg_177__0_ ( .D(n19201), .CP(wclk), .Q(ram[14960]) );
  DFF ram_reg_185__7_ ( .D(n19144), .CP(wclk), .Q(ram[14903]) );
  DFF ram_reg_185__6_ ( .D(n19143), .CP(wclk), .Q(ram[14902]) );
  DFF ram_reg_185__5_ ( .D(n19142), .CP(wclk), .Q(ram[14901]) );
  DFF ram_reg_185__4_ ( .D(n19141), .CP(wclk), .Q(ram[14900]) );
  DFF ram_reg_185__3_ ( .D(n19140), .CP(wclk), .Q(ram[14899]) );
  DFF ram_reg_185__2_ ( .D(n19139), .CP(wclk), .Q(ram[14898]) );
  DFF ram_reg_185__1_ ( .D(n19138), .CP(wclk), .Q(ram[14897]) );
  DFF ram_reg_185__0_ ( .D(n19137), .CP(wclk), .Q(ram[14896]) );
  DFF ram_reg_189__7_ ( .D(n19112), .CP(wclk), .Q(ram[14871]) );
  DFF ram_reg_189__6_ ( .D(n19111), .CP(wclk), .Q(ram[14870]) );
  DFF ram_reg_189__5_ ( .D(n19110), .CP(wclk), .Q(ram[14869]) );
  DFF ram_reg_189__4_ ( .D(n19109), .CP(wclk), .Q(ram[14868]) );
  DFF ram_reg_189__3_ ( .D(n19108), .CP(wclk), .Q(ram[14867]) );
  DFF ram_reg_189__2_ ( .D(n19107), .CP(wclk), .Q(ram[14866]) );
  DFF ram_reg_189__1_ ( .D(n19106), .CP(wclk), .Q(ram[14865]) );
  DFF ram_reg_189__0_ ( .D(n19105), .CP(wclk), .Q(ram[14864]) );
  DFF ram_reg_201__7_ ( .D(n19016), .CP(wclk), .Q(ram[14775]) );
  DFF ram_reg_201__6_ ( .D(n19015), .CP(wclk), .Q(ram[14774]) );
  DFF ram_reg_201__5_ ( .D(n19014), .CP(wclk), .Q(ram[14773]) );
  DFF ram_reg_201__4_ ( .D(n19013), .CP(wclk), .Q(ram[14772]) );
  DFF ram_reg_201__3_ ( .D(n19012), .CP(wclk), .Q(ram[14771]) );
  DFF ram_reg_201__2_ ( .D(n19011), .CP(wclk), .Q(ram[14770]) );
  DFF ram_reg_201__1_ ( .D(n19010), .CP(wclk), .Q(ram[14769]) );
  DFF ram_reg_201__0_ ( .D(n19009), .CP(wclk), .Q(ram[14768]) );
  DFF ram_reg_205__7_ ( .D(n18984), .CP(wclk), .Q(ram[14743]) );
  DFF ram_reg_205__6_ ( .D(n18983), .CP(wclk), .Q(ram[14742]) );
  DFF ram_reg_205__5_ ( .D(n18982), .CP(wclk), .Q(ram[14741]) );
  DFF ram_reg_205__4_ ( .D(n18981), .CP(wclk), .Q(ram[14740]) );
  DFF ram_reg_205__3_ ( .D(n18980), .CP(wclk), .Q(ram[14739]) );
  DFF ram_reg_205__2_ ( .D(n18979), .CP(wclk), .Q(ram[14738]) );
  DFF ram_reg_205__1_ ( .D(n18978), .CP(wclk), .Q(ram[14737]) );
  DFF ram_reg_205__0_ ( .D(n18977), .CP(wclk), .Q(ram[14736]) );
  DFF ram_reg_217__7_ ( .D(n18888), .CP(wclk), .Q(ram[14647]) );
  DFF ram_reg_217__6_ ( .D(n18887), .CP(wclk), .Q(ram[14646]) );
  DFF ram_reg_217__5_ ( .D(n18886), .CP(wclk), .Q(ram[14645]) );
  DFF ram_reg_217__4_ ( .D(n18885), .CP(wclk), .Q(ram[14644]) );
  DFF ram_reg_217__3_ ( .D(n18884), .CP(wclk), .Q(ram[14643]) );
  DFF ram_reg_217__2_ ( .D(n18883), .CP(wclk), .Q(ram[14642]) );
  DFF ram_reg_217__1_ ( .D(n18882), .CP(wclk), .Q(ram[14641]) );
  DFF ram_reg_217__0_ ( .D(n18881), .CP(wclk), .Q(ram[14640]) );
  DFF ram_reg_221__7_ ( .D(n18856), .CP(wclk), .Q(ram[14615]) );
  DFF ram_reg_221__6_ ( .D(n18855), .CP(wclk), .Q(ram[14614]) );
  DFF ram_reg_221__5_ ( .D(n18854), .CP(wclk), .Q(ram[14613]) );
  DFF ram_reg_221__4_ ( .D(n18853), .CP(wclk), .Q(ram[14612]) );
  DFF ram_reg_221__3_ ( .D(n18852), .CP(wclk), .Q(ram[14611]) );
  DFF ram_reg_221__2_ ( .D(n18851), .CP(wclk), .Q(ram[14610]) );
  DFF ram_reg_221__1_ ( .D(n18850), .CP(wclk), .Q(ram[14609]) );
  DFF ram_reg_221__0_ ( .D(n18849), .CP(wclk), .Q(ram[14608]) );
  DFF ram_reg_225__7_ ( .D(n18824), .CP(wclk), .Q(ram[14583]) );
  DFF ram_reg_225__6_ ( .D(n18823), .CP(wclk), .Q(ram[14582]) );
  DFF ram_reg_225__5_ ( .D(n18822), .CP(wclk), .Q(ram[14581]) );
  DFF ram_reg_225__4_ ( .D(n18821), .CP(wclk), .Q(ram[14580]) );
  DFF ram_reg_225__3_ ( .D(n18820), .CP(wclk), .Q(ram[14579]) );
  DFF ram_reg_225__2_ ( .D(n18819), .CP(wclk), .Q(ram[14578]) );
  DFF ram_reg_225__1_ ( .D(n18818), .CP(wclk), .Q(ram[14577]) );
  DFF ram_reg_225__0_ ( .D(n18817), .CP(wclk), .Q(ram[14576]) );
  DFF ram_reg_233__7_ ( .D(n18760), .CP(wclk), .Q(ram[14519]) );
  DFF ram_reg_233__6_ ( .D(n18759), .CP(wclk), .Q(ram[14518]) );
  DFF ram_reg_233__5_ ( .D(n18758), .CP(wclk), .Q(ram[14517]) );
  DFF ram_reg_233__4_ ( .D(n18757), .CP(wclk), .Q(ram[14516]) );
  DFF ram_reg_233__3_ ( .D(n18756), .CP(wclk), .Q(ram[14515]) );
  DFF ram_reg_233__2_ ( .D(n18755), .CP(wclk), .Q(ram[14514]) );
  DFF ram_reg_233__1_ ( .D(n18754), .CP(wclk), .Q(ram[14513]) );
  DFF ram_reg_233__0_ ( .D(n18753), .CP(wclk), .Q(ram[14512]) );
  DFF ram_reg_237__7_ ( .D(n18728), .CP(wclk), .Q(ram[14487]) );
  DFF ram_reg_237__6_ ( .D(n18727), .CP(wclk), .Q(ram[14486]) );
  DFF ram_reg_237__5_ ( .D(n18726), .CP(wclk), .Q(ram[14485]) );
  DFF ram_reg_237__4_ ( .D(n18725), .CP(wclk), .Q(ram[14484]) );
  DFF ram_reg_237__3_ ( .D(n18724), .CP(wclk), .Q(ram[14483]) );
  DFF ram_reg_237__2_ ( .D(n18723), .CP(wclk), .Q(ram[14482]) );
  DFF ram_reg_237__1_ ( .D(n18722), .CP(wclk), .Q(ram[14481]) );
  DFF ram_reg_237__0_ ( .D(n18721), .CP(wclk), .Q(ram[14480]) );
  DFF ram_reg_241__7_ ( .D(n18696), .CP(wclk), .Q(ram[14455]) );
  DFF ram_reg_241__6_ ( .D(n18695), .CP(wclk), .Q(ram[14454]) );
  DFF ram_reg_241__5_ ( .D(n18694), .CP(wclk), .Q(ram[14453]) );
  DFF ram_reg_241__4_ ( .D(n18693), .CP(wclk), .Q(ram[14452]) );
  DFF ram_reg_241__3_ ( .D(n18692), .CP(wclk), .Q(ram[14451]) );
  DFF ram_reg_241__2_ ( .D(n18691), .CP(wclk), .Q(ram[14450]) );
  DFF ram_reg_241__1_ ( .D(n18690), .CP(wclk), .Q(ram[14449]) );
  DFF ram_reg_241__0_ ( .D(n18689), .CP(wclk), .Q(ram[14448]) );
  DFF ram_reg_249__7_ ( .D(n18632), .CP(wclk), .Q(ram[14391]) );
  DFF ram_reg_249__6_ ( .D(n18631), .CP(wclk), .Q(ram[14390]) );
  DFF ram_reg_249__5_ ( .D(n18630), .CP(wclk), .Q(ram[14389]) );
  DFF ram_reg_249__4_ ( .D(n18629), .CP(wclk), .Q(ram[14388]) );
  DFF ram_reg_249__3_ ( .D(n18628), .CP(wclk), .Q(ram[14387]) );
  DFF ram_reg_249__2_ ( .D(n18627), .CP(wclk), .Q(ram[14386]) );
  DFF ram_reg_249__1_ ( .D(n18626), .CP(wclk), .Q(ram[14385]) );
  DFF ram_reg_249__0_ ( .D(n18625), .CP(wclk), .Q(ram[14384]) );
  DFF ram_reg_253__7_ ( .D(n18600), .CP(wclk), .Q(ram[14359]) );
  DFF ram_reg_253__6_ ( .D(n18599), .CP(wclk), .Q(ram[14358]) );
  DFF ram_reg_253__5_ ( .D(n18598), .CP(wclk), .Q(ram[14357]) );
  DFF ram_reg_253__4_ ( .D(n18597), .CP(wclk), .Q(ram[14356]) );
  DFF ram_reg_253__3_ ( .D(n18596), .CP(wclk), .Q(ram[14355]) );
  DFF ram_reg_253__2_ ( .D(n18595), .CP(wclk), .Q(ram[14354]) );
  DFF ram_reg_253__1_ ( .D(n18594), .CP(wclk), .Q(ram[14353]) );
  DFF ram_reg_253__0_ ( .D(n18593), .CP(wclk), .Q(ram[14352]) );
  DFF ram_reg_265__7_ ( .D(n18504), .CP(wclk), .Q(ram[14263]) );
  DFF ram_reg_265__6_ ( .D(n18503), .CP(wclk), .Q(ram[14262]) );
  DFF ram_reg_265__5_ ( .D(n18502), .CP(wclk), .Q(ram[14261]) );
  DFF ram_reg_265__4_ ( .D(n18501), .CP(wclk), .Q(ram[14260]) );
  DFF ram_reg_265__3_ ( .D(n18500), .CP(wclk), .Q(ram[14259]) );
  DFF ram_reg_265__2_ ( .D(n18499), .CP(wclk), .Q(ram[14258]) );
  DFF ram_reg_265__1_ ( .D(n18498), .CP(wclk), .Q(ram[14257]) );
  DFF ram_reg_265__0_ ( .D(n18497), .CP(wclk), .Q(ram[14256]) );
  DFF ram_reg_297__7_ ( .D(n18248), .CP(wclk), .Q(ram[14007]) );
  DFF ram_reg_297__6_ ( .D(n18247), .CP(wclk), .Q(ram[14006]) );
  DFF ram_reg_297__5_ ( .D(n18246), .CP(wclk), .Q(ram[14005]) );
  DFF ram_reg_297__4_ ( .D(n18245), .CP(wclk), .Q(ram[14004]) );
  DFF ram_reg_297__3_ ( .D(n18244), .CP(wclk), .Q(ram[14003]) );
  DFF ram_reg_297__2_ ( .D(n18243), .CP(wclk), .Q(ram[14002]) );
  DFF ram_reg_297__1_ ( .D(n18242), .CP(wclk), .Q(ram[14001]) );
  DFF ram_reg_297__0_ ( .D(n18241), .CP(wclk), .Q(ram[14000]) );
  DFF ram_reg_301__7_ ( .D(n18216), .CP(wclk), .Q(ram[13975]) );
  DFF ram_reg_301__6_ ( .D(n18215), .CP(wclk), .Q(ram[13974]) );
  DFF ram_reg_301__5_ ( .D(n18214), .CP(wclk), .Q(ram[13973]) );
  DFF ram_reg_301__4_ ( .D(n18213), .CP(wclk), .Q(ram[13972]) );
  DFF ram_reg_301__3_ ( .D(n18212), .CP(wclk), .Q(ram[13971]) );
  DFF ram_reg_301__2_ ( .D(n18211), .CP(wclk), .Q(ram[13970]) );
  DFF ram_reg_301__1_ ( .D(n18210), .CP(wclk), .Q(ram[13969]) );
  DFF ram_reg_301__0_ ( .D(n18209), .CP(wclk), .Q(ram[13968]) );
  DFF ram_reg_313__7_ ( .D(n18120), .CP(wclk), .Q(ram[13879]) );
  DFF ram_reg_313__6_ ( .D(n18119), .CP(wclk), .Q(ram[13878]) );
  DFF ram_reg_313__5_ ( .D(n18118), .CP(wclk), .Q(ram[13877]) );
  DFF ram_reg_313__4_ ( .D(n18117), .CP(wclk), .Q(ram[13876]) );
  DFF ram_reg_313__3_ ( .D(n18116), .CP(wclk), .Q(ram[13875]) );
  DFF ram_reg_313__2_ ( .D(n18115), .CP(wclk), .Q(ram[13874]) );
  DFF ram_reg_313__1_ ( .D(n18114), .CP(wclk), .Q(ram[13873]) );
  DFF ram_reg_313__0_ ( .D(n18113), .CP(wclk), .Q(ram[13872]) );
  DFF ram_reg_317__7_ ( .D(n18088), .CP(wclk), .Q(ram[13847]) );
  DFF ram_reg_317__6_ ( .D(n18087), .CP(wclk), .Q(ram[13846]) );
  DFF ram_reg_317__5_ ( .D(n18086), .CP(wclk), .Q(ram[13845]) );
  DFF ram_reg_317__4_ ( .D(n18085), .CP(wclk), .Q(ram[13844]) );
  DFF ram_reg_317__3_ ( .D(n18084), .CP(wclk), .Q(ram[13843]) );
  DFF ram_reg_317__2_ ( .D(n18083), .CP(wclk), .Q(ram[13842]) );
  DFF ram_reg_317__1_ ( .D(n18082), .CP(wclk), .Q(ram[13841]) );
  DFF ram_reg_317__0_ ( .D(n18081), .CP(wclk), .Q(ram[13840]) );
  DFF ram_reg_377__7_ ( .D(n17608), .CP(wclk), .Q(ram[13367]) );
  DFF ram_reg_377__6_ ( .D(n17607), .CP(wclk), .Q(ram[13366]) );
  DFF ram_reg_377__5_ ( .D(n17606), .CP(wclk), .Q(ram[13365]) );
  DFF ram_reg_377__4_ ( .D(n17605), .CP(wclk), .Q(ram[13364]) );
  DFF ram_reg_377__3_ ( .D(n17604), .CP(wclk), .Q(ram[13363]) );
  DFF ram_reg_377__2_ ( .D(n17603), .CP(wclk), .Q(ram[13362]) );
  DFF ram_reg_377__1_ ( .D(n17602), .CP(wclk), .Q(ram[13361]) );
  DFF ram_reg_377__0_ ( .D(n17601), .CP(wclk), .Q(ram[13360]) );
  DFF ram_reg_385__7_ ( .D(n17544), .CP(wclk), .Q(ram[13303]) );
  DFF ram_reg_385__6_ ( .D(n17543), .CP(wclk), .Q(ram[13302]) );
  DFF ram_reg_385__5_ ( .D(n17542), .CP(wclk), .Q(ram[13301]) );
  DFF ram_reg_385__4_ ( .D(n17541), .CP(wclk), .Q(ram[13300]) );
  DFF ram_reg_385__3_ ( .D(n17540), .CP(wclk), .Q(ram[13299]) );
  DFF ram_reg_385__2_ ( .D(n17539), .CP(wclk), .Q(ram[13298]) );
  DFF ram_reg_385__1_ ( .D(n17538), .CP(wclk), .Q(ram[13297]) );
  DFF ram_reg_385__0_ ( .D(n17537), .CP(wclk), .Q(ram[13296]) );
  DFF ram_reg_393__7_ ( .D(n17480), .CP(wclk), .Q(ram[13239]) );
  DFF ram_reg_393__6_ ( .D(n17479), .CP(wclk), .Q(ram[13238]) );
  DFF ram_reg_393__5_ ( .D(n17478), .CP(wclk), .Q(ram[13237]) );
  DFF ram_reg_393__4_ ( .D(n17477), .CP(wclk), .Q(ram[13236]) );
  DFF ram_reg_393__3_ ( .D(n17476), .CP(wclk), .Q(ram[13235]) );
  DFF ram_reg_393__2_ ( .D(n17475), .CP(wclk), .Q(ram[13234]) );
  DFF ram_reg_393__1_ ( .D(n17474), .CP(wclk), .Q(ram[13233]) );
  DFF ram_reg_393__0_ ( .D(n17473), .CP(wclk), .Q(ram[13232]) );
  DFF ram_reg_397__7_ ( .D(n17448), .CP(wclk), .Q(ram[13207]) );
  DFF ram_reg_397__6_ ( .D(n17447), .CP(wclk), .Q(ram[13206]) );
  DFF ram_reg_397__5_ ( .D(n17446), .CP(wclk), .Q(ram[13205]) );
  DFF ram_reg_397__4_ ( .D(n17445), .CP(wclk), .Q(ram[13204]) );
  DFF ram_reg_397__3_ ( .D(n17444), .CP(wclk), .Q(ram[13203]) );
  DFF ram_reg_397__2_ ( .D(n17443), .CP(wclk), .Q(ram[13202]) );
  DFF ram_reg_397__1_ ( .D(n17442), .CP(wclk), .Q(ram[13201]) );
  DFF ram_reg_397__0_ ( .D(n17441), .CP(wclk), .Q(ram[13200]) );
  DFF ram_reg_409__7_ ( .D(n17352), .CP(wclk), .Q(ram[13111]) );
  DFF ram_reg_409__6_ ( .D(n17351), .CP(wclk), .Q(ram[13110]) );
  DFF ram_reg_409__5_ ( .D(n17350), .CP(wclk), .Q(ram[13109]) );
  DFF ram_reg_409__4_ ( .D(n17349), .CP(wclk), .Q(ram[13108]) );
  DFF ram_reg_409__3_ ( .D(n17348), .CP(wclk), .Q(ram[13107]) );
  DFF ram_reg_409__2_ ( .D(n17347), .CP(wclk), .Q(ram[13106]) );
  DFF ram_reg_409__1_ ( .D(n17346), .CP(wclk), .Q(ram[13105]) );
  DFF ram_reg_409__0_ ( .D(n17345), .CP(wclk), .Q(ram[13104]) );
  DFF ram_reg_413__7_ ( .D(n17320), .CP(wclk), .Q(ram[13079]) );
  DFF ram_reg_413__6_ ( .D(n17319), .CP(wclk), .Q(ram[13078]) );
  DFF ram_reg_413__5_ ( .D(n17318), .CP(wclk), .Q(ram[13077]) );
  DFF ram_reg_413__4_ ( .D(n17317), .CP(wclk), .Q(ram[13076]) );
  DFF ram_reg_413__3_ ( .D(n17316), .CP(wclk), .Q(ram[13075]) );
  DFF ram_reg_413__2_ ( .D(n17315), .CP(wclk), .Q(ram[13074]) );
  DFF ram_reg_413__1_ ( .D(n17314), .CP(wclk), .Q(ram[13073]) );
  DFF ram_reg_413__0_ ( .D(n17313), .CP(wclk), .Q(ram[13072]) );
  DFF ram_reg_417__7_ ( .D(n17288), .CP(wclk), .Q(ram[13047]) );
  DFF ram_reg_417__6_ ( .D(n17287), .CP(wclk), .Q(ram[13046]) );
  DFF ram_reg_417__5_ ( .D(n17286), .CP(wclk), .Q(ram[13045]) );
  DFF ram_reg_417__4_ ( .D(n17285), .CP(wclk), .Q(ram[13044]) );
  DFF ram_reg_417__3_ ( .D(n17284), .CP(wclk), .Q(ram[13043]) );
  DFF ram_reg_417__2_ ( .D(n17283), .CP(wclk), .Q(ram[13042]) );
  DFF ram_reg_417__1_ ( .D(n17282), .CP(wclk), .Q(ram[13041]) );
  DFF ram_reg_417__0_ ( .D(n17281), .CP(wclk), .Q(ram[13040]) );
  DFF ram_reg_425__7_ ( .D(n17224), .CP(wclk), .Q(ram[12983]) );
  DFF ram_reg_425__6_ ( .D(n17223), .CP(wclk), .Q(ram[12982]) );
  DFF ram_reg_425__5_ ( .D(n17222), .CP(wclk), .Q(ram[12981]) );
  DFF ram_reg_425__4_ ( .D(n17221), .CP(wclk), .Q(ram[12980]) );
  DFF ram_reg_425__3_ ( .D(n17220), .CP(wclk), .Q(ram[12979]) );
  DFF ram_reg_425__2_ ( .D(n17219), .CP(wclk), .Q(ram[12978]) );
  DFF ram_reg_425__1_ ( .D(n17218), .CP(wclk), .Q(ram[12977]) );
  DFF ram_reg_425__0_ ( .D(n17217), .CP(wclk), .Q(ram[12976]) );
  DFF ram_reg_429__7_ ( .D(n17192), .CP(wclk), .Q(ram[12951]) );
  DFF ram_reg_429__6_ ( .D(n17191), .CP(wclk), .Q(ram[12950]) );
  DFF ram_reg_429__5_ ( .D(n17190), .CP(wclk), .Q(ram[12949]) );
  DFF ram_reg_429__4_ ( .D(n17189), .CP(wclk), .Q(ram[12948]) );
  DFF ram_reg_429__3_ ( .D(n17188), .CP(wclk), .Q(ram[12947]) );
  DFF ram_reg_429__2_ ( .D(n17187), .CP(wclk), .Q(ram[12946]) );
  DFF ram_reg_429__1_ ( .D(n17186), .CP(wclk), .Q(ram[12945]) );
  DFF ram_reg_429__0_ ( .D(n17185), .CP(wclk), .Q(ram[12944]) );
  DFF ram_reg_433__7_ ( .D(n17160), .CP(wclk), .Q(ram[12919]) );
  DFF ram_reg_433__6_ ( .D(n17159), .CP(wclk), .Q(ram[12918]) );
  DFF ram_reg_433__5_ ( .D(n17158), .CP(wclk), .Q(ram[12917]) );
  DFF ram_reg_433__4_ ( .D(n17157), .CP(wclk), .Q(ram[12916]) );
  DFF ram_reg_433__3_ ( .D(n17156), .CP(wclk), .Q(ram[12915]) );
  DFF ram_reg_433__2_ ( .D(n17155), .CP(wclk), .Q(ram[12914]) );
  DFF ram_reg_433__1_ ( .D(n17154), .CP(wclk), .Q(ram[12913]) );
  DFF ram_reg_433__0_ ( .D(n17153), .CP(wclk), .Q(ram[12912]) );
  DFF ram_reg_437__7_ ( .D(n17128), .CP(wclk), .Q(ram[12887]) );
  DFF ram_reg_437__6_ ( .D(n17127), .CP(wclk), .Q(ram[12886]) );
  DFF ram_reg_437__5_ ( .D(n17126), .CP(wclk), .Q(ram[12885]) );
  DFF ram_reg_437__4_ ( .D(n17125), .CP(wclk), .Q(ram[12884]) );
  DFF ram_reg_437__3_ ( .D(n17124), .CP(wclk), .Q(ram[12883]) );
  DFF ram_reg_437__2_ ( .D(n17123), .CP(wclk), .Q(ram[12882]) );
  DFF ram_reg_437__1_ ( .D(n17122), .CP(wclk), .Q(ram[12881]) );
  DFF ram_reg_437__0_ ( .D(n17121), .CP(wclk), .Q(ram[12880]) );
  DFF ram_reg_441__7_ ( .D(n17096), .CP(wclk), .Q(ram[12855]) );
  DFF ram_reg_441__6_ ( .D(n17095), .CP(wclk), .Q(ram[12854]) );
  DFF ram_reg_441__5_ ( .D(n17094), .CP(wclk), .Q(ram[12853]) );
  DFF ram_reg_441__4_ ( .D(n17093), .CP(wclk), .Q(ram[12852]) );
  DFF ram_reg_441__3_ ( .D(n17092), .CP(wclk), .Q(ram[12851]) );
  DFF ram_reg_441__2_ ( .D(n17091), .CP(wclk), .Q(ram[12850]) );
  DFF ram_reg_441__1_ ( .D(n17090), .CP(wclk), .Q(ram[12849]) );
  DFF ram_reg_441__0_ ( .D(n17089), .CP(wclk), .Q(ram[12848]) );
  DFF ram_reg_445__7_ ( .D(n17064), .CP(wclk), .Q(ram[12823]) );
  DFF ram_reg_445__6_ ( .D(n17063), .CP(wclk), .Q(ram[12822]) );
  DFF ram_reg_445__5_ ( .D(n17062), .CP(wclk), .Q(ram[12821]) );
  DFF ram_reg_445__4_ ( .D(n17061), .CP(wclk), .Q(ram[12820]) );
  DFF ram_reg_445__3_ ( .D(n17060), .CP(wclk), .Q(ram[12819]) );
  DFF ram_reg_445__2_ ( .D(n17059), .CP(wclk), .Q(ram[12818]) );
  DFF ram_reg_445__1_ ( .D(n17058), .CP(wclk), .Q(ram[12817]) );
  DFF ram_reg_445__0_ ( .D(n17057), .CP(wclk), .Q(ram[12816]) );
  DFF ram_reg_457__7_ ( .D(n16968), .CP(wclk), .Q(ram[12727]) );
  DFF ram_reg_457__6_ ( .D(n16967), .CP(wclk), .Q(ram[12726]) );
  DFF ram_reg_457__5_ ( .D(n16966), .CP(wclk), .Q(ram[12725]) );
  DFF ram_reg_457__4_ ( .D(n16965), .CP(wclk), .Q(ram[12724]) );
  DFF ram_reg_457__3_ ( .D(n16964), .CP(wclk), .Q(ram[12723]) );
  DFF ram_reg_457__2_ ( .D(n16963), .CP(wclk), .Q(ram[12722]) );
  DFF ram_reg_457__1_ ( .D(n16962), .CP(wclk), .Q(ram[12721]) );
  DFF ram_reg_457__0_ ( .D(n16961), .CP(wclk), .Q(ram[12720]) );
  DFF ram_reg_461__7_ ( .D(n16936), .CP(wclk), .Q(ram[12695]) );
  DFF ram_reg_461__6_ ( .D(n16935), .CP(wclk), .Q(ram[12694]) );
  DFF ram_reg_461__5_ ( .D(n16934), .CP(wclk), .Q(ram[12693]) );
  DFF ram_reg_461__4_ ( .D(n16933), .CP(wclk), .Q(ram[12692]) );
  DFF ram_reg_461__3_ ( .D(n16932), .CP(wclk), .Q(ram[12691]) );
  DFF ram_reg_461__2_ ( .D(n16931), .CP(wclk), .Q(ram[12690]) );
  DFF ram_reg_461__1_ ( .D(n16930), .CP(wclk), .Q(ram[12689]) );
  DFF ram_reg_461__0_ ( .D(n16929), .CP(wclk), .Q(ram[12688]) );
  DFF ram_reg_473__7_ ( .D(n16840), .CP(wclk), .Q(ram[12599]) );
  DFF ram_reg_473__6_ ( .D(n16839), .CP(wclk), .Q(ram[12598]) );
  DFF ram_reg_473__5_ ( .D(n16838), .CP(wclk), .Q(ram[12597]) );
  DFF ram_reg_473__4_ ( .D(n16837), .CP(wclk), .Q(ram[12596]) );
  DFF ram_reg_473__3_ ( .D(n16836), .CP(wclk), .Q(ram[12595]) );
  DFF ram_reg_473__2_ ( .D(n16835), .CP(wclk), .Q(ram[12594]) );
  DFF ram_reg_473__1_ ( .D(n16834), .CP(wclk), .Q(ram[12593]) );
  DFF ram_reg_473__0_ ( .D(n16833), .CP(wclk), .Q(ram[12592]) );
  DFF ram_reg_477__7_ ( .D(n16808), .CP(wclk), .Q(ram[12567]) );
  DFF ram_reg_477__6_ ( .D(n16807), .CP(wclk), .Q(ram[12566]) );
  DFF ram_reg_477__5_ ( .D(n16806), .CP(wclk), .Q(ram[12565]) );
  DFF ram_reg_477__4_ ( .D(n16805), .CP(wclk), .Q(ram[12564]) );
  DFF ram_reg_477__3_ ( .D(n16804), .CP(wclk), .Q(ram[12563]) );
  DFF ram_reg_477__2_ ( .D(n16803), .CP(wclk), .Q(ram[12562]) );
  DFF ram_reg_477__1_ ( .D(n16802), .CP(wclk), .Q(ram[12561]) );
  DFF ram_reg_477__0_ ( .D(n16801), .CP(wclk), .Q(ram[12560]) );
  DFF ram_reg_481__7_ ( .D(n16776), .CP(wclk), .Q(ram[12535]) );
  DFF ram_reg_481__6_ ( .D(n16775), .CP(wclk), .Q(ram[12534]) );
  DFF ram_reg_481__5_ ( .D(n16774), .CP(wclk), .Q(ram[12533]) );
  DFF ram_reg_481__4_ ( .D(n16773), .CP(wclk), .Q(ram[12532]) );
  DFF ram_reg_481__3_ ( .D(n16772), .CP(wclk), .Q(ram[12531]) );
  DFF ram_reg_481__2_ ( .D(n16771), .CP(wclk), .Q(ram[12530]) );
  DFF ram_reg_481__1_ ( .D(n16770), .CP(wclk), .Q(ram[12529]) );
  DFF ram_reg_481__0_ ( .D(n16769), .CP(wclk), .Q(ram[12528]) );
  DFF ram_reg_489__7_ ( .D(n16712), .CP(wclk), .Q(ram[12471]) );
  DFF ram_reg_489__6_ ( .D(n16711), .CP(wclk), .Q(ram[12470]) );
  DFF ram_reg_489__5_ ( .D(n16710), .CP(wclk), .Q(ram[12469]) );
  DFF ram_reg_489__4_ ( .D(n16709), .CP(wclk), .Q(ram[12468]) );
  DFF ram_reg_489__3_ ( .D(n16708), .CP(wclk), .Q(ram[12467]) );
  DFF ram_reg_489__2_ ( .D(n16707), .CP(wclk), .Q(ram[12466]) );
  DFF ram_reg_489__1_ ( .D(n16706), .CP(wclk), .Q(ram[12465]) );
  DFF ram_reg_489__0_ ( .D(n16705), .CP(wclk), .Q(ram[12464]) );
  DFF ram_reg_493__7_ ( .D(n16680), .CP(wclk), .Q(ram[12439]) );
  DFF ram_reg_493__6_ ( .D(n16679), .CP(wclk), .Q(ram[12438]) );
  DFF ram_reg_493__5_ ( .D(n16678), .CP(wclk), .Q(ram[12437]) );
  DFF ram_reg_493__4_ ( .D(n16677), .CP(wclk), .Q(ram[12436]) );
  DFF ram_reg_493__3_ ( .D(n16676), .CP(wclk), .Q(ram[12435]) );
  DFF ram_reg_493__2_ ( .D(n16675), .CP(wclk), .Q(ram[12434]) );
  DFF ram_reg_493__1_ ( .D(n16674), .CP(wclk), .Q(ram[12433]) );
  DFF ram_reg_493__0_ ( .D(n16673), .CP(wclk), .Q(ram[12432]) );
  DFF ram_reg_497__7_ ( .D(n16648), .CP(wclk), .Q(ram[12407]) );
  DFF ram_reg_497__6_ ( .D(n16647), .CP(wclk), .Q(ram[12406]) );
  DFF ram_reg_497__5_ ( .D(n16646), .CP(wclk), .Q(ram[12405]) );
  DFF ram_reg_497__4_ ( .D(n16645), .CP(wclk), .Q(ram[12404]) );
  DFF ram_reg_497__3_ ( .D(n16644), .CP(wclk), .Q(ram[12403]) );
  DFF ram_reg_497__2_ ( .D(n16643), .CP(wclk), .Q(ram[12402]) );
  DFF ram_reg_497__1_ ( .D(n16642), .CP(wclk), .Q(ram[12401]) );
  DFF ram_reg_497__0_ ( .D(n16641), .CP(wclk), .Q(ram[12400]) );
  DFF ram_reg_505__7_ ( .D(n16584), .CP(wclk), .Q(ram[12343]) );
  DFF ram_reg_505__6_ ( .D(n16583), .CP(wclk), .Q(ram[12342]) );
  DFF ram_reg_505__5_ ( .D(n16582), .CP(wclk), .Q(ram[12341]) );
  DFF ram_reg_505__4_ ( .D(n16581), .CP(wclk), .Q(ram[12340]) );
  DFF ram_reg_505__3_ ( .D(n16580), .CP(wclk), .Q(ram[12339]) );
  DFF ram_reg_505__2_ ( .D(n16579), .CP(wclk), .Q(ram[12338]) );
  DFF ram_reg_505__1_ ( .D(n16578), .CP(wclk), .Q(ram[12337]) );
  DFF ram_reg_505__0_ ( .D(n16577), .CP(wclk), .Q(ram[12336]) );
  DFF ram_reg_509__7_ ( .D(n16552), .CP(wclk), .Q(ram[12311]) );
  DFF ram_reg_509__6_ ( .D(n16551), .CP(wclk), .Q(ram[12310]) );
  DFF ram_reg_509__5_ ( .D(n16550), .CP(wclk), .Q(ram[12309]) );
  DFF ram_reg_509__4_ ( .D(n16549), .CP(wclk), .Q(ram[12308]) );
  DFF ram_reg_509__3_ ( .D(n16548), .CP(wclk), .Q(ram[12307]) );
  DFF ram_reg_509__2_ ( .D(n16547), .CP(wclk), .Q(ram[12306]) );
  DFF ram_reg_509__1_ ( .D(n16546), .CP(wclk), .Q(ram[12305]) );
  DFF ram_reg_509__0_ ( .D(n16545), .CP(wclk), .Q(ram[12304]) );
  DFF ram_reg_521__7_ ( .D(n16456), .CP(wclk), .Q(ram[12215]) );
  DFF ram_reg_521__6_ ( .D(n16455), .CP(wclk), .Q(ram[12214]) );
  DFF ram_reg_521__5_ ( .D(n16454), .CP(wclk), .Q(ram[12213]) );
  DFF ram_reg_521__4_ ( .D(n16453), .CP(wclk), .Q(ram[12212]) );
  DFF ram_reg_521__3_ ( .D(n16452), .CP(wclk), .Q(ram[12211]) );
  DFF ram_reg_521__2_ ( .D(n16451), .CP(wclk), .Q(ram[12210]) );
  DFF ram_reg_521__1_ ( .D(n16450), .CP(wclk), .Q(ram[12209]) );
  DFF ram_reg_521__0_ ( .D(n16449), .CP(wclk), .Q(ram[12208]) );
  DFF ram_reg_525__7_ ( .D(n16424), .CP(wclk), .Q(ram[12183]) );
  DFF ram_reg_525__6_ ( .D(n16423), .CP(wclk), .Q(ram[12182]) );
  DFF ram_reg_525__5_ ( .D(n16422), .CP(wclk), .Q(ram[12181]) );
  DFF ram_reg_525__4_ ( .D(n16421), .CP(wclk), .Q(ram[12180]) );
  DFF ram_reg_525__3_ ( .D(n16420), .CP(wclk), .Q(ram[12179]) );
  DFF ram_reg_525__2_ ( .D(n16419), .CP(wclk), .Q(ram[12178]) );
  DFF ram_reg_525__1_ ( .D(n16418), .CP(wclk), .Q(ram[12177]) );
  DFF ram_reg_525__0_ ( .D(n16417), .CP(wclk), .Q(ram[12176]) );
  DFF ram_reg_537__7_ ( .D(n16328), .CP(wclk), .Q(ram[12087]) );
  DFF ram_reg_537__6_ ( .D(n16327), .CP(wclk), .Q(ram[12086]) );
  DFF ram_reg_537__5_ ( .D(n16326), .CP(wclk), .Q(ram[12085]) );
  DFF ram_reg_537__4_ ( .D(n16325), .CP(wclk), .Q(ram[12084]) );
  DFF ram_reg_537__3_ ( .D(n16324), .CP(wclk), .Q(ram[12083]) );
  DFF ram_reg_537__2_ ( .D(n16323), .CP(wclk), .Q(ram[12082]) );
  DFF ram_reg_537__1_ ( .D(n16322), .CP(wclk), .Q(ram[12081]) );
  DFF ram_reg_537__0_ ( .D(n16321), .CP(wclk), .Q(ram[12080]) );
  DFF ram_reg_541__7_ ( .D(n16296), .CP(wclk), .Q(ram[12055]) );
  DFF ram_reg_541__6_ ( .D(n16295), .CP(wclk), .Q(ram[12054]) );
  DFF ram_reg_541__5_ ( .D(n16294), .CP(wclk), .Q(ram[12053]) );
  DFF ram_reg_541__4_ ( .D(n16293), .CP(wclk), .Q(ram[12052]) );
  DFF ram_reg_541__3_ ( .D(n16292), .CP(wclk), .Q(ram[12051]) );
  DFF ram_reg_541__2_ ( .D(n16291), .CP(wclk), .Q(ram[12050]) );
  DFF ram_reg_541__1_ ( .D(n16290), .CP(wclk), .Q(ram[12049]) );
  DFF ram_reg_541__0_ ( .D(n16289), .CP(wclk), .Q(ram[12048]) );
  DFF ram_reg_545__7_ ( .D(n16264), .CP(wclk), .Q(ram[12023]) );
  DFF ram_reg_545__6_ ( .D(n16263), .CP(wclk), .Q(ram[12022]) );
  DFF ram_reg_545__5_ ( .D(n16262), .CP(wclk), .Q(ram[12021]) );
  DFF ram_reg_545__4_ ( .D(n16261), .CP(wclk), .Q(ram[12020]) );
  DFF ram_reg_545__3_ ( .D(n16260), .CP(wclk), .Q(ram[12019]) );
  DFF ram_reg_545__2_ ( .D(n16259), .CP(wclk), .Q(ram[12018]) );
  DFF ram_reg_545__1_ ( .D(n16258), .CP(wclk), .Q(ram[12017]) );
  DFF ram_reg_545__0_ ( .D(n16257), .CP(wclk), .Q(ram[12016]) );
  DFF ram_reg_553__7_ ( .D(n16200), .CP(wclk), .Q(ram[11959]) );
  DFF ram_reg_553__6_ ( .D(n16199), .CP(wclk), .Q(ram[11958]) );
  DFF ram_reg_553__5_ ( .D(n16198), .CP(wclk), .Q(ram[11957]) );
  DFF ram_reg_553__4_ ( .D(n16197), .CP(wclk), .Q(ram[11956]) );
  DFF ram_reg_553__3_ ( .D(n16196), .CP(wclk), .Q(ram[11955]) );
  DFF ram_reg_553__2_ ( .D(n16195), .CP(wclk), .Q(ram[11954]) );
  DFF ram_reg_553__1_ ( .D(n16194), .CP(wclk), .Q(ram[11953]) );
  DFF ram_reg_553__0_ ( .D(n16193), .CP(wclk), .Q(ram[11952]) );
  DFF ram_reg_557__7_ ( .D(n16168), .CP(wclk), .Q(ram[11927]) );
  DFF ram_reg_557__6_ ( .D(n16167), .CP(wclk), .Q(ram[11926]) );
  DFF ram_reg_557__5_ ( .D(n16166), .CP(wclk), .Q(ram[11925]) );
  DFF ram_reg_557__4_ ( .D(n16165), .CP(wclk), .Q(ram[11924]) );
  DFF ram_reg_557__3_ ( .D(n16164), .CP(wclk), .Q(ram[11923]) );
  DFF ram_reg_557__2_ ( .D(n16163), .CP(wclk), .Q(ram[11922]) );
  DFF ram_reg_557__1_ ( .D(n16162), .CP(wclk), .Q(ram[11921]) );
  DFF ram_reg_557__0_ ( .D(n16161), .CP(wclk), .Q(ram[11920]) );
  DFF ram_reg_561__7_ ( .D(n16136), .CP(wclk), .Q(ram[11895]) );
  DFF ram_reg_561__6_ ( .D(n16135), .CP(wclk), .Q(ram[11894]) );
  DFF ram_reg_561__5_ ( .D(n16134), .CP(wclk), .Q(ram[11893]) );
  DFF ram_reg_561__4_ ( .D(n16133), .CP(wclk), .Q(ram[11892]) );
  DFF ram_reg_561__3_ ( .D(n16132), .CP(wclk), .Q(ram[11891]) );
  DFF ram_reg_561__2_ ( .D(n16131), .CP(wclk), .Q(ram[11890]) );
  DFF ram_reg_561__1_ ( .D(n16130), .CP(wclk), .Q(ram[11889]) );
  DFF ram_reg_561__0_ ( .D(n16129), .CP(wclk), .Q(ram[11888]) );
  DFF ram_reg_569__7_ ( .D(n16072), .CP(wclk), .Q(ram[11831]) );
  DFF ram_reg_569__6_ ( .D(n16071), .CP(wclk), .Q(ram[11830]) );
  DFF ram_reg_569__5_ ( .D(n16070), .CP(wclk), .Q(ram[11829]) );
  DFF ram_reg_569__4_ ( .D(n16069), .CP(wclk), .Q(ram[11828]) );
  DFF ram_reg_569__3_ ( .D(n16068), .CP(wclk), .Q(ram[11827]) );
  DFF ram_reg_569__2_ ( .D(n16067), .CP(wclk), .Q(ram[11826]) );
  DFF ram_reg_569__1_ ( .D(n16066), .CP(wclk), .Q(ram[11825]) );
  DFF ram_reg_569__0_ ( .D(n16065), .CP(wclk), .Q(ram[11824]) );
  DFF ram_reg_573__7_ ( .D(n16040), .CP(wclk), .Q(ram[11799]) );
  DFF ram_reg_573__6_ ( .D(n16039), .CP(wclk), .Q(ram[11798]) );
  DFF ram_reg_573__5_ ( .D(n16038), .CP(wclk), .Q(ram[11797]) );
  DFF ram_reg_573__4_ ( .D(n16037), .CP(wclk), .Q(ram[11796]) );
  DFF ram_reg_573__3_ ( .D(n16036), .CP(wclk), .Q(ram[11795]) );
  DFF ram_reg_573__2_ ( .D(n16035), .CP(wclk), .Q(ram[11794]) );
  DFF ram_reg_573__1_ ( .D(n16034), .CP(wclk), .Q(ram[11793]) );
  DFF ram_reg_573__0_ ( .D(n16033), .CP(wclk), .Q(ram[11792]) );
  DFF ram_reg_585__7_ ( .D(n15944), .CP(wclk), .Q(ram[11703]) );
  DFF ram_reg_585__6_ ( .D(n15943), .CP(wclk), .Q(ram[11702]) );
  DFF ram_reg_585__5_ ( .D(n15942), .CP(wclk), .Q(ram[11701]) );
  DFF ram_reg_585__4_ ( .D(n15941), .CP(wclk), .Q(ram[11700]) );
  DFF ram_reg_585__3_ ( .D(n15940), .CP(wclk), .Q(ram[11699]) );
  DFF ram_reg_585__2_ ( .D(n15939), .CP(wclk), .Q(ram[11698]) );
  DFF ram_reg_585__1_ ( .D(n15938), .CP(wclk), .Q(ram[11697]) );
  DFF ram_reg_585__0_ ( .D(n15937), .CP(wclk), .Q(ram[11696]) );
  DFF ram_reg_617__7_ ( .D(n15688), .CP(wclk), .Q(ram[11447]) );
  DFF ram_reg_617__6_ ( .D(n15687), .CP(wclk), .Q(ram[11446]) );
  DFF ram_reg_617__5_ ( .D(n15686), .CP(wclk), .Q(ram[11445]) );
  DFF ram_reg_617__4_ ( .D(n15685), .CP(wclk), .Q(ram[11444]) );
  DFF ram_reg_617__3_ ( .D(n15684), .CP(wclk), .Q(ram[11443]) );
  DFF ram_reg_617__2_ ( .D(n15683), .CP(wclk), .Q(ram[11442]) );
  DFF ram_reg_617__1_ ( .D(n15682), .CP(wclk), .Q(ram[11441]) );
  DFF ram_reg_617__0_ ( .D(n15681), .CP(wclk), .Q(ram[11440]) );
  DFF ram_reg_621__7_ ( .D(n15656), .CP(wclk), .Q(ram[11415]) );
  DFF ram_reg_621__6_ ( .D(n15655), .CP(wclk), .Q(ram[11414]) );
  DFF ram_reg_621__5_ ( .D(n15654), .CP(wclk), .Q(ram[11413]) );
  DFF ram_reg_621__4_ ( .D(n15653), .CP(wclk), .Q(ram[11412]) );
  DFF ram_reg_621__3_ ( .D(n15652), .CP(wclk), .Q(ram[11411]) );
  DFF ram_reg_621__2_ ( .D(n15651), .CP(wclk), .Q(ram[11410]) );
  DFF ram_reg_621__1_ ( .D(n15650), .CP(wclk), .Q(ram[11409]) );
  DFF ram_reg_621__0_ ( .D(n15649), .CP(wclk), .Q(ram[11408]) );
  DFF ram_reg_633__7_ ( .D(n15560), .CP(wclk), .Q(ram[11319]) );
  DFF ram_reg_633__6_ ( .D(n15559), .CP(wclk), .Q(ram[11318]) );
  DFF ram_reg_633__5_ ( .D(n15558), .CP(wclk), .Q(ram[11317]) );
  DFF ram_reg_633__4_ ( .D(n15557), .CP(wclk), .Q(ram[11316]) );
  DFF ram_reg_633__3_ ( .D(n15556), .CP(wclk), .Q(ram[11315]) );
  DFF ram_reg_633__2_ ( .D(n15555), .CP(wclk), .Q(ram[11314]) );
  DFF ram_reg_633__1_ ( .D(n15554), .CP(wclk), .Q(ram[11313]) );
  DFF ram_reg_633__0_ ( .D(n15553), .CP(wclk), .Q(ram[11312]) );
  DFF ram_reg_637__7_ ( .D(n15528), .CP(wclk), .Q(ram[11287]) );
  DFF ram_reg_637__6_ ( .D(n15527), .CP(wclk), .Q(ram[11286]) );
  DFF ram_reg_637__5_ ( .D(n15526), .CP(wclk), .Q(ram[11285]) );
  DFF ram_reg_637__4_ ( .D(n15525), .CP(wclk), .Q(ram[11284]) );
  DFF ram_reg_637__3_ ( .D(n15524), .CP(wclk), .Q(ram[11283]) );
  DFF ram_reg_637__2_ ( .D(n15523), .CP(wclk), .Q(ram[11282]) );
  DFF ram_reg_637__1_ ( .D(n15522), .CP(wclk), .Q(ram[11281]) );
  DFF ram_reg_637__0_ ( .D(n15521), .CP(wclk), .Q(ram[11280]) );
  DFF ram_reg_641__7_ ( .D(n15496), .CP(wclk), .Q(ram[11255]) );
  DFF ram_reg_641__6_ ( .D(n15495), .CP(wclk), .Q(ram[11254]) );
  DFF ram_reg_641__5_ ( .D(n15494), .CP(wclk), .Q(ram[11253]) );
  DFF ram_reg_641__4_ ( .D(n15493), .CP(wclk), .Q(ram[11252]) );
  DFF ram_reg_641__3_ ( .D(n15492), .CP(wclk), .Q(ram[11251]) );
  DFF ram_reg_641__2_ ( .D(n15491), .CP(wclk), .Q(ram[11250]) );
  DFF ram_reg_641__1_ ( .D(n15490), .CP(wclk), .Q(ram[11249]) );
  DFF ram_reg_641__0_ ( .D(n15489), .CP(wclk), .Q(ram[11248]) );
  DFF ram_reg_645__7_ ( .D(n15464), .CP(wclk), .Q(ram[11223]) );
  DFF ram_reg_645__6_ ( .D(n15463), .CP(wclk), .Q(ram[11222]) );
  DFF ram_reg_645__5_ ( .D(n15462), .CP(wclk), .Q(ram[11221]) );
  DFF ram_reg_645__4_ ( .D(n15461), .CP(wclk), .Q(ram[11220]) );
  DFF ram_reg_645__3_ ( .D(n15460), .CP(wclk), .Q(ram[11219]) );
  DFF ram_reg_645__2_ ( .D(n15459), .CP(wclk), .Q(ram[11218]) );
  DFF ram_reg_645__1_ ( .D(n15458), .CP(wclk), .Q(ram[11217]) );
  DFF ram_reg_645__0_ ( .D(n15457), .CP(wclk), .Q(ram[11216]) );
  DFF ram_reg_649__7_ ( .D(n15432), .CP(wclk), .Q(ram[11191]) );
  DFF ram_reg_649__6_ ( .D(n15431), .CP(wclk), .Q(ram[11190]) );
  DFF ram_reg_649__5_ ( .D(n15430), .CP(wclk), .Q(ram[11189]) );
  DFF ram_reg_649__4_ ( .D(n15429), .CP(wclk), .Q(ram[11188]) );
  DFF ram_reg_649__3_ ( .D(n15428), .CP(wclk), .Q(ram[11187]) );
  DFF ram_reg_649__2_ ( .D(n15427), .CP(wclk), .Q(ram[11186]) );
  DFF ram_reg_649__1_ ( .D(n15426), .CP(wclk), .Q(ram[11185]) );
  DFF ram_reg_649__0_ ( .D(n15425), .CP(wclk), .Q(ram[11184]) );
  DFF ram_reg_653__7_ ( .D(n15400), .CP(wclk), .Q(ram[11159]) );
  DFF ram_reg_653__6_ ( .D(n15399), .CP(wclk), .Q(ram[11158]) );
  DFF ram_reg_653__5_ ( .D(n15398), .CP(wclk), .Q(ram[11157]) );
  DFF ram_reg_653__4_ ( .D(n15397), .CP(wclk), .Q(ram[11156]) );
  DFF ram_reg_653__3_ ( .D(n15396), .CP(wclk), .Q(ram[11155]) );
  DFF ram_reg_653__2_ ( .D(n15395), .CP(wclk), .Q(ram[11154]) );
  DFF ram_reg_653__1_ ( .D(n15394), .CP(wclk), .Q(ram[11153]) );
  DFF ram_reg_653__0_ ( .D(n15393), .CP(wclk), .Q(ram[11152]) );
  DFF ram_reg_657__7_ ( .D(n15368), .CP(wclk), .Q(ram[11127]) );
  DFF ram_reg_657__6_ ( .D(n15367), .CP(wclk), .Q(ram[11126]) );
  DFF ram_reg_657__5_ ( .D(n15366), .CP(wclk), .Q(ram[11125]) );
  DFF ram_reg_657__4_ ( .D(n15365), .CP(wclk), .Q(ram[11124]) );
  DFF ram_reg_657__3_ ( .D(n15364), .CP(wclk), .Q(ram[11123]) );
  DFF ram_reg_657__2_ ( .D(n15363), .CP(wclk), .Q(ram[11122]) );
  DFF ram_reg_657__1_ ( .D(n15362), .CP(wclk), .Q(ram[11121]) );
  DFF ram_reg_657__0_ ( .D(n15361), .CP(wclk), .Q(ram[11120]) );
  DFF ram_reg_665__7_ ( .D(n15304), .CP(wclk), .Q(ram[11063]) );
  DFF ram_reg_665__6_ ( .D(n15303), .CP(wclk), .Q(ram[11062]) );
  DFF ram_reg_665__5_ ( .D(n15302), .CP(wclk), .Q(ram[11061]) );
  DFF ram_reg_665__4_ ( .D(n15301), .CP(wclk), .Q(ram[11060]) );
  DFF ram_reg_665__3_ ( .D(n15300), .CP(wclk), .Q(ram[11059]) );
  DFF ram_reg_665__2_ ( .D(n15299), .CP(wclk), .Q(ram[11058]) );
  DFF ram_reg_665__1_ ( .D(n15298), .CP(wclk), .Q(ram[11057]) );
  DFF ram_reg_665__0_ ( .D(n15297), .CP(wclk), .Q(ram[11056]) );
  DFF ram_reg_669__7_ ( .D(n15272), .CP(wclk), .Q(ram[11031]) );
  DFF ram_reg_669__6_ ( .D(n15271), .CP(wclk), .Q(ram[11030]) );
  DFF ram_reg_669__5_ ( .D(n15270), .CP(wclk), .Q(ram[11029]) );
  DFF ram_reg_669__4_ ( .D(n15269), .CP(wclk), .Q(ram[11028]) );
  DFF ram_reg_669__3_ ( .D(n15268), .CP(wclk), .Q(ram[11027]) );
  DFF ram_reg_669__2_ ( .D(n15267), .CP(wclk), .Q(ram[11026]) );
  DFF ram_reg_669__1_ ( .D(n15266), .CP(wclk), .Q(ram[11025]) );
  DFF ram_reg_669__0_ ( .D(n15265), .CP(wclk), .Q(ram[11024]) );
  DFF ram_reg_673__7_ ( .D(n15240), .CP(wclk), .Q(ram[10999]) );
  DFF ram_reg_673__6_ ( .D(n15239), .CP(wclk), .Q(ram[10998]) );
  DFF ram_reg_673__5_ ( .D(n15238), .CP(wclk), .Q(ram[10997]) );
  DFF ram_reg_673__4_ ( .D(n15237), .CP(wclk), .Q(ram[10996]) );
  DFF ram_reg_673__3_ ( .D(n15236), .CP(wclk), .Q(ram[10995]) );
  DFF ram_reg_673__2_ ( .D(n15235), .CP(wclk), .Q(ram[10994]) );
  DFF ram_reg_673__1_ ( .D(n15234), .CP(wclk), .Q(ram[10993]) );
  DFF ram_reg_673__0_ ( .D(n15233), .CP(wclk), .Q(ram[10992]) );
  DFF ram_reg_677__7_ ( .D(n15208), .CP(wclk), .Q(ram[10967]) );
  DFF ram_reg_677__6_ ( .D(n15207), .CP(wclk), .Q(ram[10966]) );
  DFF ram_reg_677__5_ ( .D(n15206), .CP(wclk), .Q(ram[10965]) );
  DFF ram_reg_677__4_ ( .D(n15205), .CP(wclk), .Q(ram[10964]) );
  DFF ram_reg_677__3_ ( .D(n15204), .CP(wclk), .Q(ram[10963]) );
  DFF ram_reg_677__2_ ( .D(n15203), .CP(wclk), .Q(ram[10962]) );
  DFF ram_reg_677__1_ ( .D(n15202), .CP(wclk), .Q(ram[10961]) );
  DFF ram_reg_677__0_ ( .D(n15201), .CP(wclk), .Q(ram[10960]) );
  DFF ram_reg_681__7_ ( .D(n15176), .CP(wclk), .Q(ram[10935]) );
  DFF ram_reg_681__6_ ( .D(n15175), .CP(wclk), .Q(ram[10934]) );
  DFF ram_reg_681__5_ ( .D(n15174), .CP(wclk), .Q(ram[10933]) );
  DFF ram_reg_681__4_ ( .D(n15173), .CP(wclk), .Q(ram[10932]) );
  DFF ram_reg_681__3_ ( .D(n15172), .CP(wclk), .Q(ram[10931]) );
  DFF ram_reg_681__2_ ( .D(n15171), .CP(wclk), .Q(ram[10930]) );
  DFF ram_reg_681__1_ ( .D(n15170), .CP(wclk), .Q(ram[10929]) );
  DFF ram_reg_681__0_ ( .D(n15169), .CP(wclk), .Q(ram[10928]) );
  DFF ram_reg_685__7_ ( .D(n15144), .CP(wclk), .Q(ram[10903]) );
  DFF ram_reg_685__6_ ( .D(n15143), .CP(wclk), .Q(ram[10902]) );
  DFF ram_reg_685__5_ ( .D(n15142), .CP(wclk), .Q(ram[10901]) );
  DFF ram_reg_685__4_ ( .D(n15141), .CP(wclk), .Q(ram[10900]) );
  DFF ram_reg_685__3_ ( .D(n15140), .CP(wclk), .Q(ram[10899]) );
  DFF ram_reg_685__2_ ( .D(n15139), .CP(wclk), .Q(ram[10898]) );
  DFF ram_reg_685__1_ ( .D(n15138), .CP(wclk), .Q(ram[10897]) );
  DFF ram_reg_685__0_ ( .D(n15137), .CP(wclk), .Q(ram[10896]) );
  DFF ram_reg_689__7_ ( .D(n15112), .CP(wclk), .Q(ram[10871]) );
  DFF ram_reg_689__6_ ( .D(n15111), .CP(wclk), .Q(ram[10870]) );
  DFF ram_reg_689__5_ ( .D(n15110), .CP(wclk), .Q(ram[10869]) );
  DFF ram_reg_689__4_ ( .D(n15109), .CP(wclk), .Q(ram[10868]) );
  DFF ram_reg_689__3_ ( .D(n15108), .CP(wclk), .Q(ram[10867]) );
  DFF ram_reg_689__2_ ( .D(n15107), .CP(wclk), .Q(ram[10866]) );
  DFF ram_reg_689__1_ ( .D(n15106), .CP(wclk), .Q(ram[10865]) );
  DFF ram_reg_689__0_ ( .D(n15105), .CP(wclk), .Q(ram[10864]) );
  DFF ram_reg_693__7_ ( .D(n15080), .CP(wclk), .Q(ram[10839]) );
  DFF ram_reg_693__6_ ( .D(n15079), .CP(wclk), .Q(ram[10838]) );
  DFF ram_reg_693__5_ ( .D(n15078), .CP(wclk), .Q(ram[10837]) );
  DFF ram_reg_693__4_ ( .D(n15077), .CP(wclk), .Q(ram[10836]) );
  DFF ram_reg_693__3_ ( .D(n15076), .CP(wclk), .Q(ram[10835]) );
  DFF ram_reg_693__2_ ( .D(n15075), .CP(wclk), .Q(ram[10834]) );
  DFF ram_reg_693__1_ ( .D(n15074), .CP(wclk), .Q(ram[10833]) );
  DFF ram_reg_693__0_ ( .D(n15073), .CP(wclk), .Q(ram[10832]) );
  DFF ram_reg_697__7_ ( .D(n15048), .CP(wclk), .Q(ram[10807]) );
  DFF ram_reg_697__6_ ( .D(n15047), .CP(wclk), .Q(ram[10806]) );
  DFF ram_reg_697__5_ ( .D(n15046), .CP(wclk), .Q(ram[10805]) );
  DFF ram_reg_697__4_ ( .D(n15045), .CP(wclk), .Q(ram[10804]) );
  DFF ram_reg_697__3_ ( .D(n15044), .CP(wclk), .Q(ram[10803]) );
  DFF ram_reg_697__2_ ( .D(n15043), .CP(wclk), .Q(ram[10802]) );
  DFF ram_reg_697__1_ ( .D(n15042), .CP(wclk), .Q(ram[10801]) );
  DFF ram_reg_697__0_ ( .D(n15041), .CP(wclk), .Q(ram[10800]) );
  DFF ram_reg_701__7_ ( .D(n15016), .CP(wclk), .Q(ram[10775]) );
  DFF ram_reg_701__6_ ( .D(n15015), .CP(wclk), .Q(ram[10774]) );
  DFF ram_reg_701__5_ ( .D(n15014), .CP(wclk), .Q(ram[10773]) );
  DFF ram_reg_701__4_ ( .D(n15013), .CP(wclk), .Q(ram[10772]) );
  DFF ram_reg_701__3_ ( .D(n15012), .CP(wclk), .Q(ram[10771]) );
  DFF ram_reg_701__2_ ( .D(n15011), .CP(wclk), .Q(ram[10770]) );
  DFF ram_reg_701__1_ ( .D(n15010), .CP(wclk), .Q(ram[10769]) );
  DFF ram_reg_701__0_ ( .D(n15009), .CP(wclk), .Q(ram[10768]) );
  DFF ram_reg_705__7_ ( .D(n14984), .CP(wclk), .Q(ram[10743]) );
  DFF ram_reg_705__6_ ( .D(n14983), .CP(wclk), .Q(ram[10742]) );
  DFF ram_reg_705__5_ ( .D(n14982), .CP(wclk), .Q(ram[10741]) );
  DFF ram_reg_705__4_ ( .D(n14981), .CP(wclk), .Q(ram[10740]) );
  DFF ram_reg_705__3_ ( .D(n14980), .CP(wclk), .Q(ram[10739]) );
  DFF ram_reg_705__2_ ( .D(n14979), .CP(wclk), .Q(ram[10738]) );
  DFF ram_reg_705__1_ ( .D(n14978), .CP(wclk), .Q(ram[10737]) );
  DFF ram_reg_705__0_ ( .D(n14977), .CP(wclk), .Q(ram[10736]) );
  DFF ram_reg_713__7_ ( .D(n14920), .CP(wclk), .Q(ram[10679]) );
  DFF ram_reg_713__6_ ( .D(n14919), .CP(wclk), .Q(ram[10678]) );
  DFF ram_reg_713__5_ ( .D(n14918), .CP(wclk), .Q(ram[10677]) );
  DFF ram_reg_713__4_ ( .D(n14917), .CP(wclk), .Q(ram[10676]) );
  DFF ram_reg_713__3_ ( .D(n14916), .CP(wclk), .Q(ram[10675]) );
  DFF ram_reg_713__2_ ( .D(n14915), .CP(wclk), .Q(ram[10674]) );
  DFF ram_reg_713__1_ ( .D(n14914), .CP(wclk), .Q(ram[10673]) );
  DFF ram_reg_713__0_ ( .D(n14913), .CP(wclk), .Q(ram[10672]) );
  DFF ram_reg_717__7_ ( .D(n14888), .CP(wclk), .Q(ram[10647]) );
  DFF ram_reg_717__6_ ( .D(n14887), .CP(wclk), .Q(ram[10646]) );
  DFF ram_reg_717__5_ ( .D(n14886), .CP(wclk), .Q(ram[10645]) );
  DFF ram_reg_717__4_ ( .D(n14885), .CP(wclk), .Q(ram[10644]) );
  DFF ram_reg_717__3_ ( .D(n14884), .CP(wclk), .Q(ram[10643]) );
  DFF ram_reg_717__2_ ( .D(n14883), .CP(wclk), .Q(ram[10642]) );
  DFF ram_reg_717__1_ ( .D(n14882), .CP(wclk), .Q(ram[10641]) );
  DFF ram_reg_717__0_ ( .D(n14881), .CP(wclk), .Q(ram[10640]) );
  DFF ram_reg_721__7_ ( .D(n14856), .CP(wclk), .Q(ram[10615]) );
  DFF ram_reg_721__6_ ( .D(n14855), .CP(wclk), .Q(ram[10614]) );
  DFF ram_reg_721__5_ ( .D(n14854), .CP(wclk), .Q(ram[10613]) );
  DFF ram_reg_721__4_ ( .D(n14853), .CP(wclk), .Q(ram[10612]) );
  DFF ram_reg_721__3_ ( .D(n14852), .CP(wclk), .Q(ram[10611]) );
  DFF ram_reg_721__2_ ( .D(n14851), .CP(wclk), .Q(ram[10610]) );
  DFF ram_reg_721__1_ ( .D(n14850), .CP(wclk), .Q(ram[10609]) );
  DFF ram_reg_721__0_ ( .D(n14849), .CP(wclk), .Q(ram[10608]) );
  DFF ram_reg_729__7_ ( .D(n14792), .CP(wclk), .Q(ram[10551]) );
  DFF ram_reg_729__6_ ( .D(n14791), .CP(wclk), .Q(ram[10550]) );
  DFF ram_reg_729__5_ ( .D(n14790), .CP(wclk), .Q(ram[10549]) );
  DFF ram_reg_729__4_ ( .D(n14789), .CP(wclk), .Q(ram[10548]) );
  DFF ram_reg_729__3_ ( .D(n14788), .CP(wclk), .Q(ram[10547]) );
  DFF ram_reg_729__2_ ( .D(n14787), .CP(wclk), .Q(ram[10546]) );
  DFF ram_reg_729__1_ ( .D(n14786), .CP(wclk), .Q(ram[10545]) );
  DFF ram_reg_729__0_ ( .D(n14785), .CP(wclk), .Q(ram[10544]) );
  DFF ram_reg_733__7_ ( .D(n14760), .CP(wclk), .Q(ram[10519]) );
  DFF ram_reg_733__6_ ( .D(n14759), .CP(wclk), .Q(ram[10518]) );
  DFF ram_reg_733__5_ ( .D(n14758), .CP(wclk), .Q(ram[10517]) );
  DFF ram_reg_733__4_ ( .D(n14757), .CP(wclk), .Q(ram[10516]) );
  DFF ram_reg_733__3_ ( .D(n14756), .CP(wclk), .Q(ram[10515]) );
  DFF ram_reg_733__2_ ( .D(n14755), .CP(wclk), .Q(ram[10514]) );
  DFF ram_reg_733__1_ ( .D(n14754), .CP(wclk), .Q(ram[10513]) );
  DFF ram_reg_733__0_ ( .D(n14753), .CP(wclk), .Q(ram[10512]) );
  DFF ram_reg_737__7_ ( .D(n14728), .CP(wclk), .Q(ram[10487]) );
  DFF ram_reg_737__6_ ( .D(n14727), .CP(wclk), .Q(ram[10486]) );
  DFF ram_reg_737__5_ ( .D(n14726), .CP(wclk), .Q(ram[10485]) );
  DFF ram_reg_737__4_ ( .D(n14725), .CP(wclk), .Q(ram[10484]) );
  DFF ram_reg_737__3_ ( .D(n14724), .CP(wclk), .Q(ram[10483]) );
  DFF ram_reg_737__2_ ( .D(n14723), .CP(wclk), .Q(ram[10482]) );
  DFF ram_reg_737__1_ ( .D(n14722), .CP(wclk), .Q(ram[10481]) );
  DFF ram_reg_737__0_ ( .D(n14721), .CP(wclk), .Q(ram[10480]) );
  DFF ram_reg_741__7_ ( .D(n14696), .CP(wclk), .Q(ram[10455]) );
  DFF ram_reg_741__6_ ( .D(n14695), .CP(wclk), .Q(ram[10454]) );
  DFF ram_reg_741__5_ ( .D(n14694), .CP(wclk), .Q(ram[10453]) );
  DFF ram_reg_741__4_ ( .D(n14693), .CP(wclk), .Q(ram[10452]) );
  DFF ram_reg_741__3_ ( .D(n14692), .CP(wclk), .Q(ram[10451]) );
  DFF ram_reg_741__2_ ( .D(n14691), .CP(wclk), .Q(ram[10450]) );
  DFF ram_reg_741__1_ ( .D(n14690), .CP(wclk), .Q(ram[10449]) );
  DFF ram_reg_741__0_ ( .D(n14689), .CP(wclk), .Q(ram[10448]) );
  DFF ram_reg_745__7_ ( .D(n14664), .CP(wclk), .Q(ram[10423]) );
  DFF ram_reg_745__6_ ( .D(n14663), .CP(wclk), .Q(ram[10422]) );
  DFF ram_reg_745__5_ ( .D(n14662), .CP(wclk), .Q(ram[10421]) );
  DFF ram_reg_745__4_ ( .D(n14661), .CP(wclk), .Q(ram[10420]) );
  DFF ram_reg_745__3_ ( .D(n14660), .CP(wclk), .Q(ram[10419]) );
  DFF ram_reg_745__2_ ( .D(n14659), .CP(wclk), .Q(ram[10418]) );
  DFF ram_reg_745__1_ ( .D(n14658), .CP(wclk), .Q(ram[10417]) );
  DFF ram_reg_745__0_ ( .D(n14657), .CP(wclk), .Q(ram[10416]) );
  DFF ram_reg_749__7_ ( .D(n14632), .CP(wclk), .Q(ram[10391]) );
  DFF ram_reg_749__6_ ( .D(n14631), .CP(wclk), .Q(ram[10390]) );
  DFF ram_reg_749__5_ ( .D(n14630), .CP(wclk), .Q(ram[10389]) );
  DFF ram_reg_749__4_ ( .D(n14629), .CP(wclk), .Q(ram[10388]) );
  DFF ram_reg_749__3_ ( .D(n14628), .CP(wclk), .Q(ram[10387]) );
  DFF ram_reg_749__2_ ( .D(n14627), .CP(wclk), .Q(ram[10386]) );
  DFF ram_reg_749__1_ ( .D(n14626), .CP(wclk), .Q(ram[10385]) );
  DFF ram_reg_749__0_ ( .D(n14625), .CP(wclk), .Q(ram[10384]) );
  DFF ram_reg_753__7_ ( .D(n14600), .CP(wclk), .Q(ram[10359]) );
  DFF ram_reg_753__6_ ( .D(n14599), .CP(wclk), .Q(ram[10358]) );
  DFF ram_reg_753__5_ ( .D(n14598), .CP(wclk), .Q(ram[10357]) );
  DFF ram_reg_753__4_ ( .D(n14597), .CP(wclk), .Q(ram[10356]) );
  DFF ram_reg_753__3_ ( .D(n14596), .CP(wclk), .Q(ram[10355]) );
  DFF ram_reg_753__2_ ( .D(n14595), .CP(wclk), .Q(ram[10354]) );
  DFF ram_reg_753__1_ ( .D(n14594), .CP(wclk), .Q(ram[10353]) );
  DFF ram_reg_753__0_ ( .D(n14593), .CP(wclk), .Q(ram[10352]) );
  DFF ram_reg_757__7_ ( .D(n14568), .CP(wclk), .Q(ram[10327]) );
  DFF ram_reg_757__6_ ( .D(n14567), .CP(wclk), .Q(ram[10326]) );
  DFF ram_reg_757__5_ ( .D(n14566), .CP(wclk), .Q(ram[10325]) );
  DFF ram_reg_757__4_ ( .D(n14565), .CP(wclk), .Q(ram[10324]) );
  DFF ram_reg_757__3_ ( .D(n14564), .CP(wclk), .Q(ram[10323]) );
  DFF ram_reg_757__2_ ( .D(n14563), .CP(wclk), .Q(ram[10322]) );
  DFF ram_reg_757__1_ ( .D(n14562), .CP(wclk), .Q(ram[10321]) );
  DFF ram_reg_757__0_ ( .D(n14561), .CP(wclk), .Q(ram[10320]) );
  DFF ram_reg_761__7_ ( .D(n14536), .CP(wclk), .Q(ram[10295]) );
  DFF ram_reg_761__6_ ( .D(n14535), .CP(wclk), .Q(ram[10294]) );
  DFF ram_reg_761__5_ ( .D(n14534), .CP(wclk), .Q(ram[10293]) );
  DFF ram_reg_761__4_ ( .D(n14533), .CP(wclk), .Q(ram[10292]) );
  DFF ram_reg_761__3_ ( .D(n14532), .CP(wclk), .Q(ram[10291]) );
  DFF ram_reg_761__2_ ( .D(n14531), .CP(wclk), .Q(ram[10290]) );
  DFF ram_reg_761__1_ ( .D(n14530), .CP(wclk), .Q(ram[10289]) );
  DFF ram_reg_761__0_ ( .D(n14529), .CP(wclk), .Q(ram[10288]) );
  DFF ram_reg_765__7_ ( .D(n14504), .CP(wclk), .Q(ram[10263]) );
  DFF ram_reg_765__6_ ( .D(n14503), .CP(wclk), .Q(ram[10262]) );
  DFF ram_reg_765__5_ ( .D(n14502), .CP(wclk), .Q(ram[10261]) );
  DFF ram_reg_765__4_ ( .D(n14501), .CP(wclk), .Q(ram[10260]) );
  DFF ram_reg_765__3_ ( .D(n14500), .CP(wclk), .Q(ram[10259]) );
  DFF ram_reg_765__2_ ( .D(n14499), .CP(wclk), .Q(ram[10258]) );
  DFF ram_reg_765__1_ ( .D(n14498), .CP(wclk), .Q(ram[10257]) );
  DFF ram_reg_765__0_ ( .D(n14497), .CP(wclk), .Q(ram[10256]) );
  DFF ram_reg_777__7_ ( .D(n14408), .CP(wclk), .Q(ram[10167]) );
  DFF ram_reg_777__6_ ( .D(n14407), .CP(wclk), .Q(ram[10166]) );
  DFF ram_reg_777__5_ ( .D(n14406), .CP(wclk), .Q(ram[10165]) );
  DFF ram_reg_777__4_ ( .D(n14405), .CP(wclk), .Q(ram[10164]) );
  DFF ram_reg_777__3_ ( .D(n14404), .CP(wclk), .Q(ram[10163]) );
  DFF ram_reg_777__2_ ( .D(n14403), .CP(wclk), .Q(ram[10162]) );
  DFF ram_reg_777__1_ ( .D(n14402), .CP(wclk), .Q(ram[10161]) );
  DFF ram_reg_777__0_ ( .D(n14401), .CP(wclk), .Q(ram[10160]) );
  DFF ram_reg_781__7_ ( .D(n14376), .CP(wclk), .Q(ram[10135]) );
  DFF ram_reg_781__6_ ( .D(n14375), .CP(wclk), .Q(ram[10134]) );
  DFF ram_reg_781__5_ ( .D(n14374), .CP(wclk), .Q(ram[10133]) );
  DFF ram_reg_781__4_ ( .D(n14373), .CP(wclk), .Q(ram[10132]) );
  DFF ram_reg_781__3_ ( .D(n14372), .CP(wclk), .Q(ram[10131]) );
  DFF ram_reg_781__2_ ( .D(n14371), .CP(wclk), .Q(ram[10130]) );
  DFF ram_reg_781__1_ ( .D(n14370), .CP(wclk), .Q(ram[10129]) );
  DFF ram_reg_781__0_ ( .D(n14369), .CP(wclk), .Q(ram[10128]) );
  DFF ram_reg_793__7_ ( .D(n14280), .CP(wclk), .Q(ram[10039]) );
  DFF ram_reg_793__6_ ( .D(n14279), .CP(wclk), .Q(ram[10038]) );
  DFF ram_reg_793__5_ ( .D(n14278), .CP(wclk), .Q(ram[10037]) );
  DFF ram_reg_793__4_ ( .D(n14277), .CP(wclk), .Q(ram[10036]) );
  DFF ram_reg_793__3_ ( .D(n14276), .CP(wclk), .Q(ram[10035]) );
  DFF ram_reg_793__2_ ( .D(n14275), .CP(wclk), .Q(ram[10034]) );
  DFF ram_reg_793__1_ ( .D(n14274), .CP(wclk), .Q(ram[10033]) );
  DFF ram_reg_793__0_ ( .D(n14273), .CP(wclk), .Q(ram[10032]) );
  DFF ram_reg_797__7_ ( .D(n14248), .CP(wclk), .Q(ram[10007]) );
  DFF ram_reg_797__6_ ( .D(n14247), .CP(wclk), .Q(ram[10006]) );
  DFF ram_reg_797__5_ ( .D(n14246), .CP(wclk), .Q(ram[10005]) );
  DFF ram_reg_797__4_ ( .D(n14245), .CP(wclk), .Q(ram[10004]) );
  DFF ram_reg_797__3_ ( .D(n14244), .CP(wclk), .Q(ram[10003]) );
  DFF ram_reg_797__2_ ( .D(n14243), .CP(wclk), .Q(ram[10002]) );
  DFF ram_reg_797__1_ ( .D(n14242), .CP(wclk), .Q(ram[10001]) );
  DFF ram_reg_797__0_ ( .D(n14241), .CP(wclk), .Q(ram[10000]) );
  DFF ram_reg_801__7_ ( .D(n14216), .CP(wclk), .Q(ram[9975]) );
  DFF ram_reg_801__6_ ( .D(n14215), .CP(wclk), .Q(ram[9974]) );
  DFF ram_reg_801__5_ ( .D(n14214), .CP(wclk), .Q(ram[9973]) );
  DFF ram_reg_801__4_ ( .D(n14213), .CP(wclk), .Q(ram[9972]) );
  DFF ram_reg_801__3_ ( .D(n14212), .CP(wclk), .Q(ram[9971]) );
  DFF ram_reg_801__2_ ( .D(n14211), .CP(wclk), .Q(ram[9970]) );
  DFF ram_reg_801__1_ ( .D(n14210), .CP(wclk), .Q(ram[9969]) );
  DFF ram_reg_801__0_ ( .D(n14209), .CP(wclk), .Q(ram[9968]) );
  DFF ram_reg_809__7_ ( .D(n14152), .CP(wclk), .Q(ram[9911]) );
  DFF ram_reg_809__6_ ( .D(n14151), .CP(wclk), .Q(ram[9910]) );
  DFF ram_reg_809__5_ ( .D(n14150), .CP(wclk), .Q(ram[9909]) );
  DFF ram_reg_809__4_ ( .D(n14149), .CP(wclk), .Q(ram[9908]) );
  DFF ram_reg_809__3_ ( .D(n14148), .CP(wclk), .Q(ram[9907]) );
  DFF ram_reg_809__2_ ( .D(n14147), .CP(wclk), .Q(ram[9906]) );
  DFF ram_reg_809__1_ ( .D(n14146), .CP(wclk), .Q(ram[9905]) );
  DFF ram_reg_809__0_ ( .D(n14145), .CP(wclk), .Q(ram[9904]) );
  DFF ram_reg_813__7_ ( .D(n14120), .CP(wclk), .Q(ram[9879]) );
  DFF ram_reg_813__6_ ( .D(n14119), .CP(wclk), .Q(ram[9878]) );
  DFF ram_reg_813__5_ ( .D(n14118), .CP(wclk), .Q(ram[9877]) );
  DFF ram_reg_813__4_ ( .D(n14117), .CP(wclk), .Q(ram[9876]) );
  DFF ram_reg_813__3_ ( .D(n14116), .CP(wclk), .Q(ram[9875]) );
  DFF ram_reg_813__2_ ( .D(n14115), .CP(wclk), .Q(ram[9874]) );
  DFF ram_reg_813__1_ ( .D(n14114), .CP(wclk), .Q(ram[9873]) );
  DFF ram_reg_813__0_ ( .D(n14113), .CP(wclk), .Q(ram[9872]) );
  DFF ram_reg_817__7_ ( .D(n14088), .CP(wclk), .Q(ram[9847]) );
  DFF ram_reg_817__6_ ( .D(n14087), .CP(wclk), .Q(ram[9846]) );
  DFF ram_reg_817__5_ ( .D(n14086), .CP(wclk), .Q(ram[9845]) );
  DFF ram_reg_817__4_ ( .D(n14085), .CP(wclk), .Q(ram[9844]) );
  DFF ram_reg_817__3_ ( .D(n14084), .CP(wclk), .Q(ram[9843]) );
  DFF ram_reg_817__2_ ( .D(n14083), .CP(wclk), .Q(ram[9842]) );
  DFF ram_reg_817__1_ ( .D(n14082), .CP(wclk), .Q(ram[9841]) );
  DFF ram_reg_817__0_ ( .D(n14081), .CP(wclk), .Q(ram[9840]) );
  DFF ram_reg_825__7_ ( .D(n14024), .CP(wclk), .Q(ram[9783]) );
  DFF ram_reg_825__6_ ( .D(n14023), .CP(wclk), .Q(ram[9782]) );
  DFF ram_reg_825__5_ ( .D(n14022), .CP(wclk), .Q(ram[9781]) );
  DFF ram_reg_825__4_ ( .D(n14021), .CP(wclk), .Q(ram[9780]) );
  DFF ram_reg_825__3_ ( .D(n14020), .CP(wclk), .Q(ram[9779]) );
  DFF ram_reg_825__2_ ( .D(n14019), .CP(wclk), .Q(ram[9778]) );
  DFF ram_reg_825__1_ ( .D(n14018), .CP(wclk), .Q(ram[9777]) );
  DFF ram_reg_825__0_ ( .D(n14017), .CP(wclk), .Q(ram[9776]) );
  DFF ram_reg_829__7_ ( .D(n13992), .CP(wclk), .Q(ram[9751]) );
  DFF ram_reg_829__6_ ( .D(n13991), .CP(wclk), .Q(ram[9750]) );
  DFF ram_reg_829__5_ ( .D(n13990), .CP(wclk), .Q(ram[9749]) );
  DFF ram_reg_829__4_ ( .D(n13989), .CP(wclk), .Q(ram[9748]) );
  DFF ram_reg_829__3_ ( .D(n13988), .CP(wclk), .Q(ram[9747]) );
  DFF ram_reg_829__2_ ( .D(n13987), .CP(wclk), .Q(ram[9746]) );
  DFF ram_reg_829__1_ ( .D(n13986), .CP(wclk), .Q(ram[9745]) );
  DFF ram_reg_829__0_ ( .D(n13985), .CP(wclk), .Q(ram[9744]) );
  DFF ram_reg_841__7_ ( .D(n13896), .CP(wclk), .Q(ram[9655]) );
  DFF ram_reg_841__6_ ( .D(n13895), .CP(wclk), .Q(ram[9654]) );
  DFF ram_reg_841__5_ ( .D(n13894), .CP(wclk), .Q(ram[9653]) );
  DFF ram_reg_841__4_ ( .D(n13893), .CP(wclk), .Q(ram[9652]) );
  DFF ram_reg_841__3_ ( .D(n13892), .CP(wclk), .Q(ram[9651]) );
  DFF ram_reg_841__2_ ( .D(n13891), .CP(wclk), .Q(ram[9650]) );
  DFF ram_reg_841__1_ ( .D(n13890), .CP(wclk), .Q(ram[9649]) );
  DFF ram_reg_841__0_ ( .D(n13889), .CP(wclk), .Q(ram[9648]) );
  DFF ram_reg_873__7_ ( .D(n13640), .CP(wclk), .Q(ram[9399]) );
  DFF ram_reg_873__6_ ( .D(n13639), .CP(wclk), .Q(ram[9398]) );
  DFF ram_reg_873__5_ ( .D(n13638), .CP(wclk), .Q(ram[9397]) );
  DFF ram_reg_873__4_ ( .D(n13637), .CP(wclk), .Q(ram[9396]) );
  DFF ram_reg_873__3_ ( .D(n13636), .CP(wclk), .Q(ram[9395]) );
  DFF ram_reg_873__2_ ( .D(n13635), .CP(wclk), .Q(ram[9394]) );
  DFF ram_reg_873__1_ ( .D(n13634), .CP(wclk), .Q(ram[9393]) );
  DFF ram_reg_873__0_ ( .D(n13633), .CP(wclk), .Q(ram[9392]) );
  DFF ram_reg_877__7_ ( .D(n13608), .CP(wclk), .Q(ram[9367]) );
  DFF ram_reg_877__6_ ( .D(n13607), .CP(wclk), .Q(ram[9366]) );
  DFF ram_reg_877__5_ ( .D(n13606), .CP(wclk), .Q(ram[9365]) );
  DFF ram_reg_877__4_ ( .D(n13605), .CP(wclk), .Q(ram[9364]) );
  DFF ram_reg_877__3_ ( .D(n13604), .CP(wclk), .Q(ram[9363]) );
  DFF ram_reg_877__2_ ( .D(n13603), .CP(wclk), .Q(ram[9362]) );
  DFF ram_reg_877__1_ ( .D(n13602), .CP(wclk), .Q(ram[9361]) );
  DFF ram_reg_877__0_ ( .D(n13601), .CP(wclk), .Q(ram[9360]) );
  DFF ram_reg_889__7_ ( .D(n13512), .CP(wclk), .Q(ram[9271]) );
  DFF ram_reg_889__6_ ( .D(n13511), .CP(wclk), .Q(ram[9270]) );
  DFF ram_reg_889__5_ ( .D(n13510), .CP(wclk), .Q(ram[9269]) );
  DFF ram_reg_889__4_ ( .D(n13509), .CP(wclk), .Q(ram[9268]) );
  DFF ram_reg_889__3_ ( .D(n13508), .CP(wclk), .Q(ram[9267]) );
  DFF ram_reg_889__2_ ( .D(n13507), .CP(wclk), .Q(ram[9266]) );
  DFF ram_reg_889__1_ ( .D(n13506), .CP(wclk), .Q(ram[9265]) );
  DFF ram_reg_889__0_ ( .D(n13505), .CP(wclk), .Q(ram[9264]) );
  DFF ram_reg_893__7_ ( .D(n13480), .CP(wclk), .Q(ram[9239]) );
  DFF ram_reg_893__6_ ( .D(n13479), .CP(wclk), .Q(ram[9238]) );
  DFF ram_reg_893__5_ ( .D(n13478), .CP(wclk), .Q(ram[9237]) );
  DFF ram_reg_893__4_ ( .D(n13477), .CP(wclk), .Q(ram[9236]) );
  DFF ram_reg_893__3_ ( .D(n13476), .CP(wclk), .Q(ram[9235]) );
  DFF ram_reg_893__2_ ( .D(n13475), .CP(wclk), .Q(ram[9234]) );
  DFF ram_reg_893__1_ ( .D(n13474), .CP(wclk), .Q(ram[9233]) );
  DFF ram_reg_893__0_ ( .D(n13473), .CP(wclk), .Q(ram[9232]) );
  DFF ram_reg_897__7_ ( .D(n13448), .CP(wclk), .Q(ram[9207]) );
  DFF ram_reg_897__6_ ( .D(n13447), .CP(wclk), .Q(ram[9206]) );
  DFF ram_reg_897__5_ ( .D(n13446), .CP(wclk), .Q(ram[9205]) );
  DFF ram_reg_897__4_ ( .D(n13445), .CP(wclk), .Q(ram[9204]) );
  DFF ram_reg_897__3_ ( .D(n13444), .CP(wclk), .Q(ram[9203]) );
  DFF ram_reg_897__2_ ( .D(n13443), .CP(wclk), .Q(ram[9202]) );
  DFF ram_reg_897__1_ ( .D(n13442), .CP(wclk), .Q(ram[9201]) );
  DFF ram_reg_897__0_ ( .D(n13441), .CP(wclk), .Q(ram[9200]) );
  DFF ram_reg_901__7_ ( .D(n13416), .CP(wclk), .Q(ram[9175]) );
  DFF ram_reg_901__6_ ( .D(n13415), .CP(wclk), .Q(ram[9174]) );
  DFF ram_reg_901__5_ ( .D(n13414), .CP(wclk), .Q(ram[9173]) );
  DFF ram_reg_901__4_ ( .D(n13413), .CP(wclk), .Q(ram[9172]) );
  DFF ram_reg_901__3_ ( .D(n13412), .CP(wclk), .Q(ram[9171]) );
  DFF ram_reg_901__2_ ( .D(n13411), .CP(wclk), .Q(ram[9170]) );
  DFF ram_reg_901__1_ ( .D(n13410), .CP(wclk), .Q(ram[9169]) );
  DFF ram_reg_901__0_ ( .D(n13409), .CP(wclk), .Q(ram[9168]) );
  DFF ram_reg_905__7_ ( .D(n13384), .CP(wclk), .Q(ram[9143]) );
  DFF ram_reg_905__6_ ( .D(n13383), .CP(wclk), .Q(ram[9142]) );
  DFF ram_reg_905__5_ ( .D(n13382), .CP(wclk), .Q(ram[9141]) );
  DFF ram_reg_905__4_ ( .D(n13381), .CP(wclk), .Q(ram[9140]) );
  DFF ram_reg_905__3_ ( .D(n13380), .CP(wclk), .Q(ram[9139]) );
  DFF ram_reg_905__2_ ( .D(n13379), .CP(wclk), .Q(ram[9138]) );
  DFF ram_reg_905__1_ ( .D(n13378), .CP(wclk), .Q(ram[9137]) );
  DFF ram_reg_905__0_ ( .D(n13377), .CP(wclk), .Q(ram[9136]) );
  DFF ram_reg_909__7_ ( .D(n13352), .CP(wclk), .Q(ram[9111]) );
  DFF ram_reg_909__6_ ( .D(n13351), .CP(wclk), .Q(ram[9110]) );
  DFF ram_reg_909__5_ ( .D(n13350), .CP(wclk), .Q(ram[9109]) );
  DFF ram_reg_909__4_ ( .D(n13349), .CP(wclk), .Q(ram[9108]) );
  DFF ram_reg_909__3_ ( .D(n13348), .CP(wclk), .Q(ram[9107]) );
  DFF ram_reg_909__2_ ( .D(n13347), .CP(wclk), .Q(ram[9106]) );
  DFF ram_reg_909__1_ ( .D(n13346), .CP(wclk), .Q(ram[9105]) );
  DFF ram_reg_909__0_ ( .D(n13345), .CP(wclk), .Q(ram[9104]) );
  DFF ram_reg_913__7_ ( .D(n13320), .CP(wclk), .Q(ram[9079]) );
  DFF ram_reg_913__6_ ( .D(n13319), .CP(wclk), .Q(ram[9078]) );
  DFF ram_reg_913__5_ ( .D(n13318), .CP(wclk), .Q(ram[9077]) );
  DFF ram_reg_913__4_ ( .D(n13317), .CP(wclk), .Q(ram[9076]) );
  DFF ram_reg_913__3_ ( .D(n13316), .CP(wclk), .Q(ram[9075]) );
  DFF ram_reg_913__2_ ( .D(n13315), .CP(wclk), .Q(ram[9074]) );
  DFF ram_reg_913__1_ ( .D(n13314), .CP(wclk), .Q(ram[9073]) );
  DFF ram_reg_913__0_ ( .D(n13313), .CP(wclk), .Q(ram[9072]) );
  DFF ram_reg_921__7_ ( .D(n13256), .CP(wclk), .Q(ram[9015]) );
  DFF ram_reg_921__6_ ( .D(n13255), .CP(wclk), .Q(ram[9014]) );
  DFF ram_reg_921__5_ ( .D(n13254), .CP(wclk), .Q(ram[9013]) );
  DFF ram_reg_921__4_ ( .D(n13253), .CP(wclk), .Q(ram[9012]) );
  DFF ram_reg_921__3_ ( .D(n13252), .CP(wclk), .Q(ram[9011]) );
  DFF ram_reg_921__2_ ( .D(n13251), .CP(wclk), .Q(ram[9010]) );
  DFF ram_reg_921__1_ ( .D(n13250), .CP(wclk), .Q(ram[9009]) );
  DFF ram_reg_921__0_ ( .D(n13249), .CP(wclk), .Q(ram[9008]) );
  DFF ram_reg_925__7_ ( .D(n13224), .CP(wclk), .Q(ram[8983]) );
  DFF ram_reg_925__6_ ( .D(n13223), .CP(wclk), .Q(ram[8982]) );
  DFF ram_reg_925__5_ ( .D(n13222), .CP(wclk), .Q(ram[8981]) );
  DFF ram_reg_925__4_ ( .D(n13221), .CP(wclk), .Q(ram[8980]) );
  DFF ram_reg_925__3_ ( .D(n13220), .CP(wclk), .Q(ram[8979]) );
  DFF ram_reg_925__2_ ( .D(n13219), .CP(wclk), .Q(ram[8978]) );
  DFF ram_reg_925__1_ ( .D(n13218), .CP(wclk), .Q(ram[8977]) );
  DFF ram_reg_925__0_ ( .D(n13217), .CP(wclk), .Q(ram[8976]) );
  DFF ram_reg_929__7_ ( .D(n13192), .CP(wclk), .Q(ram[8951]) );
  DFF ram_reg_929__6_ ( .D(n13191), .CP(wclk), .Q(ram[8950]) );
  DFF ram_reg_929__5_ ( .D(n13190), .CP(wclk), .Q(ram[8949]) );
  DFF ram_reg_929__4_ ( .D(n13189), .CP(wclk), .Q(ram[8948]) );
  DFF ram_reg_929__3_ ( .D(n13188), .CP(wclk), .Q(ram[8947]) );
  DFF ram_reg_929__2_ ( .D(n13187), .CP(wclk), .Q(ram[8946]) );
  DFF ram_reg_929__1_ ( .D(n13186), .CP(wclk), .Q(ram[8945]) );
  DFF ram_reg_929__0_ ( .D(n13185), .CP(wclk), .Q(ram[8944]) );
  DFF ram_reg_933__7_ ( .D(n13160), .CP(wclk), .Q(ram[8919]) );
  DFF ram_reg_933__6_ ( .D(n13159), .CP(wclk), .Q(ram[8918]) );
  DFF ram_reg_933__5_ ( .D(n13158), .CP(wclk), .Q(ram[8917]) );
  DFF ram_reg_933__4_ ( .D(n13157), .CP(wclk), .Q(ram[8916]) );
  DFF ram_reg_933__3_ ( .D(n13156), .CP(wclk), .Q(ram[8915]) );
  DFF ram_reg_933__2_ ( .D(n13155), .CP(wclk), .Q(ram[8914]) );
  DFF ram_reg_933__1_ ( .D(n13154), .CP(wclk), .Q(ram[8913]) );
  DFF ram_reg_933__0_ ( .D(n13153), .CP(wclk), .Q(ram[8912]) );
  DFF ram_reg_937__7_ ( .D(n13128), .CP(wclk), .Q(ram[8887]) );
  DFF ram_reg_937__6_ ( .D(n13127), .CP(wclk), .Q(ram[8886]) );
  DFF ram_reg_937__5_ ( .D(n13126), .CP(wclk), .Q(ram[8885]) );
  DFF ram_reg_937__4_ ( .D(n13125), .CP(wclk), .Q(ram[8884]) );
  DFF ram_reg_937__3_ ( .D(n13124), .CP(wclk), .Q(ram[8883]) );
  DFF ram_reg_937__2_ ( .D(n13123), .CP(wclk), .Q(ram[8882]) );
  DFF ram_reg_937__1_ ( .D(n13122), .CP(wclk), .Q(ram[8881]) );
  DFF ram_reg_937__0_ ( .D(n13121), .CP(wclk), .Q(ram[8880]) );
  DFF ram_reg_941__7_ ( .D(n13096), .CP(wclk), .Q(ram[8855]) );
  DFF ram_reg_941__6_ ( .D(n13095), .CP(wclk), .Q(ram[8854]) );
  DFF ram_reg_941__5_ ( .D(n13094), .CP(wclk), .Q(ram[8853]) );
  DFF ram_reg_941__4_ ( .D(n13093), .CP(wclk), .Q(ram[8852]) );
  DFF ram_reg_941__3_ ( .D(n13092), .CP(wclk), .Q(ram[8851]) );
  DFF ram_reg_941__2_ ( .D(n13091), .CP(wclk), .Q(ram[8850]) );
  DFF ram_reg_941__1_ ( .D(n13090), .CP(wclk), .Q(ram[8849]) );
  DFF ram_reg_941__0_ ( .D(n13089), .CP(wclk), .Q(ram[8848]) );
  DFF ram_reg_945__7_ ( .D(n13064), .CP(wclk), .Q(ram[8823]) );
  DFF ram_reg_945__6_ ( .D(n13063), .CP(wclk), .Q(ram[8822]) );
  DFF ram_reg_945__5_ ( .D(n13062), .CP(wclk), .Q(ram[8821]) );
  DFF ram_reg_945__4_ ( .D(n13061), .CP(wclk), .Q(ram[8820]) );
  DFF ram_reg_945__3_ ( .D(n13060), .CP(wclk), .Q(ram[8819]) );
  DFF ram_reg_945__2_ ( .D(n13059), .CP(wclk), .Q(ram[8818]) );
  DFF ram_reg_945__1_ ( .D(n13058), .CP(wclk), .Q(ram[8817]) );
  DFF ram_reg_945__0_ ( .D(n13057), .CP(wclk), .Q(ram[8816]) );
  DFF ram_reg_949__7_ ( .D(n13032), .CP(wclk), .Q(ram[8791]) );
  DFF ram_reg_949__6_ ( .D(n13031), .CP(wclk), .Q(ram[8790]) );
  DFF ram_reg_949__5_ ( .D(n13030), .CP(wclk), .Q(ram[8789]) );
  DFF ram_reg_949__4_ ( .D(n13029), .CP(wclk), .Q(ram[8788]) );
  DFF ram_reg_949__3_ ( .D(n13028), .CP(wclk), .Q(ram[8787]) );
  DFF ram_reg_949__2_ ( .D(n13027), .CP(wclk), .Q(ram[8786]) );
  DFF ram_reg_949__1_ ( .D(n13026), .CP(wclk), .Q(ram[8785]) );
  DFF ram_reg_949__0_ ( .D(n13025), .CP(wclk), .Q(ram[8784]) );
  DFF ram_reg_953__7_ ( .D(n13000), .CP(wclk), .Q(ram[8759]) );
  DFF ram_reg_953__6_ ( .D(n12999), .CP(wclk), .Q(ram[8758]) );
  DFF ram_reg_953__5_ ( .D(n12998), .CP(wclk), .Q(ram[8757]) );
  DFF ram_reg_953__4_ ( .D(n12997), .CP(wclk), .Q(ram[8756]) );
  DFF ram_reg_953__3_ ( .D(n12996), .CP(wclk), .Q(ram[8755]) );
  DFF ram_reg_953__2_ ( .D(n12995), .CP(wclk), .Q(ram[8754]) );
  DFF ram_reg_953__1_ ( .D(n12994), .CP(wclk), .Q(ram[8753]) );
  DFF ram_reg_953__0_ ( .D(n12993), .CP(wclk), .Q(ram[8752]) );
  DFF ram_reg_957__7_ ( .D(n12968), .CP(wclk), .Q(ram[8727]) );
  DFF ram_reg_957__6_ ( .D(n12967), .CP(wclk), .Q(ram[8726]) );
  DFF ram_reg_957__5_ ( .D(n12966), .CP(wclk), .Q(ram[8725]) );
  DFF ram_reg_957__4_ ( .D(n12965), .CP(wclk), .Q(ram[8724]) );
  DFF ram_reg_957__3_ ( .D(n12964), .CP(wclk), .Q(ram[8723]) );
  DFF ram_reg_957__2_ ( .D(n12963), .CP(wclk), .Q(ram[8722]) );
  DFF ram_reg_957__1_ ( .D(n12962), .CP(wclk), .Q(ram[8721]) );
  DFF ram_reg_957__0_ ( .D(n12961), .CP(wclk), .Q(ram[8720]) );
  DFF ram_reg_961__7_ ( .D(n12936), .CP(wclk), .Q(ram[8695]) );
  DFF ram_reg_961__6_ ( .D(n12935), .CP(wclk), .Q(ram[8694]) );
  DFF ram_reg_961__5_ ( .D(n12934), .CP(wclk), .Q(ram[8693]) );
  DFF ram_reg_961__4_ ( .D(n12933), .CP(wclk), .Q(ram[8692]) );
  DFF ram_reg_961__3_ ( .D(n12932), .CP(wclk), .Q(ram[8691]) );
  DFF ram_reg_961__2_ ( .D(n12931), .CP(wclk), .Q(ram[8690]) );
  DFF ram_reg_961__1_ ( .D(n12930), .CP(wclk), .Q(ram[8689]) );
  DFF ram_reg_961__0_ ( .D(n12929), .CP(wclk), .Q(ram[8688]) );
  DFF ram_reg_969__7_ ( .D(n12872), .CP(wclk), .Q(ram[8631]) );
  DFF ram_reg_969__6_ ( .D(n12871), .CP(wclk), .Q(ram[8630]) );
  DFF ram_reg_969__5_ ( .D(n12870), .CP(wclk), .Q(ram[8629]) );
  DFF ram_reg_969__4_ ( .D(n12869), .CP(wclk), .Q(ram[8628]) );
  DFF ram_reg_969__3_ ( .D(n12868), .CP(wclk), .Q(ram[8627]) );
  DFF ram_reg_969__2_ ( .D(n12867), .CP(wclk), .Q(ram[8626]) );
  DFF ram_reg_969__1_ ( .D(n12866), .CP(wclk), .Q(ram[8625]) );
  DFF ram_reg_969__0_ ( .D(n12865), .CP(wclk), .Q(ram[8624]) );
  DFF ram_reg_973__7_ ( .D(n12840), .CP(wclk), .Q(ram[8599]) );
  DFF ram_reg_973__6_ ( .D(n12839), .CP(wclk), .Q(ram[8598]) );
  DFF ram_reg_973__5_ ( .D(n12838), .CP(wclk), .Q(ram[8597]) );
  DFF ram_reg_973__4_ ( .D(n12837), .CP(wclk), .Q(ram[8596]) );
  DFF ram_reg_973__3_ ( .D(n12836), .CP(wclk), .Q(ram[8595]) );
  DFF ram_reg_973__2_ ( .D(n12835), .CP(wclk), .Q(ram[8594]) );
  DFF ram_reg_973__1_ ( .D(n12834), .CP(wclk), .Q(ram[8593]) );
  DFF ram_reg_973__0_ ( .D(n12833), .CP(wclk), .Q(ram[8592]) );
  DFF ram_reg_977__7_ ( .D(n12808), .CP(wclk), .Q(ram[8567]) );
  DFF ram_reg_977__6_ ( .D(n12807), .CP(wclk), .Q(ram[8566]) );
  DFF ram_reg_977__5_ ( .D(n12806), .CP(wclk), .Q(ram[8565]) );
  DFF ram_reg_977__4_ ( .D(n12805), .CP(wclk), .Q(ram[8564]) );
  DFF ram_reg_977__3_ ( .D(n12804), .CP(wclk), .Q(ram[8563]) );
  DFF ram_reg_977__2_ ( .D(n12803), .CP(wclk), .Q(ram[8562]) );
  DFF ram_reg_977__1_ ( .D(n12802), .CP(wclk), .Q(ram[8561]) );
  DFF ram_reg_977__0_ ( .D(n12801), .CP(wclk), .Q(ram[8560]) );
  DFF ram_reg_985__7_ ( .D(n12744), .CP(wclk), .Q(ram[8503]) );
  DFF ram_reg_985__6_ ( .D(n12743), .CP(wclk), .Q(ram[8502]) );
  DFF ram_reg_985__5_ ( .D(n12742), .CP(wclk), .Q(ram[8501]) );
  DFF ram_reg_985__4_ ( .D(n12741), .CP(wclk), .Q(ram[8500]) );
  DFF ram_reg_985__3_ ( .D(n12740), .CP(wclk), .Q(ram[8499]) );
  DFF ram_reg_985__2_ ( .D(n12739), .CP(wclk), .Q(ram[8498]) );
  DFF ram_reg_985__1_ ( .D(n12738), .CP(wclk), .Q(ram[8497]) );
  DFF ram_reg_985__0_ ( .D(n12737), .CP(wclk), .Q(ram[8496]) );
  DFF ram_reg_989__7_ ( .D(n12712), .CP(wclk), .Q(ram[8471]) );
  DFF ram_reg_989__6_ ( .D(n12711), .CP(wclk), .Q(ram[8470]) );
  DFF ram_reg_989__5_ ( .D(n12710), .CP(wclk), .Q(ram[8469]) );
  DFF ram_reg_989__4_ ( .D(n12709), .CP(wclk), .Q(ram[8468]) );
  DFF ram_reg_989__3_ ( .D(n12708), .CP(wclk), .Q(ram[8467]) );
  DFF ram_reg_989__2_ ( .D(n12707), .CP(wclk), .Q(ram[8466]) );
  DFF ram_reg_989__1_ ( .D(n12706), .CP(wclk), .Q(ram[8465]) );
  DFF ram_reg_989__0_ ( .D(n12705), .CP(wclk), .Q(ram[8464]) );
  DFF ram_reg_993__7_ ( .D(n12680), .CP(wclk), .Q(ram[8439]) );
  DFF ram_reg_993__6_ ( .D(n12679), .CP(wclk), .Q(ram[8438]) );
  DFF ram_reg_993__5_ ( .D(n12678), .CP(wclk), .Q(ram[8437]) );
  DFF ram_reg_993__4_ ( .D(n12677), .CP(wclk), .Q(ram[8436]) );
  DFF ram_reg_993__3_ ( .D(n12676), .CP(wclk), .Q(ram[8435]) );
  DFF ram_reg_993__2_ ( .D(n12675), .CP(wclk), .Q(ram[8434]) );
  DFF ram_reg_993__1_ ( .D(n12674), .CP(wclk), .Q(ram[8433]) );
  DFF ram_reg_993__0_ ( .D(n12673), .CP(wclk), .Q(ram[8432]) );
  DFF ram_reg_997__7_ ( .D(n12648), .CP(wclk), .Q(ram[8407]) );
  DFF ram_reg_997__6_ ( .D(n12647), .CP(wclk), .Q(ram[8406]) );
  DFF ram_reg_997__5_ ( .D(n12646), .CP(wclk), .Q(ram[8405]) );
  DFF ram_reg_997__4_ ( .D(n12645), .CP(wclk), .Q(ram[8404]) );
  DFF ram_reg_997__3_ ( .D(n12644), .CP(wclk), .Q(ram[8403]) );
  DFF ram_reg_997__2_ ( .D(n12643), .CP(wclk), .Q(ram[8402]) );
  DFF ram_reg_997__1_ ( .D(n12642), .CP(wclk), .Q(ram[8401]) );
  DFF ram_reg_997__0_ ( .D(n12641), .CP(wclk), .Q(ram[8400]) );
  DFF ram_reg_1001__7_ ( .D(n12616), .CP(wclk), .Q(ram[8375]) );
  DFF ram_reg_1001__6_ ( .D(n12615), .CP(wclk), .Q(ram[8374]) );
  DFF ram_reg_1001__5_ ( .D(n12614), .CP(wclk), .Q(ram[8373]) );
  DFF ram_reg_1001__4_ ( .D(n12613), .CP(wclk), .Q(ram[8372]) );
  DFF ram_reg_1001__3_ ( .D(n12612), .CP(wclk), .Q(ram[8371]) );
  DFF ram_reg_1001__2_ ( .D(n12611), .CP(wclk), .Q(ram[8370]) );
  DFF ram_reg_1001__1_ ( .D(n12610), .CP(wclk), .Q(ram[8369]) );
  DFF ram_reg_1001__0_ ( .D(n12609), .CP(wclk), .Q(ram[8368]) );
  DFF ram_reg_1005__7_ ( .D(n12584), .CP(wclk), .Q(ram[8343]) );
  DFF ram_reg_1005__6_ ( .D(n12583), .CP(wclk), .Q(ram[8342]) );
  DFF ram_reg_1005__5_ ( .D(n12582), .CP(wclk), .Q(ram[8341]) );
  DFF ram_reg_1005__4_ ( .D(n12581), .CP(wclk), .Q(ram[8340]) );
  DFF ram_reg_1005__3_ ( .D(n12580), .CP(wclk), .Q(ram[8339]) );
  DFF ram_reg_1005__2_ ( .D(n12579), .CP(wclk), .Q(ram[8338]) );
  DFF ram_reg_1005__1_ ( .D(n12578), .CP(wclk), .Q(ram[8337]) );
  DFF ram_reg_1005__0_ ( .D(n12577), .CP(wclk), .Q(ram[8336]) );
  DFF ram_reg_1009__7_ ( .D(n12552), .CP(wclk), .Q(ram[8311]) );
  DFF ram_reg_1009__6_ ( .D(n12551), .CP(wclk), .Q(ram[8310]) );
  DFF ram_reg_1009__5_ ( .D(n12550), .CP(wclk), .Q(ram[8309]) );
  DFF ram_reg_1009__4_ ( .D(n12549), .CP(wclk), .Q(ram[8308]) );
  DFF ram_reg_1009__3_ ( .D(n12548), .CP(wclk), .Q(ram[8307]) );
  DFF ram_reg_1009__2_ ( .D(n12547), .CP(wclk), .Q(ram[8306]) );
  DFF ram_reg_1009__1_ ( .D(n12546), .CP(wclk), .Q(ram[8305]) );
  DFF ram_reg_1009__0_ ( .D(n12545), .CP(wclk), .Q(ram[8304]) );
  DFF ram_reg_1013__7_ ( .D(n12520), .CP(wclk), .Q(ram[8279]) );
  DFF ram_reg_1013__6_ ( .D(n12519), .CP(wclk), .Q(ram[8278]) );
  DFF ram_reg_1013__5_ ( .D(n12518), .CP(wclk), .Q(ram[8277]) );
  DFF ram_reg_1013__4_ ( .D(n12517), .CP(wclk), .Q(ram[8276]) );
  DFF ram_reg_1013__3_ ( .D(n12516), .CP(wclk), .Q(ram[8275]) );
  DFF ram_reg_1013__2_ ( .D(n12515), .CP(wclk), .Q(ram[8274]) );
  DFF ram_reg_1013__1_ ( .D(n12514), .CP(wclk), .Q(ram[8273]) );
  DFF ram_reg_1013__0_ ( .D(n12513), .CP(wclk), .Q(ram[8272]) );
  DFF ram_reg_1017__7_ ( .D(n12488), .CP(wclk), .Q(ram[8247]) );
  DFF ram_reg_1017__6_ ( .D(n12487), .CP(wclk), .Q(ram[8246]) );
  DFF ram_reg_1017__5_ ( .D(n12486), .CP(wclk), .Q(ram[8245]) );
  DFF ram_reg_1017__4_ ( .D(n12485), .CP(wclk), .Q(ram[8244]) );
  DFF ram_reg_1017__3_ ( .D(n12484), .CP(wclk), .Q(ram[8243]) );
  DFF ram_reg_1017__2_ ( .D(n12483), .CP(wclk), .Q(ram[8242]) );
  DFF ram_reg_1017__1_ ( .D(n12482), .CP(wclk), .Q(ram[8241]) );
  DFF ram_reg_1017__0_ ( .D(n12481), .CP(wclk), .Q(ram[8240]) );
  DFF ram_reg_1021__7_ ( .D(n12456), .CP(wclk), .Q(ram[8215]) );
  DFF ram_reg_1021__6_ ( .D(n12455), .CP(wclk), .Q(ram[8214]) );
  DFF ram_reg_1021__5_ ( .D(n12454), .CP(wclk), .Q(ram[8213]) );
  DFF ram_reg_1021__4_ ( .D(n12453), .CP(wclk), .Q(ram[8212]) );
  DFF ram_reg_1021__3_ ( .D(n12452), .CP(wclk), .Q(ram[8211]) );
  DFF ram_reg_1021__2_ ( .D(n12451), .CP(wclk), .Q(ram[8210]) );
  DFF ram_reg_1021__1_ ( .D(n12450), .CP(wclk), .Q(ram[8209]) );
  DFF ram_reg_1021__0_ ( .D(n12449), .CP(wclk), .Q(ram[8208]) );
  DFF ram_reg_1033__7_ ( .D(n12360), .CP(wclk), .Q(ram[8119]) );
  DFF ram_reg_1033__6_ ( .D(n12359), .CP(wclk), .Q(ram[8118]) );
  DFF ram_reg_1033__5_ ( .D(n12358), .CP(wclk), .Q(ram[8117]) );
  DFF ram_reg_1033__4_ ( .D(n12357), .CP(wclk), .Q(ram[8116]) );
  DFF ram_reg_1033__3_ ( .D(n12356), .CP(wclk), .Q(ram[8115]) );
  DFF ram_reg_1033__2_ ( .D(n12355), .CP(wclk), .Q(ram[8114]) );
  DFF ram_reg_1033__1_ ( .D(n12354), .CP(wclk), .Q(ram[8113]) );
  DFF ram_reg_1033__0_ ( .D(n12353), .CP(wclk), .Q(ram[8112]) );
  DFF ram_reg_1037__7_ ( .D(n12328), .CP(wclk), .Q(ram[8087]) );
  DFF ram_reg_1037__6_ ( .D(n12327), .CP(wclk), .Q(ram[8086]) );
  DFF ram_reg_1037__5_ ( .D(n12326), .CP(wclk), .Q(ram[8085]) );
  DFF ram_reg_1037__4_ ( .D(n12325), .CP(wclk), .Q(ram[8084]) );
  DFF ram_reg_1037__3_ ( .D(n12324), .CP(wclk), .Q(ram[8083]) );
  DFF ram_reg_1037__2_ ( .D(n12323), .CP(wclk), .Q(ram[8082]) );
  DFF ram_reg_1037__1_ ( .D(n12322), .CP(wclk), .Q(ram[8081]) );
  DFF ram_reg_1037__0_ ( .D(n12321), .CP(wclk), .Q(ram[8080]) );
  DFF ram_reg_1049__7_ ( .D(n12232), .CP(wclk), .Q(ram[7991]) );
  DFF ram_reg_1049__6_ ( .D(n12231), .CP(wclk), .Q(ram[7990]) );
  DFF ram_reg_1049__5_ ( .D(n12230), .CP(wclk), .Q(ram[7989]) );
  DFF ram_reg_1049__4_ ( .D(n12229), .CP(wclk), .Q(ram[7988]) );
  DFF ram_reg_1049__3_ ( .D(n12228), .CP(wclk), .Q(ram[7987]) );
  DFF ram_reg_1049__2_ ( .D(n12227), .CP(wclk), .Q(ram[7986]) );
  DFF ram_reg_1049__1_ ( .D(n12226), .CP(wclk), .Q(ram[7985]) );
  DFF ram_reg_1049__0_ ( .D(n12225), .CP(wclk), .Q(ram[7984]) );
  DFF ram_reg_1065__7_ ( .D(n12104), .CP(wclk), .Q(ram[7863]) );
  DFF ram_reg_1065__6_ ( .D(n12103), .CP(wclk), .Q(ram[7862]) );
  DFF ram_reg_1065__5_ ( .D(n12102), .CP(wclk), .Q(ram[7861]) );
  DFF ram_reg_1065__4_ ( .D(n12101), .CP(wclk), .Q(ram[7860]) );
  DFF ram_reg_1065__3_ ( .D(n12100), .CP(wclk), .Q(ram[7859]) );
  DFF ram_reg_1065__2_ ( .D(n12099), .CP(wclk), .Q(ram[7858]) );
  DFF ram_reg_1065__1_ ( .D(n12098), .CP(wclk), .Q(ram[7857]) );
  DFF ram_reg_1065__0_ ( .D(n12097), .CP(wclk), .Q(ram[7856]) );
  DFF ram_reg_1069__7_ ( .D(n12072), .CP(wclk), .Q(ram[7831]) );
  DFF ram_reg_1069__6_ ( .D(n12071), .CP(wclk), .Q(ram[7830]) );
  DFF ram_reg_1069__5_ ( .D(n12070), .CP(wclk), .Q(ram[7829]) );
  DFF ram_reg_1069__4_ ( .D(n12069), .CP(wclk), .Q(ram[7828]) );
  DFF ram_reg_1069__3_ ( .D(n12068), .CP(wclk), .Q(ram[7827]) );
  DFF ram_reg_1069__2_ ( .D(n12067), .CP(wclk), .Q(ram[7826]) );
  DFF ram_reg_1069__1_ ( .D(n12066), .CP(wclk), .Q(ram[7825]) );
  DFF ram_reg_1069__0_ ( .D(n12065), .CP(wclk), .Q(ram[7824]) );
  DFF ram_reg_1073__7_ ( .D(n12040), .CP(wclk), .Q(ram[7799]) );
  DFF ram_reg_1073__6_ ( .D(n12039), .CP(wclk), .Q(ram[7798]) );
  DFF ram_reg_1073__5_ ( .D(n12038), .CP(wclk), .Q(ram[7797]) );
  DFF ram_reg_1073__4_ ( .D(n12037), .CP(wclk), .Q(ram[7796]) );
  DFF ram_reg_1073__3_ ( .D(n12036), .CP(wclk), .Q(ram[7795]) );
  DFF ram_reg_1073__2_ ( .D(n12035), .CP(wclk), .Q(ram[7794]) );
  DFF ram_reg_1073__1_ ( .D(n12034), .CP(wclk), .Q(ram[7793]) );
  DFF ram_reg_1073__0_ ( .D(n12033), .CP(wclk), .Q(ram[7792]) );
  DFF ram_reg_1081__7_ ( .D(n11976), .CP(wclk), .Q(ram[7735]) );
  DFF ram_reg_1081__6_ ( .D(n11975), .CP(wclk), .Q(ram[7734]) );
  DFF ram_reg_1081__5_ ( .D(n11974), .CP(wclk), .Q(ram[7733]) );
  DFF ram_reg_1081__4_ ( .D(n11973), .CP(wclk), .Q(ram[7732]) );
  DFF ram_reg_1081__3_ ( .D(n11972), .CP(wclk), .Q(ram[7731]) );
  DFF ram_reg_1081__2_ ( .D(n11971), .CP(wclk), .Q(ram[7730]) );
  DFF ram_reg_1081__1_ ( .D(n11970), .CP(wclk), .Q(ram[7729]) );
  DFF ram_reg_1081__0_ ( .D(n11969), .CP(wclk), .Q(ram[7728]) );
  DFF ram_reg_1085__7_ ( .D(n11944), .CP(wclk), .Q(ram[7703]) );
  DFF ram_reg_1085__6_ ( .D(n11943), .CP(wclk), .Q(ram[7702]) );
  DFF ram_reg_1085__5_ ( .D(n11942), .CP(wclk), .Q(ram[7701]) );
  DFF ram_reg_1085__4_ ( .D(n11941), .CP(wclk), .Q(ram[7700]) );
  DFF ram_reg_1085__3_ ( .D(n11940), .CP(wclk), .Q(ram[7699]) );
  DFF ram_reg_1085__2_ ( .D(n11939), .CP(wclk), .Q(ram[7698]) );
  DFF ram_reg_1085__1_ ( .D(n11938), .CP(wclk), .Q(ram[7697]) );
  DFF ram_reg_1085__0_ ( .D(n11937), .CP(wclk), .Q(ram[7696]) );
  DFF ram_reg_1129__7_ ( .D(n11592), .CP(wclk), .Q(ram[7351]) );
  DFF ram_reg_1129__6_ ( .D(n11591), .CP(wclk), .Q(ram[7350]) );
  DFF ram_reg_1129__5_ ( .D(n11590), .CP(wclk), .Q(ram[7349]) );
  DFF ram_reg_1129__4_ ( .D(n11589), .CP(wclk), .Q(ram[7348]) );
  DFF ram_reg_1129__3_ ( .D(n11588), .CP(wclk), .Q(ram[7347]) );
  DFF ram_reg_1129__2_ ( .D(n11587), .CP(wclk), .Q(ram[7346]) );
  DFF ram_reg_1129__1_ ( .D(n11586), .CP(wclk), .Q(ram[7345]) );
  DFF ram_reg_1129__0_ ( .D(n11585), .CP(wclk), .Q(ram[7344]) );
  DFF ram_reg_1145__7_ ( .D(n11464), .CP(wclk), .Q(ram[7223]) );
  DFF ram_reg_1145__6_ ( .D(n11463), .CP(wclk), .Q(ram[7222]) );
  DFF ram_reg_1145__5_ ( .D(n11462), .CP(wclk), .Q(ram[7221]) );
  DFF ram_reg_1145__4_ ( .D(n11461), .CP(wclk), .Q(ram[7220]) );
  DFF ram_reg_1145__3_ ( .D(n11460), .CP(wclk), .Q(ram[7219]) );
  DFF ram_reg_1145__2_ ( .D(n11459), .CP(wclk), .Q(ram[7218]) );
  DFF ram_reg_1145__1_ ( .D(n11458), .CP(wclk), .Q(ram[7217]) );
  DFF ram_reg_1145__0_ ( .D(n11457), .CP(wclk), .Q(ram[7216]) );
  DFF ram_reg_1153__7_ ( .D(n11400), .CP(wclk), .Q(ram[7159]) );
  DFF ram_reg_1153__6_ ( .D(n11399), .CP(wclk), .Q(ram[7158]) );
  DFF ram_reg_1153__5_ ( .D(n11398), .CP(wclk), .Q(ram[7157]) );
  DFF ram_reg_1153__4_ ( .D(n11397), .CP(wclk), .Q(ram[7156]) );
  DFF ram_reg_1153__3_ ( .D(n11396), .CP(wclk), .Q(ram[7155]) );
  DFF ram_reg_1153__2_ ( .D(n11395), .CP(wclk), .Q(ram[7154]) );
  DFF ram_reg_1153__1_ ( .D(n11394), .CP(wclk), .Q(ram[7153]) );
  DFF ram_reg_1153__0_ ( .D(n11393), .CP(wclk), .Q(ram[7152]) );
  DFF ram_reg_1161__7_ ( .D(n11336), .CP(wclk), .Q(ram[7095]) );
  DFF ram_reg_1161__6_ ( .D(n11335), .CP(wclk), .Q(ram[7094]) );
  DFF ram_reg_1161__5_ ( .D(n11334), .CP(wclk), .Q(ram[7093]) );
  DFF ram_reg_1161__4_ ( .D(n11333), .CP(wclk), .Q(ram[7092]) );
  DFF ram_reg_1161__3_ ( .D(n11332), .CP(wclk), .Q(ram[7091]) );
  DFF ram_reg_1161__2_ ( .D(n11331), .CP(wclk), .Q(ram[7090]) );
  DFF ram_reg_1161__1_ ( .D(n11330), .CP(wclk), .Q(ram[7089]) );
  DFF ram_reg_1161__0_ ( .D(n11329), .CP(wclk), .Q(ram[7088]) );
  DFF ram_reg_1165__7_ ( .D(n11304), .CP(wclk), .Q(ram[7063]) );
  DFF ram_reg_1165__6_ ( .D(n11303), .CP(wclk), .Q(ram[7062]) );
  DFF ram_reg_1165__5_ ( .D(n11302), .CP(wclk), .Q(ram[7061]) );
  DFF ram_reg_1165__4_ ( .D(n11301), .CP(wclk), .Q(ram[7060]) );
  DFF ram_reg_1165__3_ ( .D(n11300), .CP(wclk), .Q(ram[7059]) );
  DFF ram_reg_1165__2_ ( .D(n11299), .CP(wclk), .Q(ram[7058]) );
  DFF ram_reg_1165__1_ ( .D(n11298), .CP(wclk), .Q(ram[7057]) );
  DFF ram_reg_1165__0_ ( .D(n11297), .CP(wclk), .Q(ram[7056]) );
  DFF ram_reg_1169__7_ ( .D(n11272), .CP(wclk), .Q(ram[7031]) );
  DFF ram_reg_1169__6_ ( .D(n11271), .CP(wclk), .Q(ram[7030]) );
  DFF ram_reg_1169__5_ ( .D(n11270), .CP(wclk), .Q(ram[7029]) );
  DFF ram_reg_1169__4_ ( .D(n11269), .CP(wclk), .Q(ram[7028]) );
  DFF ram_reg_1169__3_ ( .D(n11268), .CP(wclk), .Q(ram[7027]) );
  DFF ram_reg_1169__2_ ( .D(n11267), .CP(wclk), .Q(ram[7026]) );
  DFF ram_reg_1169__1_ ( .D(n11266), .CP(wclk), .Q(ram[7025]) );
  DFF ram_reg_1169__0_ ( .D(n11265), .CP(wclk), .Q(ram[7024]) );
  DFF ram_reg_1177__7_ ( .D(n11208), .CP(wclk), .Q(ram[6967]) );
  DFF ram_reg_1177__6_ ( .D(n11207), .CP(wclk), .Q(ram[6966]) );
  DFF ram_reg_1177__5_ ( .D(n11206), .CP(wclk), .Q(ram[6965]) );
  DFF ram_reg_1177__4_ ( .D(n11205), .CP(wclk), .Q(ram[6964]) );
  DFF ram_reg_1177__3_ ( .D(n11204), .CP(wclk), .Q(ram[6963]) );
  DFF ram_reg_1177__2_ ( .D(n11203), .CP(wclk), .Q(ram[6962]) );
  DFF ram_reg_1177__1_ ( .D(n11202), .CP(wclk), .Q(ram[6961]) );
  DFF ram_reg_1177__0_ ( .D(n11201), .CP(wclk), .Q(ram[6960]) );
  DFF ram_reg_1181__7_ ( .D(n11176), .CP(wclk), .Q(ram[6935]) );
  DFF ram_reg_1181__6_ ( .D(n11175), .CP(wclk), .Q(ram[6934]) );
  DFF ram_reg_1181__5_ ( .D(n11174), .CP(wclk), .Q(ram[6933]) );
  DFF ram_reg_1181__4_ ( .D(n11173), .CP(wclk), .Q(ram[6932]) );
  DFF ram_reg_1181__3_ ( .D(n11172), .CP(wclk), .Q(ram[6931]) );
  DFF ram_reg_1181__2_ ( .D(n11171), .CP(wclk), .Q(ram[6930]) );
  DFF ram_reg_1181__1_ ( .D(n11170), .CP(wclk), .Q(ram[6929]) );
  DFF ram_reg_1181__0_ ( .D(n11169), .CP(wclk), .Q(ram[6928]) );
  DFF ram_reg_1185__7_ ( .D(n11144), .CP(wclk), .Q(ram[6903]) );
  DFF ram_reg_1185__6_ ( .D(n11143), .CP(wclk), .Q(ram[6902]) );
  DFF ram_reg_1185__5_ ( .D(n11142), .CP(wclk), .Q(ram[6901]) );
  DFF ram_reg_1185__4_ ( .D(n11141), .CP(wclk), .Q(ram[6900]) );
  DFF ram_reg_1185__3_ ( .D(n11140), .CP(wclk), .Q(ram[6899]) );
  DFF ram_reg_1185__2_ ( .D(n11139), .CP(wclk), .Q(ram[6898]) );
  DFF ram_reg_1185__1_ ( .D(n11138), .CP(wclk), .Q(ram[6897]) );
  DFF ram_reg_1185__0_ ( .D(n11137), .CP(wclk), .Q(ram[6896]) );
  DFF ram_reg_1189__7_ ( .D(n11112), .CP(wclk), .Q(ram[6871]) );
  DFF ram_reg_1189__6_ ( .D(n11111), .CP(wclk), .Q(ram[6870]) );
  DFF ram_reg_1189__5_ ( .D(n11110), .CP(wclk), .Q(ram[6869]) );
  DFF ram_reg_1189__4_ ( .D(n11109), .CP(wclk), .Q(ram[6868]) );
  DFF ram_reg_1189__3_ ( .D(n11108), .CP(wclk), .Q(ram[6867]) );
  DFF ram_reg_1189__2_ ( .D(n11107), .CP(wclk), .Q(ram[6866]) );
  DFF ram_reg_1189__1_ ( .D(n11106), .CP(wclk), .Q(ram[6865]) );
  DFF ram_reg_1189__0_ ( .D(n11105), .CP(wclk), .Q(ram[6864]) );
  DFF ram_reg_1193__7_ ( .D(n11080), .CP(wclk), .Q(ram[6839]) );
  DFF ram_reg_1193__6_ ( .D(n11079), .CP(wclk), .Q(ram[6838]) );
  DFF ram_reg_1193__5_ ( .D(n11078), .CP(wclk), .Q(ram[6837]) );
  DFF ram_reg_1193__4_ ( .D(n11077), .CP(wclk), .Q(ram[6836]) );
  DFF ram_reg_1193__3_ ( .D(n11076), .CP(wclk), .Q(ram[6835]) );
  DFF ram_reg_1193__2_ ( .D(n11075), .CP(wclk), .Q(ram[6834]) );
  DFF ram_reg_1193__1_ ( .D(n11074), .CP(wclk), .Q(ram[6833]) );
  DFF ram_reg_1193__0_ ( .D(n11073), .CP(wclk), .Q(ram[6832]) );
  DFF ram_reg_1197__7_ ( .D(n11048), .CP(wclk), .Q(ram[6807]) );
  DFF ram_reg_1197__6_ ( .D(n11047), .CP(wclk), .Q(ram[6806]) );
  DFF ram_reg_1197__5_ ( .D(n11046), .CP(wclk), .Q(ram[6805]) );
  DFF ram_reg_1197__4_ ( .D(n11045), .CP(wclk), .Q(ram[6804]) );
  DFF ram_reg_1197__3_ ( .D(n11044), .CP(wclk), .Q(ram[6803]) );
  DFF ram_reg_1197__2_ ( .D(n11043), .CP(wclk), .Q(ram[6802]) );
  DFF ram_reg_1197__1_ ( .D(n11042), .CP(wclk), .Q(ram[6801]) );
  DFF ram_reg_1197__0_ ( .D(n11041), .CP(wclk), .Q(ram[6800]) );
  DFF ram_reg_1201__7_ ( .D(n11016), .CP(wclk), .Q(ram[6775]) );
  DFF ram_reg_1201__6_ ( .D(n11015), .CP(wclk), .Q(ram[6774]) );
  DFF ram_reg_1201__5_ ( .D(n11014), .CP(wclk), .Q(ram[6773]) );
  DFF ram_reg_1201__4_ ( .D(n11013), .CP(wclk), .Q(ram[6772]) );
  DFF ram_reg_1201__3_ ( .D(n11012), .CP(wclk), .Q(ram[6771]) );
  DFF ram_reg_1201__2_ ( .D(n11011), .CP(wclk), .Q(ram[6770]) );
  DFF ram_reg_1201__1_ ( .D(n11010), .CP(wclk), .Q(ram[6769]) );
  DFF ram_reg_1201__0_ ( .D(n11009), .CP(wclk), .Q(ram[6768]) );
  DFF ram_reg_1205__7_ ( .D(n10984), .CP(wclk), .Q(ram[6743]) );
  DFF ram_reg_1205__6_ ( .D(n10983), .CP(wclk), .Q(ram[6742]) );
  DFF ram_reg_1205__5_ ( .D(n10982), .CP(wclk), .Q(ram[6741]) );
  DFF ram_reg_1205__4_ ( .D(n10981), .CP(wclk), .Q(ram[6740]) );
  DFF ram_reg_1205__3_ ( .D(n10980), .CP(wclk), .Q(ram[6739]) );
  DFF ram_reg_1205__2_ ( .D(n10979), .CP(wclk), .Q(ram[6738]) );
  DFF ram_reg_1205__1_ ( .D(n10978), .CP(wclk), .Q(ram[6737]) );
  DFF ram_reg_1205__0_ ( .D(n10977), .CP(wclk), .Q(ram[6736]) );
  DFF ram_reg_1209__7_ ( .D(n10952), .CP(wclk), .Q(ram[6711]) );
  DFF ram_reg_1209__6_ ( .D(n10951), .CP(wclk), .Q(ram[6710]) );
  DFF ram_reg_1209__5_ ( .D(n10950), .CP(wclk), .Q(ram[6709]) );
  DFF ram_reg_1209__4_ ( .D(n10949), .CP(wclk), .Q(ram[6708]) );
  DFF ram_reg_1209__3_ ( .D(n10948), .CP(wclk), .Q(ram[6707]) );
  DFF ram_reg_1209__2_ ( .D(n10947), .CP(wclk), .Q(ram[6706]) );
  DFF ram_reg_1209__1_ ( .D(n10946), .CP(wclk), .Q(ram[6705]) );
  DFF ram_reg_1209__0_ ( .D(n10945), .CP(wclk), .Q(ram[6704]) );
  DFF ram_reg_1213__7_ ( .D(n10920), .CP(wclk), .Q(ram[6679]) );
  DFF ram_reg_1213__6_ ( .D(n10919), .CP(wclk), .Q(ram[6678]) );
  DFF ram_reg_1213__5_ ( .D(n10918), .CP(wclk), .Q(ram[6677]) );
  DFF ram_reg_1213__4_ ( .D(n10917), .CP(wclk), .Q(ram[6676]) );
  DFF ram_reg_1213__3_ ( .D(n10916), .CP(wclk), .Q(ram[6675]) );
  DFF ram_reg_1213__2_ ( .D(n10915), .CP(wclk), .Q(ram[6674]) );
  DFF ram_reg_1213__1_ ( .D(n10914), .CP(wclk), .Q(ram[6673]) );
  DFF ram_reg_1213__0_ ( .D(n10913), .CP(wclk), .Q(ram[6672]) );
  DFF ram_reg_1217__7_ ( .D(n10888), .CP(wclk), .Q(ram[6647]) );
  DFF ram_reg_1217__6_ ( .D(n10887), .CP(wclk), .Q(ram[6646]) );
  DFF ram_reg_1217__5_ ( .D(n10886), .CP(wclk), .Q(ram[6645]) );
  DFF ram_reg_1217__4_ ( .D(n10885), .CP(wclk), .Q(ram[6644]) );
  DFF ram_reg_1217__3_ ( .D(n10884), .CP(wclk), .Q(ram[6643]) );
  DFF ram_reg_1217__2_ ( .D(n10883), .CP(wclk), .Q(ram[6642]) );
  DFF ram_reg_1217__1_ ( .D(n10882), .CP(wclk), .Q(ram[6641]) );
  DFF ram_reg_1217__0_ ( .D(n10881), .CP(wclk), .Q(ram[6640]) );
  DFF ram_reg_1225__7_ ( .D(n10824), .CP(wclk), .Q(ram[6583]) );
  DFF ram_reg_1225__6_ ( .D(n10823), .CP(wclk), .Q(ram[6582]) );
  DFF ram_reg_1225__5_ ( .D(n10822), .CP(wclk), .Q(ram[6581]) );
  DFF ram_reg_1225__4_ ( .D(n10821), .CP(wclk), .Q(ram[6580]) );
  DFF ram_reg_1225__3_ ( .D(n10820), .CP(wclk), .Q(ram[6579]) );
  DFF ram_reg_1225__2_ ( .D(n10819), .CP(wclk), .Q(ram[6578]) );
  DFF ram_reg_1225__1_ ( .D(n10818), .CP(wclk), .Q(ram[6577]) );
  DFF ram_reg_1225__0_ ( .D(n10817), .CP(wclk), .Q(ram[6576]) );
  DFF ram_reg_1229__7_ ( .D(n10792), .CP(wclk), .Q(ram[6551]) );
  DFF ram_reg_1229__6_ ( .D(n10791), .CP(wclk), .Q(ram[6550]) );
  DFF ram_reg_1229__5_ ( .D(n10790), .CP(wclk), .Q(ram[6549]) );
  DFF ram_reg_1229__4_ ( .D(n10789), .CP(wclk), .Q(ram[6548]) );
  DFF ram_reg_1229__3_ ( .D(n10788), .CP(wclk), .Q(ram[6547]) );
  DFF ram_reg_1229__2_ ( .D(n10787), .CP(wclk), .Q(ram[6546]) );
  DFF ram_reg_1229__1_ ( .D(n10786), .CP(wclk), .Q(ram[6545]) );
  DFF ram_reg_1229__0_ ( .D(n10785), .CP(wclk), .Q(ram[6544]) );
  DFF ram_reg_1241__7_ ( .D(n10696), .CP(wclk), .Q(ram[6455]) );
  DFF ram_reg_1241__6_ ( .D(n10695), .CP(wclk), .Q(ram[6454]) );
  DFF ram_reg_1241__5_ ( .D(n10694), .CP(wclk), .Q(ram[6453]) );
  DFF ram_reg_1241__4_ ( .D(n10693), .CP(wclk), .Q(ram[6452]) );
  DFF ram_reg_1241__3_ ( .D(n10692), .CP(wclk), .Q(ram[6451]) );
  DFF ram_reg_1241__2_ ( .D(n10691), .CP(wclk), .Q(ram[6450]) );
  DFF ram_reg_1241__1_ ( .D(n10690), .CP(wclk), .Q(ram[6449]) );
  DFF ram_reg_1241__0_ ( .D(n10689), .CP(wclk), .Q(ram[6448]) );
  DFF ram_reg_1245__7_ ( .D(n10664), .CP(wclk), .Q(ram[6423]) );
  DFF ram_reg_1245__6_ ( .D(n10663), .CP(wclk), .Q(ram[6422]) );
  DFF ram_reg_1245__5_ ( .D(n10662), .CP(wclk), .Q(ram[6421]) );
  DFF ram_reg_1245__4_ ( .D(n10661), .CP(wclk), .Q(ram[6420]) );
  DFF ram_reg_1245__3_ ( .D(n10660), .CP(wclk), .Q(ram[6419]) );
  DFF ram_reg_1245__2_ ( .D(n10659), .CP(wclk), .Q(ram[6418]) );
  DFF ram_reg_1245__1_ ( .D(n10658), .CP(wclk), .Q(ram[6417]) );
  DFF ram_reg_1245__0_ ( .D(n10657), .CP(wclk), .Q(ram[6416]) );
  DFF ram_reg_1249__7_ ( .D(n10632), .CP(wclk), .Q(ram[6391]) );
  DFF ram_reg_1249__6_ ( .D(n10631), .CP(wclk), .Q(ram[6390]) );
  DFF ram_reg_1249__5_ ( .D(n10630), .CP(wclk), .Q(ram[6389]) );
  DFF ram_reg_1249__4_ ( .D(n10629), .CP(wclk), .Q(ram[6388]) );
  DFF ram_reg_1249__3_ ( .D(n10628), .CP(wclk), .Q(ram[6387]) );
  DFF ram_reg_1249__2_ ( .D(n10627), .CP(wclk), .Q(ram[6386]) );
  DFF ram_reg_1249__1_ ( .D(n10626), .CP(wclk), .Q(ram[6385]) );
  DFF ram_reg_1249__0_ ( .D(n10625), .CP(wclk), .Q(ram[6384]) );
  DFF ram_reg_1257__7_ ( .D(n10568), .CP(wclk), .Q(ram[6327]) );
  DFF ram_reg_1257__6_ ( .D(n10567), .CP(wclk), .Q(ram[6326]) );
  DFF ram_reg_1257__5_ ( .D(n10566), .CP(wclk), .Q(ram[6325]) );
  DFF ram_reg_1257__4_ ( .D(n10565), .CP(wclk), .Q(ram[6324]) );
  DFF ram_reg_1257__3_ ( .D(n10564), .CP(wclk), .Q(ram[6323]) );
  DFF ram_reg_1257__2_ ( .D(n10563), .CP(wclk), .Q(ram[6322]) );
  DFF ram_reg_1257__1_ ( .D(n10562), .CP(wclk), .Q(ram[6321]) );
  DFF ram_reg_1257__0_ ( .D(n10561), .CP(wclk), .Q(ram[6320]) );
  DFF ram_reg_1261__7_ ( .D(n10536), .CP(wclk), .Q(ram[6295]) );
  DFF ram_reg_1261__6_ ( .D(n10535), .CP(wclk), .Q(ram[6294]) );
  DFF ram_reg_1261__5_ ( .D(n10534), .CP(wclk), .Q(ram[6293]) );
  DFF ram_reg_1261__4_ ( .D(n10533), .CP(wclk), .Q(ram[6292]) );
  DFF ram_reg_1261__3_ ( .D(n10532), .CP(wclk), .Q(ram[6291]) );
  DFF ram_reg_1261__2_ ( .D(n10531), .CP(wclk), .Q(ram[6290]) );
  DFF ram_reg_1261__1_ ( .D(n10530), .CP(wclk), .Q(ram[6289]) );
  DFF ram_reg_1261__0_ ( .D(n10529), .CP(wclk), .Q(ram[6288]) );
  DFF ram_reg_1265__7_ ( .D(n10504), .CP(wclk), .Q(ram[6263]) );
  DFF ram_reg_1265__6_ ( .D(n10503), .CP(wclk), .Q(ram[6262]) );
  DFF ram_reg_1265__5_ ( .D(n10502), .CP(wclk), .Q(ram[6261]) );
  DFF ram_reg_1265__4_ ( .D(n10501), .CP(wclk), .Q(ram[6260]) );
  DFF ram_reg_1265__3_ ( .D(n10500), .CP(wclk), .Q(ram[6259]) );
  DFF ram_reg_1265__2_ ( .D(n10499), .CP(wclk), .Q(ram[6258]) );
  DFF ram_reg_1265__1_ ( .D(n10498), .CP(wclk), .Q(ram[6257]) );
  DFF ram_reg_1265__0_ ( .D(n10497), .CP(wclk), .Q(ram[6256]) );
  DFF ram_reg_1273__7_ ( .D(n10440), .CP(wclk), .Q(ram[6199]) );
  DFF ram_reg_1273__6_ ( .D(n10439), .CP(wclk), .Q(ram[6198]) );
  DFF ram_reg_1273__5_ ( .D(n10438), .CP(wclk), .Q(ram[6197]) );
  DFF ram_reg_1273__4_ ( .D(n10437), .CP(wclk), .Q(ram[6196]) );
  DFF ram_reg_1273__3_ ( .D(n10436), .CP(wclk), .Q(ram[6195]) );
  DFF ram_reg_1273__2_ ( .D(n10435), .CP(wclk), .Q(ram[6194]) );
  DFF ram_reg_1273__1_ ( .D(n10434), .CP(wclk), .Q(ram[6193]) );
  DFF ram_reg_1273__0_ ( .D(n10433), .CP(wclk), .Q(ram[6192]) );
  DFF ram_reg_1277__7_ ( .D(n10408), .CP(wclk), .Q(ram[6167]) );
  DFF ram_reg_1277__6_ ( .D(n10407), .CP(wclk), .Q(ram[6166]) );
  DFF ram_reg_1277__5_ ( .D(n10406), .CP(wclk), .Q(ram[6165]) );
  DFF ram_reg_1277__4_ ( .D(n10405), .CP(wclk), .Q(ram[6164]) );
  DFF ram_reg_1277__3_ ( .D(n10404), .CP(wclk), .Q(ram[6163]) );
  DFF ram_reg_1277__2_ ( .D(n10403), .CP(wclk), .Q(ram[6162]) );
  DFF ram_reg_1277__1_ ( .D(n10402), .CP(wclk), .Q(ram[6161]) );
  DFF ram_reg_1277__0_ ( .D(n10401), .CP(wclk), .Q(ram[6160]) );
  DFF ram_reg_1281__7_ ( .D(n10376), .CP(wclk), .Q(ram[6135]) );
  DFF ram_reg_1281__6_ ( .D(n10375), .CP(wclk), .Q(ram[6134]) );
  DFF ram_reg_1281__5_ ( .D(n10374), .CP(wclk), .Q(ram[6133]) );
  DFF ram_reg_1281__4_ ( .D(n10373), .CP(wclk), .Q(ram[6132]) );
  DFF ram_reg_1281__3_ ( .D(n10372), .CP(wclk), .Q(ram[6131]) );
  DFF ram_reg_1281__2_ ( .D(n10371), .CP(wclk), .Q(ram[6130]) );
  DFF ram_reg_1281__1_ ( .D(n10370), .CP(wclk), .Q(ram[6129]) );
  DFF ram_reg_1281__0_ ( .D(n10369), .CP(wclk), .Q(ram[6128]) );
  DFF ram_reg_1289__7_ ( .D(n10312), .CP(wclk), .Q(ram[6071]) );
  DFF ram_reg_1289__6_ ( .D(n10311), .CP(wclk), .Q(ram[6070]) );
  DFF ram_reg_1289__5_ ( .D(n10310), .CP(wclk), .Q(ram[6069]) );
  DFF ram_reg_1289__4_ ( .D(n10309), .CP(wclk), .Q(ram[6068]) );
  DFF ram_reg_1289__3_ ( .D(n10308), .CP(wclk), .Q(ram[6067]) );
  DFF ram_reg_1289__2_ ( .D(n10307), .CP(wclk), .Q(ram[6066]) );
  DFF ram_reg_1289__1_ ( .D(n10306), .CP(wclk), .Q(ram[6065]) );
  DFF ram_reg_1289__0_ ( .D(n10305), .CP(wclk), .Q(ram[6064]) );
  DFF ram_reg_1293__7_ ( .D(n10280), .CP(wclk), .Q(ram[6039]) );
  DFF ram_reg_1293__6_ ( .D(n10279), .CP(wclk), .Q(ram[6038]) );
  DFF ram_reg_1293__5_ ( .D(n10278), .CP(wclk), .Q(ram[6037]) );
  DFF ram_reg_1293__4_ ( .D(n10277), .CP(wclk), .Q(ram[6036]) );
  DFF ram_reg_1293__3_ ( .D(n10276), .CP(wclk), .Q(ram[6035]) );
  DFF ram_reg_1293__2_ ( .D(n10275), .CP(wclk), .Q(ram[6034]) );
  DFF ram_reg_1293__1_ ( .D(n10274), .CP(wclk), .Q(ram[6033]) );
  DFF ram_reg_1293__0_ ( .D(n10273), .CP(wclk), .Q(ram[6032]) );
  DFF ram_reg_1305__7_ ( .D(n10184), .CP(wclk), .Q(ram[5943]) );
  DFF ram_reg_1305__6_ ( .D(n10183), .CP(wclk), .Q(ram[5942]) );
  DFF ram_reg_1305__5_ ( .D(n10182), .CP(wclk), .Q(ram[5941]) );
  DFF ram_reg_1305__4_ ( .D(n10181), .CP(wclk), .Q(ram[5940]) );
  DFF ram_reg_1305__3_ ( .D(n10180), .CP(wclk), .Q(ram[5939]) );
  DFF ram_reg_1305__2_ ( .D(n10179), .CP(wclk), .Q(ram[5938]) );
  DFF ram_reg_1305__1_ ( .D(n10178), .CP(wclk), .Q(ram[5937]) );
  DFF ram_reg_1305__0_ ( .D(n10177), .CP(wclk), .Q(ram[5936]) );
  DFF ram_reg_1309__7_ ( .D(n10152), .CP(wclk), .Q(ram[5911]) );
  DFF ram_reg_1309__6_ ( .D(n10151), .CP(wclk), .Q(ram[5910]) );
  DFF ram_reg_1309__5_ ( .D(n10150), .CP(wclk), .Q(ram[5909]) );
  DFF ram_reg_1309__4_ ( .D(n10149), .CP(wclk), .Q(ram[5908]) );
  DFF ram_reg_1309__3_ ( .D(n10148), .CP(wclk), .Q(ram[5907]) );
  DFF ram_reg_1309__2_ ( .D(n10147), .CP(wclk), .Q(ram[5906]) );
  DFF ram_reg_1309__1_ ( .D(n10146), .CP(wclk), .Q(ram[5905]) );
  DFF ram_reg_1309__0_ ( .D(n10145), .CP(wclk), .Q(ram[5904]) );
  DFF ram_reg_1313__7_ ( .D(n10120), .CP(wclk), .Q(ram[5879]) );
  DFF ram_reg_1313__6_ ( .D(n10119), .CP(wclk), .Q(ram[5878]) );
  DFF ram_reg_1313__5_ ( .D(n10118), .CP(wclk), .Q(ram[5877]) );
  DFF ram_reg_1313__4_ ( .D(n10117), .CP(wclk), .Q(ram[5876]) );
  DFF ram_reg_1313__3_ ( .D(n10116), .CP(wclk), .Q(ram[5875]) );
  DFF ram_reg_1313__2_ ( .D(n10115), .CP(wclk), .Q(ram[5874]) );
  DFF ram_reg_1313__1_ ( .D(n10114), .CP(wclk), .Q(ram[5873]) );
  DFF ram_reg_1313__0_ ( .D(n10113), .CP(wclk), .Q(ram[5872]) );
  DFF ram_reg_1321__7_ ( .D(n10056), .CP(wclk), .Q(ram[5815]) );
  DFF ram_reg_1321__6_ ( .D(n10055), .CP(wclk), .Q(ram[5814]) );
  DFF ram_reg_1321__5_ ( .D(n10054), .CP(wclk), .Q(ram[5813]) );
  DFF ram_reg_1321__4_ ( .D(n10053), .CP(wclk), .Q(ram[5812]) );
  DFF ram_reg_1321__3_ ( .D(n10052), .CP(wclk), .Q(ram[5811]) );
  DFF ram_reg_1321__2_ ( .D(n10051), .CP(wclk), .Q(ram[5810]) );
  DFF ram_reg_1321__1_ ( .D(n10050), .CP(wclk), .Q(ram[5809]) );
  DFF ram_reg_1321__0_ ( .D(n10049), .CP(wclk), .Q(ram[5808]) );
  DFF ram_reg_1325__7_ ( .D(n10024), .CP(wclk), .Q(ram[5783]) );
  DFF ram_reg_1325__6_ ( .D(n10023), .CP(wclk), .Q(ram[5782]) );
  DFF ram_reg_1325__5_ ( .D(n10022), .CP(wclk), .Q(ram[5781]) );
  DFF ram_reg_1325__4_ ( .D(n10021), .CP(wclk), .Q(ram[5780]) );
  DFF ram_reg_1325__3_ ( .D(n10020), .CP(wclk), .Q(ram[5779]) );
  DFF ram_reg_1325__2_ ( .D(n10019), .CP(wclk), .Q(ram[5778]) );
  DFF ram_reg_1325__1_ ( .D(n10018), .CP(wclk), .Q(ram[5777]) );
  DFF ram_reg_1325__0_ ( .D(n10017), .CP(wclk), .Q(ram[5776]) );
  DFF ram_reg_1329__7_ ( .D(n9992), .CP(wclk), .Q(ram[5751]) );
  DFF ram_reg_1329__6_ ( .D(n9991), .CP(wclk), .Q(ram[5750]) );
  DFF ram_reg_1329__5_ ( .D(n9990), .CP(wclk), .Q(ram[5749]) );
  DFF ram_reg_1329__4_ ( .D(n9989), .CP(wclk), .Q(ram[5748]) );
  DFF ram_reg_1329__3_ ( .D(n9988), .CP(wclk), .Q(ram[5747]) );
  DFF ram_reg_1329__2_ ( .D(n9987), .CP(wclk), .Q(ram[5746]) );
  DFF ram_reg_1329__1_ ( .D(n9986), .CP(wclk), .Q(ram[5745]) );
  DFF ram_reg_1329__0_ ( .D(n9985), .CP(wclk), .Q(ram[5744]) );
  DFF ram_reg_1337__7_ ( .D(n9928), .CP(wclk), .Q(ram[5687]) );
  DFF ram_reg_1337__6_ ( .D(n9927), .CP(wclk), .Q(ram[5686]) );
  DFF ram_reg_1337__5_ ( .D(n9926), .CP(wclk), .Q(ram[5685]) );
  DFF ram_reg_1337__4_ ( .D(n9925), .CP(wclk), .Q(ram[5684]) );
  DFF ram_reg_1337__3_ ( .D(n9924), .CP(wclk), .Q(ram[5683]) );
  DFF ram_reg_1337__2_ ( .D(n9923), .CP(wclk), .Q(ram[5682]) );
  DFF ram_reg_1337__1_ ( .D(n9922), .CP(wclk), .Q(ram[5681]) );
  DFF ram_reg_1337__0_ ( .D(n9921), .CP(wclk), .Q(ram[5680]) );
  DFF ram_reg_1341__7_ ( .D(n9896), .CP(wclk), .Q(ram[5655]) );
  DFF ram_reg_1341__6_ ( .D(n9895), .CP(wclk), .Q(ram[5654]) );
  DFF ram_reg_1341__5_ ( .D(n9894), .CP(wclk), .Q(ram[5653]) );
  DFF ram_reg_1341__4_ ( .D(n9893), .CP(wclk), .Q(ram[5652]) );
  DFF ram_reg_1341__3_ ( .D(n9892), .CP(wclk), .Q(ram[5651]) );
  DFF ram_reg_1341__2_ ( .D(n9891), .CP(wclk), .Q(ram[5650]) );
  DFF ram_reg_1341__1_ ( .D(n9890), .CP(wclk), .Q(ram[5649]) );
  DFF ram_reg_1341__0_ ( .D(n9889), .CP(wclk), .Q(ram[5648]) );
  DFF ram_reg_1353__7_ ( .D(n9800), .CP(wclk), .Q(ram[5559]) );
  DFF ram_reg_1353__6_ ( .D(n9799), .CP(wclk), .Q(ram[5558]) );
  DFF ram_reg_1353__5_ ( .D(n9798), .CP(wclk), .Q(ram[5557]) );
  DFF ram_reg_1353__4_ ( .D(n9797), .CP(wclk), .Q(ram[5556]) );
  DFF ram_reg_1353__3_ ( .D(n9796), .CP(wclk), .Q(ram[5555]) );
  DFF ram_reg_1353__2_ ( .D(n9795), .CP(wclk), .Q(ram[5554]) );
  DFF ram_reg_1353__1_ ( .D(n9794), .CP(wclk), .Q(ram[5553]) );
  DFF ram_reg_1353__0_ ( .D(n9793), .CP(wclk), .Q(ram[5552]) );
  DFF ram_reg_1357__7_ ( .D(n9768), .CP(wclk), .Q(ram[5527]) );
  DFF ram_reg_1357__6_ ( .D(n9767), .CP(wclk), .Q(ram[5526]) );
  DFF ram_reg_1357__5_ ( .D(n9766), .CP(wclk), .Q(ram[5525]) );
  DFF ram_reg_1357__4_ ( .D(n9765), .CP(wclk), .Q(ram[5524]) );
  DFF ram_reg_1357__3_ ( .D(n9764), .CP(wclk), .Q(ram[5523]) );
  DFF ram_reg_1357__2_ ( .D(n9763), .CP(wclk), .Q(ram[5522]) );
  DFF ram_reg_1357__1_ ( .D(n9762), .CP(wclk), .Q(ram[5521]) );
  DFF ram_reg_1357__0_ ( .D(n9761), .CP(wclk), .Q(ram[5520]) );
  DFF ram_reg_1369__7_ ( .D(n9672), .CP(wclk), .Q(ram[5431]) );
  DFF ram_reg_1369__6_ ( .D(n9671), .CP(wclk), .Q(ram[5430]) );
  DFF ram_reg_1369__5_ ( .D(n9670), .CP(wclk), .Q(ram[5429]) );
  DFF ram_reg_1369__4_ ( .D(n9669), .CP(wclk), .Q(ram[5428]) );
  DFF ram_reg_1369__3_ ( .D(n9668), .CP(wclk), .Q(ram[5427]) );
  DFF ram_reg_1369__2_ ( .D(n9667), .CP(wclk), .Q(ram[5426]) );
  DFF ram_reg_1369__1_ ( .D(n9666), .CP(wclk), .Q(ram[5425]) );
  DFF ram_reg_1369__0_ ( .D(n9665), .CP(wclk), .Q(ram[5424]) );
  DFF ram_reg_1385__7_ ( .D(n9544), .CP(wclk), .Q(ram[5303]) );
  DFF ram_reg_1385__6_ ( .D(n9543), .CP(wclk), .Q(ram[5302]) );
  DFF ram_reg_1385__5_ ( .D(n9542), .CP(wclk), .Q(ram[5301]) );
  DFF ram_reg_1385__4_ ( .D(n9541), .CP(wclk), .Q(ram[5300]) );
  DFF ram_reg_1385__3_ ( .D(n9540), .CP(wclk), .Q(ram[5299]) );
  DFF ram_reg_1385__2_ ( .D(n9539), .CP(wclk), .Q(ram[5298]) );
  DFF ram_reg_1385__1_ ( .D(n9538), .CP(wclk), .Q(ram[5297]) );
  DFF ram_reg_1385__0_ ( .D(n9537), .CP(wclk), .Q(ram[5296]) );
  DFF ram_reg_1389__7_ ( .D(n9512), .CP(wclk), .Q(ram[5271]) );
  DFF ram_reg_1389__6_ ( .D(n9511), .CP(wclk), .Q(ram[5270]) );
  DFF ram_reg_1389__5_ ( .D(n9510), .CP(wclk), .Q(ram[5269]) );
  DFF ram_reg_1389__4_ ( .D(n9509), .CP(wclk), .Q(ram[5268]) );
  DFF ram_reg_1389__3_ ( .D(n9508), .CP(wclk), .Q(ram[5267]) );
  DFF ram_reg_1389__2_ ( .D(n9507), .CP(wclk), .Q(ram[5266]) );
  DFF ram_reg_1389__1_ ( .D(n9506), .CP(wclk), .Q(ram[5265]) );
  DFF ram_reg_1389__0_ ( .D(n9505), .CP(wclk), .Q(ram[5264]) );
  DFF ram_reg_1401__7_ ( .D(n9416), .CP(wclk), .Q(ram[5175]) );
  DFF ram_reg_1401__6_ ( .D(n9415), .CP(wclk), .Q(ram[5174]) );
  DFF ram_reg_1401__5_ ( .D(n9414), .CP(wclk), .Q(ram[5173]) );
  DFF ram_reg_1401__4_ ( .D(n9413), .CP(wclk), .Q(ram[5172]) );
  DFF ram_reg_1401__3_ ( .D(n9412), .CP(wclk), .Q(ram[5171]) );
  DFF ram_reg_1401__2_ ( .D(n9411), .CP(wclk), .Q(ram[5170]) );
  DFF ram_reg_1401__1_ ( .D(n9410), .CP(wclk), .Q(ram[5169]) );
  DFF ram_reg_1401__0_ ( .D(n9409), .CP(wclk), .Q(ram[5168]) );
  DFF ram_reg_1405__7_ ( .D(n9384), .CP(wclk), .Q(ram[5143]) );
  DFF ram_reg_1405__6_ ( .D(n9383), .CP(wclk), .Q(ram[5142]) );
  DFF ram_reg_1405__5_ ( .D(n9382), .CP(wclk), .Q(ram[5141]) );
  DFF ram_reg_1405__4_ ( .D(n9381), .CP(wclk), .Q(ram[5140]) );
  DFF ram_reg_1405__3_ ( .D(n9380), .CP(wclk), .Q(ram[5139]) );
  DFF ram_reg_1405__2_ ( .D(n9379), .CP(wclk), .Q(ram[5138]) );
  DFF ram_reg_1405__1_ ( .D(n9378), .CP(wclk), .Q(ram[5137]) );
  DFF ram_reg_1405__0_ ( .D(n9377), .CP(wclk), .Q(ram[5136]) );
  DFF ram_reg_1409__7_ ( .D(n9352), .CP(wclk), .Q(ram[5111]) );
  DFF ram_reg_1409__6_ ( .D(n9351), .CP(wclk), .Q(ram[5110]) );
  DFF ram_reg_1409__5_ ( .D(n9350), .CP(wclk), .Q(ram[5109]) );
  DFF ram_reg_1409__4_ ( .D(n9349), .CP(wclk), .Q(ram[5108]) );
  DFF ram_reg_1409__3_ ( .D(n9348), .CP(wclk), .Q(ram[5107]) );
  DFF ram_reg_1409__2_ ( .D(n9347), .CP(wclk), .Q(ram[5106]) );
  DFF ram_reg_1409__1_ ( .D(n9346), .CP(wclk), .Q(ram[5105]) );
  DFF ram_reg_1409__0_ ( .D(n9345), .CP(wclk), .Q(ram[5104]) );
  DFF ram_reg_1413__7_ ( .D(n9320), .CP(wclk), .Q(ram[5079]) );
  DFF ram_reg_1413__6_ ( .D(n9319), .CP(wclk), .Q(ram[5078]) );
  DFF ram_reg_1413__5_ ( .D(n9318), .CP(wclk), .Q(ram[5077]) );
  DFF ram_reg_1413__4_ ( .D(n9317), .CP(wclk), .Q(ram[5076]) );
  DFF ram_reg_1413__3_ ( .D(n9316), .CP(wclk), .Q(ram[5075]) );
  DFF ram_reg_1413__2_ ( .D(n9315), .CP(wclk), .Q(ram[5074]) );
  DFF ram_reg_1413__1_ ( .D(n9314), .CP(wclk), .Q(ram[5073]) );
  DFF ram_reg_1413__0_ ( .D(n9313), .CP(wclk), .Q(ram[5072]) );
  DFF ram_reg_1417__7_ ( .D(n9288), .CP(wclk), .Q(ram[5047]) );
  DFF ram_reg_1417__6_ ( .D(n9287), .CP(wclk), .Q(ram[5046]) );
  DFF ram_reg_1417__5_ ( .D(n9286), .CP(wclk), .Q(ram[5045]) );
  DFF ram_reg_1417__4_ ( .D(n9285), .CP(wclk), .Q(ram[5044]) );
  DFF ram_reg_1417__3_ ( .D(n9284), .CP(wclk), .Q(ram[5043]) );
  DFF ram_reg_1417__2_ ( .D(n9283), .CP(wclk), .Q(ram[5042]) );
  DFF ram_reg_1417__1_ ( .D(n9282), .CP(wclk), .Q(ram[5041]) );
  DFF ram_reg_1417__0_ ( .D(n9281), .CP(wclk), .Q(ram[5040]) );
  DFF ram_reg_1421__7_ ( .D(n9256), .CP(wclk), .Q(ram[5015]) );
  DFF ram_reg_1421__6_ ( .D(n9255), .CP(wclk), .Q(ram[5014]) );
  DFF ram_reg_1421__5_ ( .D(n9254), .CP(wclk), .Q(ram[5013]) );
  DFF ram_reg_1421__4_ ( .D(n9253), .CP(wclk), .Q(ram[5012]) );
  DFF ram_reg_1421__3_ ( .D(n9252), .CP(wclk), .Q(ram[5011]) );
  DFF ram_reg_1421__2_ ( .D(n9251), .CP(wclk), .Q(ram[5010]) );
  DFF ram_reg_1421__1_ ( .D(n9250), .CP(wclk), .Q(ram[5009]) );
  DFF ram_reg_1421__0_ ( .D(n9249), .CP(wclk), .Q(ram[5008]) );
  DFF ram_reg_1425__7_ ( .D(n9224), .CP(wclk), .Q(ram[4983]) );
  DFF ram_reg_1425__6_ ( .D(n9223), .CP(wclk), .Q(ram[4982]) );
  DFF ram_reg_1425__5_ ( .D(n9222), .CP(wclk), .Q(ram[4981]) );
  DFF ram_reg_1425__4_ ( .D(n9221), .CP(wclk), .Q(ram[4980]) );
  DFF ram_reg_1425__3_ ( .D(n9220), .CP(wclk), .Q(ram[4979]) );
  DFF ram_reg_1425__2_ ( .D(n9219), .CP(wclk), .Q(ram[4978]) );
  DFF ram_reg_1425__1_ ( .D(n9218), .CP(wclk), .Q(ram[4977]) );
  DFF ram_reg_1425__0_ ( .D(n9217), .CP(wclk), .Q(ram[4976]) );
  DFF ram_reg_1429__7_ ( .D(n9192), .CP(wclk), .Q(ram[4951]) );
  DFF ram_reg_1429__6_ ( .D(n9191), .CP(wclk), .Q(ram[4950]) );
  DFF ram_reg_1429__5_ ( .D(n9190), .CP(wclk), .Q(ram[4949]) );
  DFF ram_reg_1429__4_ ( .D(n9189), .CP(wclk), .Q(ram[4948]) );
  DFF ram_reg_1429__3_ ( .D(n9188), .CP(wclk), .Q(ram[4947]) );
  DFF ram_reg_1429__2_ ( .D(n9187), .CP(wclk), .Q(ram[4946]) );
  DFF ram_reg_1429__1_ ( .D(n9186), .CP(wclk), .Q(ram[4945]) );
  DFF ram_reg_1429__0_ ( .D(n9185), .CP(wclk), .Q(ram[4944]) );
  DFF ram_reg_1433__7_ ( .D(n9160), .CP(wclk), .Q(ram[4919]) );
  DFF ram_reg_1433__6_ ( .D(n9159), .CP(wclk), .Q(ram[4918]) );
  DFF ram_reg_1433__5_ ( .D(n9158), .CP(wclk), .Q(ram[4917]) );
  DFF ram_reg_1433__4_ ( .D(n9157), .CP(wclk), .Q(ram[4916]) );
  DFF ram_reg_1433__3_ ( .D(n9156), .CP(wclk), .Q(ram[4915]) );
  DFF ram_reg_1433__2_ ( .D(n9155), .CP(wclk), .Q(ram[4914]) );
  DFF ram_reg_1433__1_ ( .D(n9154), .CP(wclk), .Q(ram[4913]) );
  DFF ram_reg_1433__0_ ( .D(n9153), .CP(wclk), .Q(ram[4912]) );
  DFF ram_reg_1437__7_ ( .D(n9128), .CP(wclk), .Q(ram[4887]) );
  DFF ram_reg_1437__6_ ( .D(n9127), .CP(wclk), .Q(ram[4886]) );
  DFF ram_reg_1437__5_ ( .D(n9126), .CP(wclk), .Q(ram[4885]) );
  DFF ram_reg_1437__4_ ( .D(n9125), .CP(wclk), .Q(ram[4884]) );
  DFF ram_reg_1437__3_ ( .D(n9124), .CP(wclk), .Q(ram[4883]) );
  DFF ram_reg_1437__2_ ( .D(n9123), .CP(wclk), .Q(ram[4882]) );
  DFF ram_reg_1437__1_ ( .D(n9122), .CP(wclk), .Q(ram[4881]) );
  DFF ram_reg_1437__0_ ( .D(n9121), .CP(wclk), .Q(ram[4880]) );
  DFF ram_reg_1441__7_ ( .D(n9096), .CP(wclk), .Q(ram[4855]) );
  DFF ram_reg_1441__6_ ( .D(n9095), .CP(wclk), .Q(ram[4854]) );
  DFF ram_reg_1441__5_ ( .D(n9094), .CP(wclk), .Q(ram[4853]) );
  DFF ram_reg_1441__4_ ( .D(n9093), .CP(wclk), .Q(ram[4852]) );
  DFF ram_reg_1441__3_ ( .D(n9092), .CP(wclk), .Q(ram[4851]) );
  DFF ram_reg_1441__2_ ( .D(n9091), .CP(wclk), .Q(ram[4850]) );
  DFF ram_reg_1441__1_ ( .D(n9090), .CP(wclk), .Q(ram[4849]) );
  DFF ram_reg_1441__0_ ( .D(n9089), .CP(wclk), .Q(ram[4848]) );
  DFF ram_reg_1445__7_ ( .D(n9064), .CP(wclk), .Q(ram[4823]) );
  DFF ram_reg_1445__6_ ( .D(n9063), .CP(wclk), .Q(ram[4822]) );
  DFF ram_reg_1445__5_ ( .D(n9062), .CP(wclk), .Q(ram[4821]) );
  DFF ram_reg_1445__4_ ( .D(n9061), .CP(wclk), .Q(ram[4820]) );
  DFF ram_reg_1445__3_ ( .D(n9060), .CP(wclk), .Q(ram[4819]) );
  DFF ram_reg_1445__2_ ( .D(n9059), .CP(wclk), .Q(ram[4818]) );
  DFF ram_reg_1445__1_ ( .D(n9058), .CP(wclk), .Q(ram[4817]) );
  DFF ram_reg_1445__0_ ( .D(n9057), .CP(wclk), .Q(ram[4816]) );
  DFF ram_reg_1449__7_ ( .D(n9032), .CP(wclk), .Q(ram[4791]) );
  DFF ram_reg_1449__6_ ( .D(n9031), .CP(wclk), .Q(ram[4790]) );
  DFF ram_reg_1449__5_ ( .D(n9030), .CP(wclk), .Q(ram[4789]) );
  DFF ram_reg_1449__4_ ( .D(n9029), .CP(wclk), .Q(ram[4788]) );
  DFF ram_reg_1449__3_ ( .D(n9028), .CP(wclk), .Q(ram[4787]) );
  DFF ram_reg_1449__2_ ( .D(n9027), .CP(wclk), .Q(ram[4786]) );
  DFF ram_reg_1449__1_ ( .D(n9026), .CP(wclk), .Q(ram[4785]) );
  DFF ram_reg_1449__0_ ( .D(n9025), .CP(wclk), .Q(ram[4784]) );
  DFF ram_reg_1453__7_ ( .D(n9000), .CP(wclk), .Q(ram[4759]) );
  DFF ram_reg_1453__6_ ( .D(n8999), .CP(wclk), .Q(ram[4758]) );
  DFF ram_reg_1453__5_ ( .D(n8998), .CP(wclk), .Q(ram[4757]) );
  DFF ram_reg_1453__4_ ( .D(n8997), .CP(wclk), .Q(ram[4756]) );
  DFF ram_reg_1453__3_ ( .D(n8996), .CP(wclk), .Q(ram[4755]) );
  DFF ram_reg_1453__2_ ( .D(n8995), .CP(wclk), .Q(ram[4754]) );
  DFF ram_reg_1453__1_ ( .D(n8994), .CP(wclk), .Q(ram[4753]) );
  DFF ram_reg_1453__0_ ( .D(n8993), .CP(wclk), .Q(ram[4752]) );
  DFF ram_reg_1457__7_ ( .D(n8968), .CP(wclk), .Q(ram[4727]) );
  DFF ram_reg_1457__6_ ( .D(n8967), .CP(wclk), .Q(ram[4726]) );
  DFF ram_reg_1457__5_ ( .D(n8966), .CP(wclk), .Q(ram[4725]) );
  DFF ram_reg_1457__4_ ( .D(n8965), .CP(wclk), .Q(ram[4724]) );
  DFF ram_reg_1457__3_ ( .D(n8964), .CP(wclk), .Q(ram[4723]) );
  DFF ram_reg_1457__2_ ( .D(n8963), .CP(wclk), .Q(ram[4722]) );
  DFF ram_reg_1457__1_ ( .D(n8962), .CP(wclk), .Q(ram[4721]) );
  DFF ram_reg_1457__0_ ( .D(n8961), .CP(wclk), .Q(ram[4720]) );
  DFF ram_reg_1461__7_ ( .D(n8936), .CP(wclk), .Q(ram[4695]) );
  DFF ram_reg_1461__6_ ( .D(n8935), .CP(wclk), .Q(ram[4694]) );
  DFF ram_reg_1461__5_ ( .D(n8934), .CP(wclk), .Q(ram[4693]) );
  DFF ram_reg_1461__4_ ( .D(n8933), .CP(wclk), .Q(ram[4692]) );
  DFF ram_reg_1461__3_ ( .D(n8932), .CP(wclk), .Q(ram[4691]) );
  DFF ram_reg_1461__2_ ( .D(n8931), .CP(wclk), .Q(ram[4690]) );
  DFF ram_reg_1461__1_ ( .D(n8930), .CP(wclk), .Q(ram[4689]) );
  DFF ram_reg_1461__0_ ( .D(n8929), .CP(wclk), .Q(ram[4688]) );
  DFF ram_reg_1465__7_ ( .D(n8904), .CP(wclk), .Q(ram[4663]) );
  DFF ram_reg_1465__6_ ( .D(n8903), .CP(wclk), .Q(ram[4662]) );
  DFF ram_reg_1465__5_ ( .D(n8902), .CP(wclk), .Q(ram[4661]) );
  DFF ram_reg_1465__4_ ( .D(n8901), .CP(wclk), .Q(ram[4660]) );
  DFF ram_reg_1465__3_ ( .D(n8900), .CP(wclk), .Q(ram[4659]) );
  DFF ram_reg_1465__2_ ( .D(n8899), .CP(wclk), .Q(ram[4658]) );
  DFF ram_reg_1465__1_ ( .D(n8898), .CP(wclk), .Q(ram[4657]) );
  DFF ram_reg_1465__0_ ( .D(n8897), .CP(wclk), .Q(ram[4656]) );
  DFF ram_reg_1469__7_ ( .D(n8872), .CP(wclk), .Q(ram[4631]) );
  DFF ram_reg_1469__6_ ( .D(n8871), .CP(wclk), .Q(ram[4630]) );
  DFF ram_reg_1469__5_ ( .D(n8870), .CP(wclk), .Q(ram[4629]) );
  DFF ram_reg_1469__4_ ( .D(n8869), .CP(wclk), .Q(ram[4628]) );
  DFF ram_reg_1469__3_ ( .D(n8868), .CP(wclk), .Q(ram[4627]) );
  DFF ram_reg_1469__2_ ( .D(n8867), .CP(wclk), .Q(ram[4626]) );
  DFF ram_reg_1469__1_ ( .D(n8866), .CP(wclk), .Q(ram[4625]) );
  DFF ram_reg_1469__0_ ( .D(n8865), .CP(wclk), .Q(ram[4624]) );
  DFF ram_reg_1473__7_ ( .D(n8840), .CP(wclk), .Q(ram[4599]) );
  DFF ram_reg_1473__6_ ( .D(n8839), .CP(wclk), .Q(ram[4598]) );
  DFF ram_reg_1473__5_ ( .D(n8838), .CP(wclk), .Q(ram[4597]) );
  DFF ram_reg_1473__4_ ( .D(n8837), .CP(wclk), .Q(ram[4596]) );
  DFF ram_reg_1473__3_ ( .D(n8836), .CP(wclk), .Q(ram[4595]) );
  DFF ram_reg_1473__2_ ( .D(n8835), .CP(wclk), .Q(ram[4594]) );
  DFF ram_reg_1473__1_ ( .D(n8834), .CP(wclk), .Q(ram[4593]) );
  DFF ram_reg_1473__0_ ( .D(n8833), .CP(wclk), .Q(ram[4592]) );
  DFF ram_reg_1477__7_ ( .D(n8808), .CP(wclk), .Q(ram[4567]) );
  DFF ram_reg_1477__6_ ( .D(n8807), .CP(wclk), .Q(ram[4566]) );
  DFF ram_reg_1477__5_ ( .D(n8806), .CP(wclk), .Q(ram[4565]) );
  DFF ram_reg_1477__4_ ( .D(n8805), .CP(wclk), .Q(ram[4564]) );
  DFF ram_reg_1477__3_ ( .D(n8804), .CP(wclk), .Q(ram[4563]) );
  DFF ram_reg_1477__2_ ( .D(n8803), .CP(wclk), .Q(ram[4562]) );
  DFF ram_reg_1477__1_ ( .D(n8802), .CP(wclk), .Q(ram[4561]) );
  DFF ram_reg_1477__0_ ( .D(n8801), .CP(wclk), .Q(ram[4560]) );
  DFF ram_reg_1481__7_ ( .D(n8776), .CP(wclk), .Q(ram[4535]) );
  DFF ram_reg_1481__6_ ( .D(n8775), .CP(wclk), .Q(ram[4534]) );
  DFF ram_reg_1481__5_ ( .D(n8774), .CP(wclk), .Q(ram[4533]) );
  DFF ram_reg_1481__4_ ( .D(n8773), .CP(wclk), .Q(ram[4532]) );
  DFF ram_reg_1481__3_ ( .D(n8772), .CP(wclk), .Q(ram[4531]) );
  DFF ram_reg_1481__2_ ( .D(n8771), .CP(wclk), .Q(ram[4530]) );
  DFF ram_reg_1481__1_ ( .D(n8770), .CP(wclk), .Q(ram[4529]) );
  DFF ram_reg_1481__0_ ( .D(n8769), .CP(wclk), .Q(ram[4528]) );
  DFF ram_reg_1485__7_ ( .D(n8744), .CP(wclk), .Q(ram[4503]) );
  DFF ram_reg_1485__6_ ( .D(n8743), .CP(wclk), .Q(ram[4502]) );
  DFF ram_reg_1485__5_ ( .D(n8742), .CP(wclk), .Q(ram[4501]) );
  DFF ram_reg_1485__4_ ( .D(n8741), .CP(wclk), .Q(ram[4500]) );
  DFF ram_reg_1485__3_ ( .D(n8740), .CP(wclk), .Q(ram[4499]) );
  DFF ram_reg_1485__2_ ( .D(n8739), .CP(wclk), .Q(ram[4498]) );
  DFF ram_reg_1485__1_ ( .D(n8738), .CP(wclk), .Q(ram[4497]) );
  DFF ram_reg_1485__0_ ( .D(n8737), .CP(wclk), .Q(ram[4496]) );
  DFF ram_reg_1489__7_ ( .D(n8712), .CP(wclk), .Q(ram[4471]) );
  DFF ram_reg_1489__6_ ( .D(n8711), .CP(wclk), .Q(ram[4470]) );
  DFF ram_reg_1489__5_ ( .D(n8710), .CP(wclk), .Q(ram[4469]) );
  DFF ram_reg_1489__4_ ( .D(n8709), .CP(wclk), .Q(ram[4468]) );
  DFF ram_reg_1489__3_ ( .D(n8708), .CP(wclk), .Q(ram[4467]) );
  DFF ram_reg_1489__2_ ( .D(n8707), .CP(wclk), .Q(ram[4466]) );
  DFF ram_reg_1489__1_ ( .D(n8706), .CP(wclk), .Q(ram[4465]) );
  DFF ram_reg_1489__0_ ( .D(n8705), .CP(wclk), .Q(ram[4464]) );
  DFF ram_reg_1497__7_ ( .D(n8648), .CP(wclk), .Q(ram[4407]) );
  DFF ram_reg_1497__6_ ( .D(n8647), .CP(wclk), .Q(ram[4406]) );
  DFF ram_reg_1497__5_ ( .D(n8646), .CP(wclk), .Q(ram[4405]) );
  DFF ram_reg_1497__4_ ( .D(n8645), .CP(wclk), .Q(ram[4404]) );
  DFF ram_reg_1497__3_ ( .D(n8644), .CP(wclk), .Q(ram[4403]) );
  DFF ram_reg_1497__2_ ( .D(n8643), .CP(wclk), .Q(ram[4402]) );
  DFF ram_reg_1497__1_ ( .D(n8642), .CP(wclk), .Q(ram[4401]) );
  DFF ram_reg_1497__0_ ( .D(n8641), .CP(wclk), .Q(ram[4400]) );
  DFF ram_reg_1501__7_ ( .D(n8616), .CP(wclk), .Q(ram[4375]) );
  DFF ram_reg_1501__6_ ( .D(n8615), .CP(wclk), .Q(ram[4374]) );
  DFF ram_reg_1501__5_ ( .D(n8614), .CP(wclk), .Q(ram[4373]) );
  DFF ram_reg_1501__4_ ( .D(n8613), .CP(wclk), .Q(ram[4372]) );
  DFF ram_reg_1501__3_ ( .D(n8612), .CP(wclk), .Q(ram[4371]) );
  DFF ram_reg_1501__2_ ( .D(n8611), .CP(wclk), .Q(ram[4370]) );
  DFF ram_reg_1501__1_ ( .D(n8610), .CP(wclk), .Q(ram[4369]) );
  DFF ram_reg_1501__0_ ( .D(n8609), .CP(wclk), .Q(ram[4368]) );
  DFF ram_reg_1505__7_ ( .D(n8584), .CP(wclk), .Q(ram[4343]) );
  DFF ram_reg_1505__6_ ( .D(n8583), .CP(wclk), .Q(ram[4342]) );
  DFF ram_reg_1505__5_ ( .D(n8582), .CP(wclk), .Q(ram[4341]) );
  DFF ram_reg_1505__4_ ( .D(n8581), .CP(wclk), .Q(ram[4340]) );
  DFF ram_reg_1505__3_ ( .D(n8580), .CP(wclk), .Q(ram[4339]) );
  DFF ram_reg_1505__2_ ( .D(n8579), .CP(wclk), .Q(ram[4338]) );
  DFF ram_reg_1505__1_ ( .D(n8578), .CP(wclk), .Q(ram[4337]) );
  DFF ram_reg_1505__0_ ( .D(n8577), .CP(wclk), .Q(ram[4336]) );
  DFF ram_reg_1509__7_ ( .D(n8552), .CP(wclk), .Q(ram[4311]) );
  DFF ram_reg_1509__6_ ( .D(n8551), .CP(wclk), .Q(ram[4310]) );
  DFF ram_reg_1509__5_ ( .D(n8550), .CP(wclk), .Q(ram[4309]) );
  DFF ram_reg_1509__4_ ( .D(n8549), .CP(wclk), .Q(ram[4308]) );
  DFF ram_reg_1509__3_ ( .D(n8548), .CP(wclk), .Q(ram[4307]) );
  DFF ram_reg_1509__2_ ( .D(n8547), .CP(wclk), .Q(ram[4306]) );
  DFF ram_reg_1509__1_ ( .D(n8546), .CP(wclk), .Q(ram[4305]) );
  DFF ram_reg_1509__0_ ( .D(n8545), .CP(wclk), .Q(ram[4304]) );
  DFF ram_reg_1513__7_ ( .D(n8520), .CP(wclk), .Q(ram[4279]) );
  DFF ram_reg_1513__6_ ( .D(n8519), .CP(wclk), .Q(ram[4278]) );
  DFF ram_reg_1513__5_ ( .D(n8518), .CP(wclk), .Q(ram[4277]) );
  DFF ram_reg_1513__4_ ( .D(n8517), .CP(wclk), .Q(ram[4276]) );
  DFF ram_reg_1513__3_ ( .D(n8516), .CP(wclk), .Q(ram[4275]) );
  DFF ram_reg_1513__2_ ( .D(n8515), .CP(wclk), .Q(ram[4274]) );
  DFF ram_reg_1513__1_ ( .D(n8514), .CP(wclk), .Q(ram[4273]) );
  DFF ram_reg_1513__0_ ( .D(n8513), .CP(wclk), .Q(ram[4272]) );
  DFF ram_reg_1517__7_ ( .D(n8488), .CP(wclk), .Q(ram[4247]) );
  DFF ram_reg_1517__6_ ( .D(n8487), .CP(wclk), .Q(ram[4246]) );
  DFF ram_reg_1517__5_ ( .D(n8486), .CP(wclk), .Q(ram[4245]) );
  DFF ram_reg_1517__4_ ( .D(n8485), .CP(wclk), .Q(ram[4244]) );
  DFF ram_reg_1517__3_ ( .D(n8484), .CP(wclk), .Q(ram[4243]) );
  DFF ram_reg_1517__2_ ( .D(n8483), .CP(wclk), .Q(ram[4242]) );
  DFF ram_reg_1517__1_ ( .D(n8482), .CP(wclk), .Q(ram[4241]) );
  DFF ram_reg_1517__0_ ( .D(n8481), .CP(wclk), .Q(ram[4240]) );
  DFF ram_reg_1521__7_ ( .D(n8456), .CP(wclk), .Q(ram[4215]) );
  DFF ram_reg_1521__6_ ( .D(n8455), .CP(wclk), .Q(ram[4214]) );
  DFF ram_reg_1521__5_ ( .D(n8454), .CP(wclk), .Q(ram[4213]) );
  DFF ram_reg_1521__4_ ( .D(n8453), .CP(wclk), .Q(ram[4212]) );
  DFF ram_reg_1521__3_ ( .D(n8452), .CP(wclk), .Q(ram[4211]) );
  DFF ram_reg_1521__2_ ( .D(n8451), .CP(wclk), .Q(ram[4210]) );
  DFF ram_reg_1521__1_ ( .D(n8450), .CP(wclk), .Q(ram[4209]) );
  DFF ram_reg_1521__0_ ( .D(n8449), .CP(wclk), .Q(ram[4208]) );
  DFF ram_reg_1525__7_ ( .D(n8424), .CP(wclk), .Q(ram[4183]) );
  DFF ram_reg_1525__6_ ( .D(n8423), .CP(wclk), .Q(ram[4182]) );
  DFF ram_reg_1525__5_ ( .D(n8422), .CP(wclk), .Q(ram[4181]) );
  DFF ram_reg_1525__4_ ( .D(n8421), .CP(wclk), .Q(ram[4180]) );
  DFF ram_reg_1525__3_ ( .D(n8420), .CP(wclk), .Q(ram[4179]) );
  DFF ram_reg_1525__2_ ( .D(n8419), .CP(wclk), .Q(ram[4178]) );
  DFF ram_reg_1525__1_ ( .D(n8418), .CP(wclk), .Q(ram[4177]) );
  DFF ram_reg_1525__0_ ( .D(n8417), .CP(wclk), .Q(ram[4176]) );
  DFF ram_reg_1529__7_ ( .D(n8392), .CP(wclk), .Q(ram[4151]) );
  DFF ram_reg_1529__6_ ( .D(n8391), .CP(wclk), .Q(ram[4150]) );
  DFF ram_reg_1529__5_ ( .D(n8390), .CP(wclk), .Q(ram[4149]) );
  DFF ram_reg_1529__4_ ( .D(n8389), .CP(wclk), .Q(ram[4148]) );
  DFF ram_reg_1529__3_ ( .D(n8388), .CP(wclk), .Q(ram[4147]) );
  DFF ram_reg_1529__2_ ( .D(n8387), .CP(wclk), .Q(ram[4146]) );
  DFF ram_reg_1529__1_ ( .D(n8386), .CP(wclk), .Q(ram[4145]) );
  DFF ram_reg_1529__0_ ( .D(n8385), .CP(wclk), .Q(ram[4144]) );
  DFF ram_reg_1533__7_ ( .D(n8360), .CP(wclk), .Q(ram[4119]) );
  DFF ram_reg_1533__6_ ( .D(n8359), .CP(wclk), .Q(ram[4118]) );
  DFF ram_reg_1533__5_ ( .D(n8358), .CP(wclk), .Q(ram[4117]) );
  DFF ram_reg_1533__4_ ( .D(n8357), .CP(wclk), .Q(ram[4116]) );
  DFF ram_reg_1533__3_ ( .D(n8356), .CP(wclk), .Q(ram[4115]) );
  DFF ram_reg_1533__2_ ( .D(n8355), .CP(wclk), .Q(ram[4114]) );
  DFF ram_reg_1533__1_ ( .D(n8354), .CP(wclk), .Q(ram[4113]) );
  DFF ram_reg_1533__0_ ( .D(n8353), .CP(wclk), .Q(ram[4112]) );
  DFF ram_reg_1545__7_ ( .D(n8264), .CP(wclk), .Q(ram[4023]) );
  DFF ram_reg_1545__6_ ( .D(n8263), .CP(wclk), .Q(ram[4022]) );
  DFF ram_reg_1545__5_ ( .D(n8262), .CP(wclk), .Q(ram[4021]) );
  DFF ram_reg_1545__4_ ( .D(n8261), .CP(wclk), .Q(ram[4020]) );
  DFF ram_reg_1545__3_ ( .D(n8260), .CP(wclk), .Q(ram[4019]) );
  DFF ram_reg_1545__2_ ( .D(n8259), .CP(wclk), .Q(ram[4018]) );
  DFF ram_reg_1545__1_ ( .D(n8258), .CP(wclk), .Q(ram[4017]) );
  DFF ram_reg_1545__0_ ( .D(n8257), .CP(wclk), .Q(ram[4016]) );
  DFF ram_reg_1549__7_ ( .D(n8232), .CP(wclk), .Q(ram[3991]) );
  DFF ram_reg_1549__6_ ( .D(n8231), .CP(wclk), .Q(ram[3990]) );
  DFF ram_reg_1549__5_ ( .D(n8230), .CP(wclk), .Q(ram[3989]) );
  DFF ram_reg_1549__4_ ( .D(n8229), .CP(wclk), .Q(ram[3988]) );
  DFF ram_reg_1549__3_ ( .D(n8228), .CP(wclk), .Q(ram[3987]) );
  DFF ram_reg_1549__2_ ( .D(n8227), .CP(wclk), .Q(ram[3986]) );
  DFF ram_reg_1549__1_ ( .D(n8226), .CP(wclk), .Q(ram[3985]) );
  DFF ram_reg_1549__0_ ( .D(n8225), .CP(wclk), .Q(ram[3984]) );
  DFF ram_reg_1561__7_ ( .D(n8136), .CP(wclk), .Q(ram[3895]) );
  DFF ram_reg_1561__6_ ( .D(n8135), .CP(wclk), .Q(ram[3894]) );
  DFF ram_reg_1561__5_ ( .D(n8134), .CP(wclk), .Q(ram[3893]) );
  DFF ram_reg_1561__4_ ( .D(n8133), .CP(wclk), .Q(ram[3892]) );
  DFF ram_reg_1561__3_ ( .D(n8132), .CP(wclk), .Q(ram[3891]) );
  DFF ram_reg_1561__2_ ( .D(n8131), .CP(wclk), .Q(ram[3890]) );
  DFF ram_reg_1561__1_ ( .D(n8130), .CP(wclk), .Q(ram[3889]) );
  DFF ram_reg_1561__0_ ( .D(n8129), .CP(wclk), .Q(ram[3888]) );
  DFF ram_reg_1577__7_ ( .D(n8008), .CP(wclk), .Q(ram[3767]) );
  DFF ram_reg_1577__6_ ( .D(n8007), .CP(wclk), .Q(ram[3766]) );
  DFF ram_reg_1577__5_ ( .D(n8006), .CP(wclk), .Q(ram[3765]) );
  DFF ram_reg_1577__4_ ( .D(n8005), .CP(wclk), .Q(ram[3764]) );
  DFF ram_reg_1577__3_ ( .D(n8004), .CP(wclk), .Q(ram[3763]) );
  DFF ram_reg_1577__2_ ( .D(n8003), .CP(wclk), .Q(ram[3762]) );
  DFF ram_reg_1577__1_ ( .D(n8002), .CP(wclk), .Q(ram[3761]) );
  DFF ram_reg_1577__0_ ( .D(n8001), .CP(wclk), .Q(ram[3760]) );
  DFF ram_reg_1581__7_ ( .D(n7976), .CP(wclk), .Q(ram[3735]) );
  DFF ram_reg_1581__6_ ( .D(n7975), .CP(wclk), .Q(ram[3734]) );
  DFF ram_reg_1581__5_ ( .D(n7974), .CP(wclk), .Q(ram[3733]) );
  DFF ram_reg_1581__4_ ( .D(n7973), .CP(wclk), .Q(ram[3732]) );
  DFF ram_reg_1581__3_ ( .D(n7972), .CP(wclk), .Q(ram[3731]) );
  DFF ram_reg_1581__2_ ( .D(n7971), .CP(wclk), .Q(ram[3730]) );
  DFF ram_reg_1581__1_ ( .D(n7970), .CP(wclk), .Q(ram[3729]) );
  DFF ram_reg_1581__0_ ( .D(n7969), .CP(wclk), .Q(ram[3728]) );
  DFF ram_reg_1585__7_ ( .D(n7944), .CP(wclk), .Q(ram[3703]) );
  DFF ram_reg_1585__6_ ( .D(n7943), .CP(wclk), .Q(ram[3702]) );
  DFF ram_reg_1585__5_ ( .D(n7942), .CP(wclk), .Q(ram[3701]) );
  DFF ram_reg_1585__4_ ( .D(n7941), .CP(wclk), .Q(ram[3700]) );
  DFF ram_reg_1585__3_ ( .D(n7940), .CP(wclk), .Q(ram[3699]) );
  DFF ram_reg_1585__2_ ( .D(n7939), .CP(wclk), .Q(ram[3698]) );
  DFF ram_reg_1585__1_ ( .D(n7938), .CP(wclk), .Q(ram[3697]) );
  DFF ram_reg_1585__0_ ( .D(n7937), .CP(wclk), .Q(ram[3696]) );
  DFF ram_reg_1593__7_ ( .D(n7880), .CP(wclk), .Q(ram[3639]) );
  DFF ram_reg_1593__6_ ( .D(n7879), .CP(wclk), .Q(ram[3638]) );
  DFF ram_reg_1593__5_ ( .D(n7878), .CP(wclk), .Q(ram[3637]) );
  DFF ram_reg_1593__4_ ( .D(n7877), .CP(wclk), .Q(ram[3636]) );
  DFF ram_reg_1593__3_ ( .D(n7876), .CP(wclk), .Q(ram[3635]) );
  DFF ram_reg_1593__2_ ( .D(n7875), .CP(wclk), .Q(ram[3634]) );
  DFF ram_reg_1593__1_ ( .D(n7874), .CP(wclk), .Q(ram[3633]) );
  DFF ram_reg_1593__0_ ( .D(n7873), .CP(wclk), .Q(ram[3632]) );
  DFF ram_reg_1597__7_ ( .D(n7848), .CP(wclk), .Q(ram[3607]) );
  DFF ram_reg_1597__6_ ( .D(n7847), .CP(wclk), .Q(ram[3606]) );
  DFF ram_reg_1597__5_ ( .D(n7846), .CP(wclk), .Q(ram[3605]) );
  DFF ram_reg_1597__4_ ( .D(n7845), .CP(wclk), .Q(ram[3604]) );
  DFF ram_reg_1597__3_ ( .D(n7844), .CP(wclk), .Q(ram[3603]) );
  DFF ram_reg_1597__2_ ( .D(n7843), .CP(wclk), .Q(ram[3602]) );
  DFF ram_reg_1597__1_ ( .D(n7842), .CP(wclk), .Q(ram[3601]) );
  DFF ram_reg_1597__0_ ( .D(n7841), .CP(wclk), .Q(ram[3600]) );
  DFF ram_reg_1641__7_ ( .D(n7496), .CP(wclk), .Q(ram[3255]) );
  DFF ram_reg_1641__6_ ( .D(n7495), .CP(wclk), .Q(ram[3254]) );
  DFF ram_reg_1641__5_ ( .D(n7494), .CP(wclk), .Q(ram[3253]) );
  DFF ram_reg_1641__4_ ( .D(n7493), .CP(wclk), .Q(ram[3252]) );
  DFF ram_reg_1641__3_ ( .D(n7492), .CP(wclk), .Q(ram[3251]) );
  DFF ram_reg_1641__2_ ( .D(n7491), .CP(wclk), .Q(ram[3250]) );
  DFF ram_reg_1641__1_ ( .D(n7490), .CP(wclk), .Q(ram[3249]) );
  DFF ram_reg_1641__0_ ( .D(n7489), .CP(wclk), .Q(ram[3248]) );
  DFF ram_reg_1657__7_ ( .D(n7368), .CP(wclk), .Q(ram[3127]) );
  DFF ram_reg_1657__6_ ( .D(n7367), .CP(wclk), .Q(ram[3126]) );
  DFF ram_reg_1657__5_ ( .D(n7366), .CP(wclk), .Q(ram[3125]) );
  DFF ram_reg_1657__4_ ( .D(n7365), .CP(wclk), .Q(ram[3124]) );
  DFF ram_reg_1657__3_ ( .D(n7364), .CP(wclk), .Q(ram[3123]) );
  DFF ram_reg_1657__2_ ( .D(n7363), .CP(wclk), .Q(ram[3122]) );
  DFF ram_reg_1657__1_ ( .D(n7362), .CP(wclk), .Q(ram[3121]) );
  DFF ram_reg_1657__0_ ( .D(n7361), .CP(wclk), .Q(ram[3120]) );
  DFF ram_reg_1665__7_ ( .D(n7304), .CP(wclk), .Q(ram[3063]) );
  DFF ram_reg_1665__6_ ( .D(n7303), .CP(wclk), .Q(ram[3062]) );
  DFF ram_reg_1665__5_ ( .D(n7302), .CP(wclk), .Q(ram[3061]) );
  DFF ram_reg_1665__4_ ( .D(n7301), .CP(wclk), .Q(ram[3060]) );
  DFF ram_reg_1665__3_ ( .D(n7300), .CP(wclk), .Q(ram[3059]) );
  DFF ram_reg_1665__2_ ( .D(n7299), .CP(wclk), .Q(ram[3058]) );
  DFF ram_reg_1665__1_ ( .D(n7298), .CP(wclk), .Q(ram[3057]) );
  DFF ram_reg_1665__0_ ( .D(n7297), .CP(wclk), .Q(ram[3056]) );
  DFF ram_reg_1673__7_ ( .D(n7240), .CP(wclk), .Q(ram[2999]) );
  DFF ram_reg_1673__6_ ( .D(n7239), .CP(wclk), .Q(ram[2998]) );
  DFF ram_reg_1673__5_ ( .D(n7238), .CP(wclk), .Q(ram[2997]) );
  DFF ram_reg_1673__4_ ( .D(n7237), .CP(wclk), .Q(ram[2996]) );
  DFF ram_reg_1673__3_ ( .D(n7236), .CP(wclk), .Q(ram[2995]) );
  DFF ram_reg_1673__2_ ( .D(n7235), .CP(wclk), .Q(ram[2994]) );
  DFF ram_reg_1673__1_ ( .D(n7234), .CP(wclk), .Q(ram[2993]) );
  DFF ram_reg_1673__0_ ( .D(n7233), .CP(wclk), .Q(ram[2992]) );
  DFF ram_reg_1677__7_ ( .D(n7208), .CP(wclk), .Q(ram[2967]) );
  DFF ram_reg_1677__6_ ( .D(n7207), .CP(wclk), .Q(ram[2966]) );
  DFF ram_reg_1677__5_ ( .D(n7206), .CP(wclk), .Q(ram[2965]) );
  DFF ram_reg_1677__4_ ( .D(n7205), .CP(wclk), .Q(ram[2964]) );
  DFF ram_reg_1677__3_ ( .D(n7204), .CP(wclk), .Q(ram[2963]) );
  DFF ram_reg_1677__2_ ( .D(n7203), .CP(wclk), .Q(ram[2962]) );
  DFF ram_reg_1677__1_ ( .D(n7202), .CP(wclk), .Q(ram[2961]) );
  DFF ram_reg_1677__0_ ( .D(n7201), .CP(wclk), .Q(ram[2960]) );
  DFF ram_reg_1681__7_ ( .D(n7176), .CP(wclk), .Q(ram[2935]) );
  DFF ram_reg_1681__6_ ( .D(n7175), .CP(wclk), .Q(ram[2934]) );
  DFF ram_reg_1681__5_ ( .D(n7174), .CP(wclk), .Q(ram[2933]) );
  DFF ram_reg_1681__4_ ( .D(n7173), .CP(wclk), .Q(ram[2932]) );
  DFF ram_reg_1681__3_ ( .D(n7172), .CP(wclk), .Q(ram[2931]) );
  DFF ram_reg_1681__2_ ( .D(n7171), .CP(wclk), .Q(ram[2930]) );
  DFF ram_reg_1681__1_ ( .D(n7170), .CP(wclk), .Q(ram[2929]) );
  DFF ram_reg_1681__0_ ( .D(n7169), .CP(wclk), .Q(ram[2928]) );
  DFF ram_reg_1689__7_ ( .D(n7112), .CP(wclk), .Q(ram[2871]) );
  DFF ram_reg_1689__6_ ( .D(n7111), .CP(wclk), .Q(ram[2870]) );
  DFF ram_reg_1689__5_ ( .D(n7110), .CP(wclk), .Q(ram[2869]) );
  DFF ram_reg_1689__4_ ( .D(n7109), .CP(wclk), .Q(ram[2868]) );
  DFF ram_reg_1689__3_ ( .D(n7108), .CP(wclk), .Q(ram[2867]) );
  DFF ram_reg_1689__2_ ( .D(n7107), .CP(wclk), .Q(ram[2866]) );
  DFF ram_reg_1689__1_ ( .D(n7106), .CP(wclk), .Q(ram[2865]) );
  DFF ram_reg_1689__0_ ( .D(n7105), .CP(wclk), .Q(ram[2864]) );
  DFF ram_reg_1693__7_ ( .D(n7080), .CP(wclk), .Q(ram[2839]) );
  DFF ram_reg_1693__6_ ( .D(n7079), .CP(wclk), .Q(ram[2838]) );
  DFF ram_reg_1693__5_ ( .D(n7078), .CP(wclk), .Q(ram[2837]) );
  DFF ram_reg_1693__4_ ( .D(n7077), .CP(wclk), .Q(ram[2836]) );
  DFF ram_reg_1693__3_ ( .D(n7076), .CP(wclk), .Q(ram[2835]) );
  DFF ram_reg_1693__2_ ( .D(n7075), .CP(wclk), .Q(ram[2834]) );
  DFF ram_reg_1693__1_ ( .D(n7074), .CP(wclk), .Q(ram[2833]) );
  DFF ram_reg_1693__0_ ( .D(n7073), .CP(wclk), .Q(ram[2832]) );
  DFF ram_reg_1697__7_ ( .D(n7048), .CP(wclk), .Q(ram[2807]) );
  DFF ram_reg_1697__6_ ( .D(n7047), .CP(wclk), .Q(ram[2806]) );
  DFF ram_reg_1697__5_ ( .D(n7046), .CP(wclk), .Q(ram[2805]) );
  DFF ram_reg_1697__4_ ( .D(n7045), .CP(wclk), .Q(ram[2804]) );
  DFF ram_reg_1697__3_ ( .D(n7044), .CP(wclk), .Q(ram[2803]) );
  DFF ram_reg_1697__2_ ( .D(n7043), .CP(wclk), .Q(ram[2802]) );
  DFF ram_reg_1697__1_ ( .D(n7042), .CP(wclk), .Q(ram[2801]) );
  DFF ram_reg_1697__0_ ( .D(n7041), .CP(wclk), .Q(ram[2800]) );
  DFF ram_reg_1701__7_ ( .D(n7016), .CP(wclk), .Q(ram[2775]) );
  DFF ram_reg_1701__6_ ( .D(n7015), .CP(wclk), .Q(ram[2774]) );
  DFF ram_reg_1701__5_ ( .D(n7014), .CP(wclk), .Q(ram[2773]) );
  DFF ram_reg_1701__4_ ( .D(n7013), .CP(wclk), .Q(ram[2772]) );
  DFF ram_reg_1701__3_ ( .D(n7012), .CP(wclk), .Q(ram[2771]) );
  DFF ram_reg_1701__2_ ( .D(n7011), .CP(wclk), .Q(ram[2770]) );
  DFF ram_reg_1701__1_ ( .D(n7010), .CP(wclk), .Q(ram[2769]) );
  DFF ram_reg_1701__0_ ( .D(n7009), .CP(wclk), .Q(ram[2768]) );
  DFF ram_reg_1705__7_ ( .D(n6984), .CP(wclk), .Q(ram[2743]) );
  DFF ram_reg_1705__6_ ( .D(n6983), .CP(wclk), .Q(ram[2742]) );
  DFF ram_reg_1705__5_ ( .D(n6982), .CP(wclk), .Q(ram[2741]) );
  DFF ram_reg_1705__4_ ( .D(n6981), .CP(wclk), .Q(ram[2740]) );
  DFF ram_reg_1705__3_ ( .D(n6980), .CP(wclk), .Q(ram[2739]) );
  DFF ram_reg_1705__2_ ( .D(n6979), .CP(wclk), .Q(ram[2738]) );
  DFF ram_reg_1705__1_ ( .D(n6978), .CP(wclk), .Q(ram[2737]) );
  DFF ram_reg_1705__0_ ( .D(n6977), .CP(wclk), .Q(ram[2736]) );
  DFF ram_reg_1709__7_ ( .D(n6952), .CP(wclk), .Q(ram[2711]) );
  DFF ram_reg_1709__6_ ( .D(n6951), .CP(wclk), .Q(ram[2710]) );
  DFF ram_reg_1709__5_ ( .D(n6950), .CP(wclk), .Q(ram[2709]) );
  DFF ram_reg_1709__4_ ( .D(n6949), .CP(wclk), .Q(ram[2708]) );
  DFF ram_reg_1709__3_ ( .D(n6948), .CP(wclk), .Q(ram[2707]) );
  DFF ram_reg_1709__2_ ( .D(n6947), .CP(wclk), .Q(ram[2706]) );
  DFF ram_reg_1709__1_ ( .D(n6946), .CP(wclk), .Q(ram[2705]) );
  DFF ram_reg_1709__0_ ( .D(n6945), .CP(wclk), .Q(ram[2704]) );
  DFF ram_reg_1713__7_ ( .D(n6920), .CP(wclk), .Q(ram[2679]) );
  DFF ram_reg_1713__6_ ( .D(n6919), .CP(wclk), .Q(ram[2678]) );
  DFF ram_reg_1713__5_ ( .D(n6918), .CP(wclk), .Q(ram[2677]) );
  DFF ram_reg_1713__4_ ( .D(n6917), .CP(wclk), .Q(ram[2676]) );
  DFF ram_reg_1713__3_ ( .D(n6916), .CP(wclk), .Q(ram[2675]) );
  DFF ram_reg_1713__2_ ( .D(n6915), .CP(wclk), .Q(ram[2674]) );
  DFF ram_reg_1713__1_ ( .D(n6914), .CP(wclk), .Q(ram[2673]) );
  DFF ram_reg_1713__0_ ( .D(n6913), .CP(wclk), .Q(ram[2672]) );
  DFF ram_reg_1717__7_ ( .D(n6888), .CP(wclk), .Q(ram[2647]) );
  DFF ram_reg_1717__6_ ( .D(n6887), .CP(wclk), .Q(ram[2646]) );
  DFF ram_reg_1717__5_ ( .D(n6886), .CP(wclk), .Q(ram[2645]) );
  DFF ram_reg_1717__4_ ( .D(n6885), .CP(wclk), .Q(ram[2644]) );
  DFF ram_reg_1717__3_ ( .D(n6884), .CP(wclk), .Q(ram[2643]) );
  DFF ram_reg_1717__2_ ( .D(n6883), .CP(wclk), .Q(ram[2642]) );
  DFF ram_reg_1717__1_ ( .D(n6882), .CP(wclk), .Q(ram[2641]) );
  DFF ram_reg_1717__0_ ( .D(n6881), .CP(wclk), .Q(ram[2640]) );
  DFF ram_reg_1721__7_ ( .D(n6856), .CP(wclk), .Q(ram[2615]) );
  DFF ram_reg_1721__6_ ( .D(n6855), .CP(wclk), .Q(ram[2614]) );
  DFF ram_reg_1721__5_ ( .D(n6854), .CP(wclk), .Q(ram[2613]) );
  DFF ram_reg_1721__4_ ( .D(n6853), .CP(wclk), .Q(ram[2612]) );
  DFF ram_reg_1721__3_ ( .D(n6852), .CP(wclk), .Q(ram[2611]) );
  DFF ram_reg_1721__2_ ( .D(n6851), .CP(wclk), .Q(ram[2610]) );
  DFF ram_reg_1721__1_ ( .D(n6850), .CP(wclk), .Q(ram[2609]) );
  DFF ram_reg_1721__0_ ( .D(n6849), .CP(wclk), .Q(ram[2608]) );
  DFF ram_reg_1725__7_ ( .D(n6824), .CP(wclk), .Q(ram[2583]) );
  DFF ram_reg_1725__6_ ( .D(n6823), .CP(wclk), .Q(ram[2582]) );
  DFF ram_reg_1725__5_ ( .D(n6822), .CP(wclk), .Q(ram[2581]) );
  DFF ram_reg_1725__4_ ( .D(n6821), .CP(wclk), .Q(ram[2580]) );
  DFF ram_reg_1725__3_ ( .D(n6820), .CP(wclk), .Q(ram[2579]) );
  DFF ram_reg_1725__2_ ( .D(n6819), .CP(wclk), .Q(ram[2578]) );
  DFF ram_reg_1725__1_ ( .D(n6818), .CP(wclk), .Q(ram[2577]) );
  DFF ram_reg_1725__0_ ( .D(n6817), .CP(wclk), .Q(ram[2576]) );
  DFF ram_reg_1729__7_ ( .D(n6792), .CP(wclk), .Q(ram[2551]) );
  DFF ram_reg_1729__6_ ( .D(n6791), .CP(wclk), .Q(ram[2550]) );
  DFF ram_reg_1729__5_ ( .D(n6790), .CP(wclk), .Q(ram[2549]) );
  DFF ram_reg_1729__4_ ( .D(n6789), .CP(wclk), .Q(ram[2548]) );
  DFF ram_reg_1729__3_ ( .D(n6788), .CP(wclk), .Q(ram[2547]) );
  DFF ram_reg_1729__2_ ( .D(n6787), .CP(wclk), .Q(ram[2546]) );
  DFF ram_reg_1729__1_ ( .D(n6786), .CP(wclk), .Q(ram[2545]) );
  DFF ram_reg_1729__0_ ( .D(n6785), .CP(wclk), .Q(ram[2544]) );
  DFF ram_reg_1737__7_ ( .D(n6728), .CP(wclk), .Q(ram[2487]) );
  DFF ram_reg_1737__6_ ( .D(n6727), .CP(wclk), .Q(ram[2486]) );
  DFF ram_reg_1737__5_ ( .D(n6726), .CP(wclk), .Q(ram[2485]) );
  DFF ram_reg_1737__4_ ( .D(n6725), .CP(wclk), .Q(ram[2484]) );
  DFF ram_reg_1737__3_ ( .D(n6724), .CP(wclk), .Q(ram[2483]) );
  DFF ram_reg_1737__2_ ( .D(n6723), .CP(wclk), .Q(ram[2482]) );
  DFF ram_reg_1737__1_ ( .D(n6722), .CP(wclk), .Q(ram[2481]) );
  DFF ram_reg_1737__0_ ( .D(n6721), .CP(wclk), .Q(ram[2480]) );
  DFF ram_reg_1741__7_ ( .D(n6696), .CP(wclk), .Q(ram[2455]) );
  DFF ram_reg_1741__6_ ( .D(n6695), .CP(wclk), .Q(ram[2454]) );
  DFF ram_reg_1741__5_ ( .D(n6694), .CP(wclk), .Q(ram[2453]) );
  DFF ram_reg_1741__4_ ( .D(n6693), .CP(wclk), .Q(ram[2452]) );
  DFF ram_reg_1741__3_ ( .D(n6692), .CP(wclk), .Q(ram[2451]) );
  DFF ram_reg_1741__2_ ( .D(n6691), .CP(wclk), .Q(ram[2450]) );
  DFF ram_reg_1741__1_ ( .D(n6690), .CP(wclk), .Q(ram[2449]) );
  DFF ram_reg_1741__0_ ( .D(n6689), .CP(wclk), .Q(ram[2448]) );
  DFF ram_reg_1753__7_ ( .D(n6600), .CP(wclk), .Q(ram[2359]) );
  DFF ram_reg_1753__6_ ( .D(n6599), .CP(wclk), .Q(ram[2358]) );
  DFF ram_reg_1753__5_ ( .D(n6598), .CP(wclk), .Q(ram[2357]) );
  DFF ram_reg_1753__4_ ( .D(n6597), .CP(wclk), .Q(ram[2356]) );
  DFF ram_reg_1753__3_ ( .D(n6596), .CP(wclk), .Q(ram[2355]) );
  DFF ram_reg_1753__2_ ( .D(n6595), .CP(wclk), .Q(ram[2354]) );
  DFF ram_reg_1753__1_ ( .D(n6594), .CP(wclk), .Q(ram[2353]) );
  DFF ram_reg_1753__0_ ( .D(n6593), .CP(wclk), .Q(ram[2352]) );
  DFF ram_reg_1757__7_ ( .D(n6568), .CP(wclk), .Q(ram[2327]) );
  DFF ram_reg_1757__6_ ( .D(n6567), .CP(wclk), .Q(ram[2326]) );
  DFF ram_reg_1757__5_ ( .D(n6566), .CP(wclk), .Q(ram[2325]) );
  DFF ram_reg_1757__4_ ( .D(n6565), .CP(wclk), .Q(ram[2324]) );
  DFF ram_reg_1757__3_ ( .D(n6564), .CP(wclk), .Q(ram[2323]) );
  DFF ram_reg_1757__2_ ( .D(n6563), .CP(wclk), .Q(ram[2322]) );
  DFF ram_reg_1757__1_ ( .D(n6562), .CP(wclk), .Q(ram[2321]) );
  DFF ram_reg_1757__0_ ( .D(n6561), .CP(wclk), .Q(ram[2320]) );
  DFF ram_reg_1761__7_ ( .D(n6536), .CP(wclk), .Q(ram[2295]) );
  DFF ram_reg_1761__6_ ( .D(n6535), .CP(wclk), .Q(ram[2294]) );
  DFF ram_reg_1761__5_ ( .D(n6534), .CP(wclk), .Q(ram[2293]) );
  DFF ram_reg_1761__4_ ( .D(n6533), .CP(wclk), .Q(ram[2292]) );
  DFF ram_reg_1761__3_ ( .D(n6532), .CP(wclk), .Q(ram[2291]) );
  DFF ram_reg_1761__2_ ( .D(n6531), .CP(wclk), .Q(ram[2290]) );
  DFF ram_reg_1761__1_ ( .D(n6530), .CP(wclk), .Q(ram[2289]) );
  DFF ram_reg_1761__0_ ( .D(n6529), .CP(wclk), .Q(ram[2288]) );
  DFF ram_reg_1769__7_ ( .D(n6472), .CP(wclk), .Q(ram[2231]) );
  DFF ram_reg_1769__6_ ( .D(n6471), .CP(wclk), .Q(ram[2230]) );
  DFF ram_reg_1769__5_ ( .D(n6470), .CP(wclk), .Q(ram[2229]) );
  DFF ram_reg_1769__4_ ( .D(n6469), .CP(wclk), .Q(ram[2228]) );
  DFF ram_reg_1769__3_ ( .D(n6468), .CP(wclk), .Q(ram[2227]) );
  DFF ram_reg_1769__2_ ( .D(n6467), .CP(wclk), .Q(ram[2226]) );
  DFF ram_reg_1769__1_ ( .D(n6466), .CP(wclk), .Q(ram[2225]) );
  DFF ram_reg_1769__0_ ( .D(n6465), .CP(wclk), .Q(ram[2224]) );
  DFF ram_reg_1773__7_ ( .D(n6440), .CP(wclk), .Q(ram[2199]) );
  DFF ram_reg_1773__6_ ( .D(n6439), .CP(wclk), .Q(ram[2198]) );
  DFF ram_reg_1773__5_ ( .D(n6438), .CP(wclk), .Q(ram[2197]) );
  DFF ram_reg_1773__4_ ( .D(n6437), .CP(wclk), .Q(ram[2196]) );
  DFF ram_reg_1773__3_ ( .D(n6436), .CP(wclk), .Q(ram[2195]) );
  DFF ram_reg_1773__2_ ( .D(n6435), .CP(wclk), .Q(ram[2194]) );
  DFF ram_reg_1773__1_ ( .D(n6434), .CP(wclk), .Q(ram[2193]) );
  DFF ram_reg_1773__0_ ( .D(n6433), .CP(wclk), .Q(ram[2192]) );
  DFF ram_reg_1777__7_ ( .D(n6408), .CP(wclk), .Q(ram[2167]) );
  DFF ram_reg_1777__6_ ( .D(n6407), .CP(wclk), .Q(ram[2166]) );
  DFF ram_reg_1777__5_ ( .D(n6406), .CP(wclk), .Q(ram[2165]) );
  DFF ram_reg_1777__4_ ( .D(n6405), .CP(wclk), .Q(ram[2164]) );
  DFF ram_reg_1777__3_ ( .D(n6404), .CP(wclk), .Q(ram[2163]) );
  DFF ram_reg_1777__2_ ( .D(n6403), .CP(wclk), .Q(ram[2162]) );
  DFF ram_reg_1777__1_ ( .D(n6402), .CP(wclk), .Q(ram[2161]) );
  DFF ram_reg_1777__0_ ( .D(n6401), .CP(wclk), .Q(ram[2160]) );
  DFF ram_reg_1785__7_ ( .D(n6344), .CP(wclk), .Q(ram[2103]) );
  DFF ram_reg_1785__6_ ( .D(n6343), .CP(wclk), .Q(ram[2102]) );
  DFF ram_reg_1785__5_ ( .D(n6342), .CP(wclk), .Q(ram[2101]) );
  DFF ram_reg_1785__4_ ( .D(n6341), .CP(wclk), .Q(ram[2100]) );
  DFF ram_reg_1785__3_ ( .D(n6340), .CP(wclk), .Q(ram[2099]) );
  DFF ram_reg_1785__2_ ( .D(n6339), .CP(wclk), .Q(ram[2098]) );
  DFF ram_reg_1785__1_ ( .D(n6338), .CP(wclk), .Q(ram[2097]) );
  DFF ram_reg_1785__0_ ( .D(n6337), .CP(wclk), .Q(ram[2096]) );
  DFF ram_reg_1789__7_ ( .D(n6312), .CP(wclk), .Q(ram[2071]) );
  DFF ram_reg_1789__6_ ( .D(n6311), .CP(wclk), .Q(ram[2070]) );
  DFF ram_reg_1789__5_ ( .D(n6310), .CP(wclk), .Q(ram[2069]) );
  DFF ram_reg_1789__4_ ( .D(n6309), .CP(wclk), .Q(ram[2068]) );
  DFF ram_reg_1789__3_ ( .D(n6308), .CP(wclk), .Q(ram[2067]) );
  DFF ram_reg_1789__2_ ( .D(n6307), .CP(wclk), .Q(ram[2066]) );
  DFF ram_reg_1789__1_ ( .D(n6306), .CP(wclk), .Q(ram[2065]) );
  DFF ram_reg_1789__0_ ( .D(n6305), .CP(wclk), .Q(ram[2064]) );
  DFF ram_reg_1801__7_ ( .D(n6216), .CP(wclk), .Q(ram[1975]) );
  DFF ram_reg_1801__6_ ( .D(n6215), .CP(wclk), .Q(ram[1974]) );
  DFF ram_reg_1801__5_ ( .D(n6214), .CP(wclk), .Q(ram[1973]) );
  DFF ram_reg_1801__4_ ( .D(n6213), .CP(wclk), .Q(ram[1972]) );
  DFF ram_reg_1801__3_ ( .D(n6212), .CP(wclk), .Q(ram[1971]) );
  DFF ram_reg_1801__2_ ( .D(n6211), .CP(wclk), .Q(ram[1970]) );
  DFF ram_reg_1801__1_ ( .D(n6210), .CP(wclk), .Q(ram[1969]) );
  DFF ram_reg_1801__0_ ( .D(n6209), .CP(wclk), .Q(ram[1968]) );
  DFF ram_reg_1805__7_ ( .D(n6184), .CP(wclk), .Q(ram[1943]) );
  DFF ram_reg_1805__6_ ( .D(n6183), .CP(wclk), .Q(ram[1942]) );
  DFF ram_reg_1805__5_ ( .D(n6182), .CP(wclk), .Q(ram[1941]) );
  DFF ram_reg_1805__4_ ( .D(n6181), .CP(wclk), .Q(ram[1940]) );
  DFF ram_reg_1805__3_ ( .D(n6180), .CP(wclk), .Q(ram[1939]) );
  DFF ram_reg_1805__2_ ( .D(n6179), .CP(wclk), .Q(ram[1938]) );
  DFF ram_reg_1805__1_ ( .D(n6178), .CP(wclk), .Q(ram[1937]) );
  DFF ram_reg_1805__0_ ( .D(n6177), .CP(wclk), .Q(ram[1936]) );
  DFF ram_reg_1817__7_ ( .D(n6088), .CP(wclk), .Q(ram[1847]) );
  DFF ram_reg_1817__6_ ( .D(n6087), .CP(wclk), .Q(ram[1846]) );
  DFF ram_reg_1817__5_ ( .D(n6086), .CP(wclk), .Q(ram[1845]) );
  DFF ram_reg_1817__4_ ( .D(n6085), .CP(wclk), .Q(ram[1844]) );
  DFF ram_reg_1817__3_ ( .D(n6084), .CP(wclk), .Q(ram[1843]) );
  DFF ram_reg_1817__2_ ( .D(n6083), .CP(wclk), .Q(ram[1842]) );
  DFF ram_reg_1817__1_ ( .D(n6082), .CP(wclk), .Q(ram[1841]) );
  DFF ram_reg_1817__0_ ( .D(n6081), .CP(wclk), .Q(ram[1840]) );
  DFF ram_reg_1825__7_ ( .D(n6024), .CP(wclk), .Q(ram[1783]) );
  DFF ram_reg_1825__6_ ( .D(n6023), .CP(wclk), .Q(ram[1782]) );
  DFF ram_reg_1825__5_ ( .D(n6022), .CP(wclk), .Q(ram[1781]) );
  DFF ram_reg_1825__4_ ( .D(n6021), .CP(wclk), .Q(ram[1780]) );
  DFF ram_reg_1825__3_ ( .D(n6020), .CP(wclk), .Q(ram[1779]) );
  DFF ram_reg_1825__2_ ( .D(n6019), .CP(wclk), .Q(ram[1778]) );
  DFF ram_reg_1825__1_ ( .D(n6018), .CP(wclk), .Q(ram[1777]) );
  DFF ram_reg_1825__0_ ( .D(n6017), .CP(wclk), .Q(ram[1776]) );
  DFF ram_reg_1833__7_ ( .D(n5960), .CP(wclk), .Q(ram[1719]) );
  DFF ram_reg_1833__6_ ( .D(n5959), .CP(wclk), .Q(ram[1718]) );
  DFF ram_reg_1833__5_ ( .D(n5958), .CP(wclk), .Q(ram[1717]) );
  DFF ram_reg_1833__4_ ( .D(n5957), .CP(wclk), .Q(ram[1716]) );
  DFF ram_reg_1833__3_ ( .D(n5956), .CP(wclk), .Q(ram[1715]) );
  DFF ram_reg_1833__2_ ( .D(n5955), .CP(wclk), .Q(ram[1714]) );
  DFF ram_reg_1833__1_ ( .D(n5954), .CP(wclk), .Q(ram[1713]) );
  DFF ram_reg_1833__0_ ( .D(n5953), .CP(wclk), .Q(ram[1712]) );
  DFF ram_reg_1837__7_ ( .D(n5928), .CP(wclk), .Q(ram[1687]) );
  DFF ram_reg_1837__6_ ( .D(n5927), .CP(wclk), .Q(ram[1686]) );
  DFF ram_reg_1837__5_ ( .D(n5926), .CP(wclk), .Q(ram[1685]) );
  DFF ram_reg_1837__4_ ( .D(n5925), .CP(wclk), .Q(ram[1684]) );
  DFF ram_reg_1837__3_ ( .D(n5924), .CP(wclk), .Q(ram[1683]) );
  DFF ram_reg_1837__2_ ( .D(n5923), .CP(wclk), .Q(ram[1682]) );
  DFF ram_reg_1837__1_ ( .D(n5922), .CP(wclk), .Q(ram[1681]) );
  DFF ram_reg_1837__0_ ( .D(n5921), .CP(wclk), .Q(ram[1680]) );
  DFF ram_reg_1841__7_ ( .D(n5896), .CP(wclk), .Q(ram[1655]) );
  DFF ram_reg_1841__6_ ( .D(n5895), .CP(wclk), .Q(ram[1654]) );
  DFF ram_reg_1841__5_ ( .D(n5894), .CP(wclk), .Q(ram[1653]) );
  DFF ram_reg_1841__4_ ( .D(n5893), .CP(wclk), .Q(ram[1652]) );
  DFF ram_reg_1841__3_ ( .D(n5892), .CP(wclk), .Q(ram[1651]) );
  DFF ram_reg_1841__2_ ( .D(n5891), .CP(wclk), .Q(ram[1650]) );
  DFF ram_reg_1841__1_ ( .D(n5890), .CP(wclk), .Q(ram[1649]) );
  DFF ram_reg_1841__0_ ( .D(n5889), .CP(wclk), .Q(ram[1648]) );
  DFF ram_reg_1849__7_ ( .D(n5832), .CP(wclk), .Q(ram[1591]) );
  DFF ram_reg_1849__6_ ( .D(n5831), .CP(wclk), .Q(ram[1590]) );
  DFF ram_reg_1849__5_ ( .D(n5830), .CP(wclk), .Q(ram[1589]) );
  DFF ram_reg_1849__4_ ( .D(n5829), .CP(wclk), .Q(ram[1588]) );
  DFF ram_reg_1849__3_ ( .D(n5828), .CP(wclk), .Q(ram[1587]) );
  DFF ram_reg_1849__2_ ( .D(n5827), .CP(wclk), .Q(ram[1586]) );
  DFF ram_reg_1849__1_ ( .D(n5826), .CP(wclk), .Q(ram[1585]) );
  DFF ram_reg_1849__0_ ( .D(n5825), .CP(wclk), .Q(ram[1584]) );
  DFF ram_reg_1853__7_ ( .D(n5800), .CP(wclk), .Q(ram[1559]) );
  DFF ram_reg_1853__6_ ( .D(n5799), .CP(wclk), .Q(ram[1558]) );
  DFF ram_reg_1853__5_ ( .D(n5798), .CP(wclk), .Q(ram[1557]) );
  DFF ram_reg_1853__4_ ( .D(n5797), .CP(wclk), .Q(ram[1556]) );
  DFF ram_reg_1853__3_ ( .D(n5796), .CP(wclk), .Q(ram[1555]) );
  DFF ram_reg_1853__2_ ( .D(n5795), .CP(wclk), .Q(ram[1554]) );
  DFF ram_reg_1853__1_ ( .D(n5794), .CP(wclk), .Q(ram[1553]) );
  DFF ram_reg_1853__0_ ( .D(n5793), .CP(wclk), .Q(ram[1552]) );
  DFF ram_reg_1897__7_ ( .D(n5448), .CP(wclk), .Q(ram[1207]) );
  DFF ram_reg_1897__6_ ( .D(n5447), .CP(wclk), .Q(ram[1206]) );
  DFF ram_reg_1897__5_ ( .D(n5446), .CP(wclk), .Q(ram[1205]) );
  DFF ram_reg_1897__4_ ( .D(n5445), .CP(wclk), .Q(ram[1204]) );
  DFF ram_reg_1897__3_ ( .D(n5444), .CP(wclk), .Q(ram[1203]) );
  DFF ram_reg_1897__2_ ( .D(n5443), .CP(wclk), .Q(ram[1202]) );
  DFF ram_reg_1897__1_ ( .D(n5442), .CP(wclk), .Q(ram[1201]) );
  DFF ram_reg_1897__0_ ( .D(n5441), .CP(wclk), .Q(ram[1200]) );
  DFF ram_reg_1913__7_ ( .D(n5320), .CP(wclk), .Q(ram[1079]) );
  DFF ram_reg_1913__6_ ( .D(n5319), .CP(wclk), .Q(ram[1078]) );
  DFF ram_reg_1913__5_ ( .D(n5318), .CP(wclk), .Q(ram[1077]) );
  DFF ram_reg_1913__4_ ( .D(n5317), .CP(wclk), .Q(ram[1076]) );
  DFF ram_reg_1913__3_ ( .D(n5316), .CP(wclk), .Q(ram[1075]) );
  DFF ram_reg_1913__2_ ( .D(n5315), .CP(wclk), .Q(ram[1074]) );
  DFF ram_reg_1913__1_ ( .D(n5314), .CP(wclk), .Q(ram[1073]) );
  DFF ram_reg_1913__0_ ( .D(n5313), .CP(wclk), .Q(ram[1072]) );
  DFF ram_reg_1917__7_ ( .D(n5288), .CP(wclk), .Q(ram[1047]) );
  DFF ram_reg_1917__6_ ( .D(n5287), .CP(wclk), .Q(ram[1046]) );
  DFF ram_reg_1917__5_ ( .D(n5286), .CP(wclk), .Q(ram[1045]) );
  DFF ram_reg_1917__4_ ( .D(n5285), .CP(wclk), .Q(ram[1044]) );
  DFF ram_reg_1917__3_ ( .D(n5284), .CP(wclk), .Q(ram[1043]) );
  DFF ram_reg_1917__2_ ( .D(n5283), .CP(wclk), .Q(ram[1042]) );
  DFF ram_reg_1917__1_ ( .D(n5282), .CP(wclk), .Q(ram[1041]) );
  DFF ram_reg_1917__0_ ( .D(n5281), .CP(wclk), .Q(ram[1040]) );
  DFF ram_reg_1921__7_ ( .D(n5256), .CP(wclk), .Q(ram[1015]) );
  DFF ram_reg_1921__6_ ( .D(n5255), .CP(wclk), .Q(ram[1014]) );
  DFF ram_reg_1921__5_ ( .D(n5254), .CP(wclk), .Q(ram[1013]) );
  DFF ram_reg_1921__4_ ( .D(n5253), .CP(wclk), .Q(ram[1012]) );
  DFF ram_reg_1921__3_ ( .D(n5252), .CP(wclk), .Q(ram[1011]) );
  DFF ram_reg_1921__2_ ( .D(n5251), .CP(wclk), .Q(ram[1010]) );
  DFF ram_reg_1921__1_ ( .D(n5250), .CP(wclk), .Q(ram[1009]) );
  DFF ram_reg_1921__0_ ( .D(n5249), .CP(wclk), .Q(ram[1008]) );
  DFF ram_reg_1929__7_ ( .D(n5192), .CP(wclk), .Q(ram[951]) );
  DFF ram_reg_1929__6_ ( .D(n5191), .CP(wclk), .Q(ram[950]) );
  DFF ram_reg_1929__5_ ( .D(n5190), .CP(wclk), .Q(ram[949]) );
  DFF ram_reg_1929__4_ ( .D(n5189), .CP(wclk), .Q(ram[948]) );
  DFF ram_reg_1929__3_ ( .D(n5188), .CP(wclk), .Q(ram[947]) );
  DFF ram_reg_1929__2_ ( .D(n5187), .CP(wclk), .Q(ram[946]) );
  DFF ram_reg_1929__1_ ( .D(n5186), .CP(wclk), .Q(ram[945]) );
  DFF ram_reg_1929__0_ ( .D(n5185), .CP(wclk), .Q(ram[944]) );
  DFF ram_reg_1933__7_ ( .D(n5160), .CP(wclk), .Q(ram[919]) );
  DFF ram_reg_1933__6_ ( .D(n5159), .CP(wclk), .Q(ram[918]) );
  DFF ram_reg_1933__5_ ( .D(n5158), .CP(wclk), .Q(ram[917]) );
  DFF ram_reg_1933__4_ ( .D(n5157), .CP(wclk), .Q(ram[916]) );
  DFF ram_reg_1933__3_ ( .D(n5156), .CP(wclk), .Q(ram[915]) );
  DFF ram_reg_1933__2_ ( .D(n5155), .CP(wclk), .Q(ram[914]) );
  DFF ram_reg_1933__1_ ( .D(n5154), .CP(wclk), .Q(ram[913]) );
  DFF ram_reg_1933__0_ ( .D(n5153), .CP(wclk), .Q(ram[912]) );
  DFF ram_reg_1937__7_ ( .D(n5128), .CP(wclk), .Q(ram[887]) );
  DFF ram_reg_1937__6_ ( .D(n5127), .CP(wclk), .Q(ram[886]) );
  DFF ram_reg_1937__5_ ( .D(n5126), .CP(wclk), .Q(ram[885]) );
  DFF ram_reg_1937__4_ ( .D(n5125), .CP(wclk), .Q(ram[884]) );
  DFF ram_reg_1937__3_ ( .D(n5124), .CP(wclk), .Q(ram[883]) );
  DFF ram_reg_1937__2_ ( .D(n5123), .CP(wclk), .Q(ram[882]) );
  DFF ram_reg_1937__1_ ( .D(n5122), .CP(wclk), .Q(ram[881]) );
  DFF ram_reg_1937__0_ ( .D(n5121), .CP(wclk), .Q(ram[880]) );
  DFF ram_reg_1945__7_ ( .D(n5064), .CP(wclk), .Q(ram[823]) );
  DFF ram_reg_1945__6_ ( .D(n5063), .CP(wclk), .Q(ram[822]) );
  DFF ram_reg_1945__5_ ( .D(n5062), .CP(wclk), .Q(ram[821]) );
  DFF ram_reg_1945__4_ ( .D(n5061), .CP(wclk), .Q(ram[820]) );
  DFF ram_reg_1945__3_ ( .D(n5060), .CP(wclk), .Q(ram[819]) );
  DFF ram_reg_1945__2_ ( .D(n5059), .CP(wclk), .Q(ram[818]) );
  DFF ram_reg_1945__1_ ( .D(n5058), .CP(wclk), .Q(ram[817]) );
  DFF ram_reg_1945__0_ ( .D(n5057), .CP(wclk), .Q(ram[816]) );
  DFF ram_reg_1949__7_ ( .D(n5032), .CP(wclk), .Q(ram[791]) );
  DFF ram_reg_1949__6_ ( .D(n5031), .CP(wclk), .Q(ram[790]) );
  DFF ram_reg_1949__5_ ( .D(n5030), .CP(wclk), .Q(ram[789]) );
  DFF ram_reg_1949__4_ ( .D(n5029), .CP(wclk), .Q(ram[788]) );
  DFF ram_reg_1949__3_ ( .D(n5028), .CP(wclk), .Q(ram[787]) );
  DFF ram_reg_1949__2_ ( .D(n5027), .CP(wclk), .Q(ram[786]) );
  DFF ram_reg_1949__1_ ( .D(n5026), .CP(wclk), .Q(ram[785]) );
  DFF ram_reg_1949__0_ ( .D(n5025), .CP(wclk), .Q(ram[784]) );
  DFF ram_reg_1953__7_ ( .D(n5000), .CP(wclk), .Q(ram[759]) );
  DFF ram_reg_1953__6_ ( .D(n4999), .CP(wclk), .Q(ram[758]) );
  DFF ram_reg_1953__5_ ( .D(n4998), .CP(wclk), .Q(ram[757]) );
  DFF ram_reg_1953__4_ ( .D(n4997), .CP(wclk), .Q(ram[756]) );
  DFF ram_reg_1953__3_ ( .D(n4996), .CP(wclk), .Q(ram[755]) );
  DFF ram_reg_1953__2_ ( .D(n4995), .CP(wclk), .Q(ram[754]) );
  DFF ram_reg_1953__1_ ( .D(n4994), .CP(wclk), .Q(ram[753]) );
  DFF ram_reg_1953__0_ ( .D(n4993), .CP(wclk), .Q(ram[752]) );
  DFF ram_reg_1957__7_ ( .D(n4968), .CP(wclk), .Q(ram[727]) );
  DFF ram_reg_1957__6_ ( .D(n4967), .CP(wclk), .Q(ram[726]) );
  DFF ram_reg_1957__5_ ( .D(n4966), .CP(wclk), .Q(ram[725]) );
  DFF ram_reg_1957__4_ ( .D(n4965), .CP(wclk), .Q(ram[724]) );
  DFF ram_reg_1957__3_ ( .D(n4964), .CP(wclk), .Q(ram[723]) );
  DFF ram_reg_1957__2_ ( .D(n4963), .CP(wclk), .Q(ram[722]) );
  DFF ram_reg_1957__1_ ( .D(n4962), .CP(wclk), .Q(ram[721]) );
  DFF ram_reg_1957__0_ ( .D(n4961), .CP(wclk), .Q(ram[720]) );
  DFF ram_reg_1961__7_ ( .D(n4936), .CP(wclk), .Q(ram[695]) );
  DFF ram_reg_1961__6_ ( .D(n4935), .CP(wclk), .Q(ram[694]) );
  DFF ram_reg_1961__5_ ( .D(n4934), .CP(wclk), .Q(ram[693]) );
  DFF ram_reg_1961__4_ ( .D(n4933), .CP(wclk), .Q(ram[692]) );
  DFF ram_reg_1961__3_ ( .D(n4932), .CP(wclk), .Q(ram[691]) );
  DFF ram_reg_1961__2_ ( .D(n4931), .CP(wclk), .Q(ram[690]) );
  DFF ram_reg_1961__1_ ( .D(n4930), .CP(wclk), .Q(ram[689]) );
  DFF ram_reg_1961__0_ ( .D(n4929), .CP(wclk), .Q(ram[688]) );
  DFF ram_reg_1965__7_ ( .D(n4904), .CP(wclk), .Q(ram[663]) );
  DFF ram_reg_1965__6_ ( .D(n4903), .CP(wclk), .Q(ram[662]) );
  DFF ram_reg_1965__5_ ( .D(n4902), .CP(wclk), .Q(ram[661]) );
  DFF ram_reg_1965__4_ ( .D(n4901), .CP(wclk), .Q(ram[660]) );
  DFF ram_reg_1965__3_ ( .D(n4900), .CP(wclk), .Q(ram[659]) );
  DFF ram_reg_1965__2_ ( .D(n4899), .CP(wclk), .Q(ram[658]) );
  DFF ram_reg_1965__1_ ( .D(n4898), .CP(wclk), .Q(ram[657]) );
  DFF ram_reg_1965__0_ ( .D(n4897), .CP(wclk), .Q(ram[656]) );
  DFF ram_reg_1969__7_ ( .D(n4872), .CP(wclk), .Q(ram[631]) );
  DFF ram_reg_1969__6_ ( .D(n4871), .CP(wclk), .Q(ram[630]) );
  DFF ram_reg_1969__5_ ( .D(n4870), .CP(wclk), .Q(ram[629]) );
  DFF ram_reg_1969__4_ ( .D(n4869), .CP(wclk), .Q(ram[628]) );
  DFF ram_reg_1969__3_ ( .D(n4868), .CP(wclk), .Q(ram[627]) );
  DFF ram_reg_1969__2_ ( .D(n4867), .CP(wclk), .Q(ram[626]) );
  DFF ram_reg_1969__1_ ( .D(n4866), .CP(wclk), .Q(ram[625]) );
  DFF ram_reg_1969__0_ ( .D(n4865), .CP(wclk), .Q(ram[624]) );
  DFF ram_reg_1973__7_ ( .D(n4840), .CP(wclk), .Q(ram[599]) );
  DFF ram_reg_1973__6_ ( .D(n4839), .CP(wclk), .Q(ram[598]) );
  DFF ram_reg_1973__5_ ( .D(n4838), .CP(wclk), .Q(ram[597]) );
  DFF ram_reg_1973__4_ ( .D(n4837), .CP(wclk), .Q(ram[596]) );
  DFF ram_reg_1973__3_ ( .D(n4836), .CP(wclk), .Q(ram[595]) );
  DFF ram_reg_1973__2_ ( .D(n4835), .CP(wclk), .Q(ram[594]) );
  DFF ram_reg_1973__1_ ( .D(n4834), .CP(wclk), .Q(ram[593]) );
  DFF ram_reg_1973__0_ ( .D(n4833), .CP(wclk), .Q(ram[592]) );
  DFF ram_reg_1977__7_ ( .D(n4808), .CP(wclk), .Q(ram[567]) );
  DFF ram_reg_1977__6_ ( .D(n4807), .CP(wclk), .Q(ram[566]) );
  DFF ram_reg_1977__5_ ( .D(n4806), .CP(wclk), .Q(ram[565]) );
  DFF ram_reg_1977__4_ ( .D(n4805), .CP(wclk), .Q(ram[564]) );
  DFF ram_reg_1977__3_ ( .D(n4804), .CP(wclk), .Q(ram[563]) );
  DFF ram_reg_1977__2_ ( .D(n4803), .CP(wclk), .Q(ram[562]) );
  DFF ram_reg_1977__1_ ( .D(n4802), .CP(wclk), .Q(ram[561]) );
  DFF ram_reg_1977__0_ ( .D(n4801), .CP(wclk), .Q(ram[560]) );
  DFF ram_reg_1981__7_ ( .D(n4776), .CP(wclk), .Q(ram[535]) );
  DFF ram_reg_1981__6_ ( .D(n4775), .CP(wclk), .Q(ram[534]) );
  DFF ram_reg_1981__5_ ( .D(n4774), .CP(wclk), .Q(ram[533]) );
  DFF ram_reg_1981__4_ ( .D(n4773), .CP(wclk), .Q(ram[532]) );
  DFF ram_reg_1981__3_ ( .D(n4772), .CP(wclk), .Q(ram[531]) );
  DFF ram_reg_1981__2_ ( .D(n4771), .CP(wclk), .Q(ram[530]) );
  DFF ram_reg_1981__1_ ( .D(n4770), .CP(wclk), .Q(ram[529]) );
  DFF ram_reg_1981__0_ ( .D(n4769), .CP(wclk), .Q(ram[528]) );
  DFF ram_reg_1985__7_ ( .D(n4744), .CP(wclk), .Q(ram[503]) );
  DFF ram_reg_1985__6_ ( .D(n4743), .CP(wclk), .Q(ram[502]) );
  DFF ram_reg_1985__5_ ( .D(n4742), .CP(wclk), .Q(ram[501]) );
  DFF ram_reg_1985__4_ ( .D(n4741), .CP(wclk), .Q(ram[500]) );
  DFF ram_reg_1985__3_ ( .D(n4740), .CP(wclk), .Q(ram[499]) );
  DFF ram_reg_1985__2_ ( .D(n4739), .CP(wclk), .Q(ram[498]) );
  DFF ram_reg_1985__1_ ( .D(n4738), .CP(wclk), .Q(ram[497]) );
  DFF ram_reg_1985__0_ ( .D(n4737), .CP(wclk), .Q(ram[496]) );
  DFF ram_reg_1993__7_ ( .D(n4680), .CP(wclk), .Q(ram[439]) );
  DFF ram_reg_1993__6_ ( .D(n4679), .CP(wclk), .Q(ram[438]) );
  DFF ram_reg_1993__5_ ( .D(n4678), .CP(wclk), .Q(ram[437]) );
  DFF ram_reg_1993__4_ ( .D(n4677), .CP(wclk), .Q(ram[436]) );
  DFF ram_reg_1993__3_ ( .D(n4676), .CP(wclk), .Q(ram[435]) );
  DFF ram_reg_1993__2_ ( .D(n4675), .CP(wclk), .Q(ram[434]) );
  DFF ram_reg_1993__1_ ( .D(n4674), .CP(wclk), .Q(ram[433]) );
  DFF ram_reg_1993__0_ ( .D(n4673), .CP(wclk), .Q(ram[432]) );
  DFF ram_reg_1997__7_ ( .D(n4648), .CP(wclk), .Q(ram[407]) );
  DFF ram_reg_1997__6_ ( .D(n4647), .CP(wclk), .Q(ram[406]) );
  DFF ram_reg_1997__5_ ( .D(n4646), .CP(wclk), .Q(ram[405]) );
  DFF ram_reg_1997__4_ ( .D(n4645), .CP(wclk), .Q(ram[404]) );
  DFF ram_reg_1997__3_ ( .D(n4644), .CP(wclk), .Q(ram[403]) );
  DFF ram_reg_1997__2_ ( .D(n4643), .CP(wclk), .Q(ram[402]) );
  DFF ram_reg_1997__1_ ( .D(n4642), .CP(wclk), .Q(ram[401]) );
  DFF ram_reg_1997__0_ ( .D(n4641), .CP(wclk), .Q(ram[400]) );
  DFF ram_reg_2009__7_ ( .D(n4552), .CP(wclk), .Q(ram[311]) );
  DFF ram_reg_2009__6_ ( .D(n4551), .CP(wclk), .Q(ram[310]) );
  DFF ram_reg_2009__5_ ( .D(n4550), .CP(wclk), .Q(ram[309]) );
  DFF ram_reg_2009__4_ ( .D(n4549), .CP(wclk), .Q(ram[308]) );
  DFF ram_reg_2009__3_ ( .D(n4548), .CP(wclk), .Q(ram[307]) );
  DFF ram_reg_2009__2_ ( .D(n4547), .CP(wclk), .Q(ram[306]) );
  DFF ram_reg_2009__1_ ( .D(n4546), .CP(wclk), .Q(ram[305]) );
  DFF ram_reg_2009__0_ ( .D(n4545), .CP(wclk), .Q(ram[304]) );
  DFF ram_reg_2013__7_ ( .D(n4520), .CP(wclk), .Q(ram[279]) );
  DFF ram_reg_2013__6_ ( .D(n4519), .CP(wclk), .Q(ram[278]) );
  DFF ram_reg_2013__5_ ( .D(n4518), .CP(wclk), .Q(ram[277]) );
  DFF ram_reg_2013__4_ ( .D(n4517), .CP(wclk), .Q(ram[276]) );
  DFF ram_reg_2013__3_ ( .D(n4516), .CP(wclk), .Q(ram[275]) );
  DFF ram_reg_2013__2_ ( .D(n4515), .CP(wclk), .Q(ram[274]) );
  DFF ram_reg_2013__1_ ( .D(n4514), .CP(wclk), .Q(ram[273]) );
  DFF ram_reg_2013__0_ ( .D(n4513), .CP(wclk), .Q(ram[272]) );
  DFF ram_reg_2017__7_ ( .D(n4488), .CP(wclk), .Q(ram[247]) );
  DFF ram_reg_2017__6_ ( .D(n4487), .CP(wclk), .Q(ram[246]) );
  DFF ram_reg_2017__5_ ( .D(n4486), .CP(wclk), .Q(ram[245]) );
  DFF ram_reg_2017__4_ ( .D(n4485), .CP(wclk), .Q(ram[244]) );
  DFF ram_reg_2017__3_ ( .D(n4484), .CP(wclk), .Q(ram[243]) );
  DFF ram_reg_2017__2_ ( .D(n4483), .CP(wclk), .Q(ram[242]) );
  DFF ram_reg_2017__1_ ( .D(n4482), .CP(wclk), .Q(ram[241]) );
  DFF ram_reg_2017__0_ ( .D(n4481), .CP(wclk), .Q(ram[240]) );
  DFF ram_reg_2025__7_ ( .D(n4424), .CP(wclk), .Q(ram[183]) );
  DFF ram_reg_2025__6_ ( .D(n4423), .CP(wclk), .Q(ram[182]) );
  DFF ram_reg_2025__5_ ( .D(n4422), .CP(wclk), .Q(ram[181]) );
  DFF ram_reg_2025__4_ ( .D(n4421), .CP(wclk), .Q(ram[180]) );
  DFF ram_reg_2025__3_ ( .D(n4420), .CP(wclk), .Q(ram[179]) );
  DFF ram_reg_2025__2_ ( .D(n4419), .CP(wclk), .Q(ram[178]) );
  DFF ram_reg_2025__1_ ( .D(n4418), .CP(wclk), .Q(ram[177]) );
  DFF ram_reg_2025__0_ ( .D(n4417), .CP(wclk), .Q(ram[176]) );
  DFF ram_reg_2029__7_ ( .D(n4392), .CP(wclk), .Q(ram[151]) );
  DFF ram_reg_2029__6_ ( .D(n4391), .CP(wclk), .Q(ram[150]) );
  DFF ram_reg_2029__5_ ( .D(n4390), .CP(wclk), .Q(ram[149]) );
  DFF ram_reg_2029__4_ ( .D(n4389), .CP(wclk), .Q(ram[148]) );
  DFF ram_reg_2029__3_ ( .D(n4388), .CP(wclk), .Q(ram[147]) );
  DFF ram_reg_2029__2_ ( .D(n4387), .CP(wclk), .Q(ram[146]) );
  DFF ram_reg_2029__1_ ( .D(n4386), .CP(wclk), .Q(ram[145]) );
  DFF ram_reg_2029__0_ ( .D(n4385), .CP(wclk), .Q(ram[144]) );
  DFF ram_reg_2033__7_ ( .D(n4360), .CP(wclk), .Q(ram[119]) );
  DFF ram_reg_2033__6_ ( .D(n4359), .CP(wclk), .Q(ram[118]) );
  DFF ram_reg_2033__5_ ( .D(n4358), .CP(wclk), .Q(ram[117]) );
  DFF ram_reg_2033__4_ ( .D(n4357), .CP(wclk), .Q(ram[116]) );
  DFF ram_reg_2033__3_ ( .D(n4356), .CP(wclk), .Q(ram[115]) );
  DFF ram_reg_2033__2_ ( .D(n4355), .CP(wclk), .Q(ram[114]) );
  DFF ram_reg_2033__1_ ( .D(n4354), .CP(wclk), .Q(ram[113]) );
  DFF ram_reg_2033__0_ ( .D(n4353), .CP(wclk), .Q(ram[112]) );
  DFF ram_reg_2037__7_ ( .D(n4328), .CP(wclk), .Q(ram[87]) );
  DFF ram_reg_2037__6_ ( .D(n4327), .CP(wclk), .Q(ram[86]) );
  DFF ram_reg_2037__5_ ( .D(n4326), .CP(wclk), .Q(ram[85]) );
  DFF ram_reg_2037__4_ ( .D(n4325), .CP(wclk), .Q(ram[84]) );
  DFF ram_reg_2037__3_ ( .D(n4324), .CP(wclk), .Q(ram[83]) );
  DFF ram_reg_2037__2_ ( .D(n4323), .CP(wclk), .Q(ram[82]) );
  DFF ram_reg_2037__1_ ( .D(n4322), .CP(wclk), .Q(ram[81]) );
  DFF ram_reg_2037__0_ ( .D(n4321), .CP(wclk), .Q(ram[80]) );
  DFF ram_reg_2041__7_ ( .D(n4296), .CP(wclk), .Q(ram[55]) );
  DFF ram_reg_2041__6_ ( .D(n4295), .CP(wclk), .Q(ram[54]) );
  DFF ram_reg_2041__5_ ( .D(n4294), .CP(wclk), .Q(ram[53]) );
  DFF ram_reg_2041__4_ ( .D(n4293), .CP(wclk), .Q(ram[52]) );
  DFF ram_reg_2041__3_ ( .D(n4292), .CP(wclk), .Q(ram[51]) );
  DFF ram_reg_2041__2_ ( .D(n4291), .CP(wclk), .Q(ram[50]) );
  DFF ram_reg_2041__1_ ( .D(n4290), .CP(wclk), .Q(ram[49]) );
  DFF ram_reg_2041__0_ ( .D(n4289), .CP(wclk), .Q(ram[48]) );
  DFF ram_reg_2045__7_ ( .D(n4264), .CP(wclk), .Q(ram[23]) );
  DFF ram_reg_2045__6_ ( .D(n4263), .CP(wclk), .Q(ram[22]) );
  DFF ram_reg_2045__5_ ( .D(n4262), .CP(wclk), .Q(ram[21]) );
  DFF ram_reg_2045__4_ ( .D(n4261), .CP(wclk), .Q(ram[20]) );
  DFF ram_reg_2045__3_ ( .D(n4260), .CP(wclk), .Q(ram[19]) );
  DFF ram_reg_2045__2_ ( .D(n4259), .CP(wclk), .Q(ram[18]) );
  DFF ram_reg_2045__1_ ( .D(n4258), .CP(wclk), .Q(ram[17]) );
  DFF ram_reg_2045__0_ ( .D(n4257), .CP(wclk), .Q(ram[16]) );
  DFF ram_reg_11__7_ ( .D(n20536), .CP(wclk), .Q(ram[16295]) );
  DFF ram_reg_11__6_ ( .D(n20535), .CP(wclk), .Q(ram[16294]) );
  DFF ram_reg_11__5_ ( .D(n20534), .CP(wclk), .Q(ram[16293]) );
  DFF ram_reg_11__4_ ( .D(n20533), .CP(wclk), .Q(ram[16292]) );
  DFF ram_reg_11__3_ ( .D(n20532), .CP(wclk), .Q(ram[16291]) );
  DFF ram_reg_11__2_ ( .D(n20531), .CP(wclk), .Q(ram[16290]) );
  DFF ram_reg_11__1_ ( .D(n20530), .CP(wclk), .Q(ram[16289]) );
  DFF ram_reg_11__0_ ( .D(n20529), .CP(wclk), .Q(ram[16288]) );
  DFF ram_reg_43__7_ ( .D(n20280), .CP(wclk), .Q(ram[16039]) );
  DFF ram_reg_43__6_ ( .D(n20279), .CP(wclk), .Q(ram[16038]) );
  DFF ram_reg_43__5_ ( .D(n20278), .CP(wclk), .Q(ram[16037]) );
  DFF ram_reg_43__4_ ( .D(n20277), .CP(wclk), .Q(ram[16036]) );
  DFF ram_reg_43__3_ ( .D(n20276), .CP(wclk), .Q(ram[16035]) );
  DFF ram_reg_43__2_ ( .D(n20275), .CP(wclk), .Q(ram[16034]) );
  DFF ram_reg_43__1_ ( .D(n20274), .CP(wclk), .Q(ram[16033]) );
  DFF ram_reg_43__0_ ( .D(n20273), .CP(wclk), .Q(ram[16032]) );
  DFF ram_reg_47__7_ ( .D(n20248), .CP(wclk), .Q(ram[16007]) );
  DFF ram_reg_47__6_ ( .D(n20247), .CP(wclk), .Q(ram[16006]) );
  DFF ram_reg_47__5_ ( .D(n20246), .CP(wclk), .Q(ram[16005]) );
  DFF ram_reg_47__4_ ( .D(n20245), .CP(wclk), .Q(ram[16004]) );
  DFF ram_reg_47__3_ ( .D(n20244), .CP(wclk), .Q(ram[16003]) );
  DFF ram_reg_47__2_ ( .D(n20243), .CP(wclk), .Q(ram[16002]) );
  DFF ram_reg_47__1_ ( .D(n20242), .CP(wclk), .Q(ram[16001]) );
  DFF ram_reg_47__0_ ( .D(n20241), .CP(wclk), .Q(ram[16000]) );
  DFF ram_reg_59__7_ ( .D(n20152), .CP(wclk), .Q(ram[15911]) );
  DFF ram_reg_59__6_ ( .D(n20151), .CP(wclk), .Q(ram[15910]) );
  DFF ram_reg_59__5_ ( .D(n20150), .CP(wclk), .Q(ram[15909]) );
  DFF ram_reg_59__4_ ( .D(n20149), .CP(wclk), .Q(ram[15908]) );
  DFF ram_reg_59__3_ ( .D(n20148), .CP(wclk), .Q(ram[15907]) );
  DFF ram_reg_59__2_ ( .D(n20147), .CP(wclk), .Q(ram[15906]) );
  DFF ram_reg_59__1_ ( .D(n20146), .CP(wclk), .Q(ram[15905]) );
  DFF ram_reg_59__0_ ( .D(n20145), .CP(wclk), .Q(ram[15904]) );
  DFF ram_reg_63__7_ ( .D(n20120), .CP(wclk), .Q(ram[15879]) );
  DFF ram_reg_63__6_ ( .D(n20119), .CP(wclk), .Q(ram[15878]) );
  DFF ram_reg_63__5_ ( .D(n20118), .CP(wclk), .Q(ram[15877]) );
  DFF ram_reg_63__4_ ( .D(n20117), .CP(wclk), .Q(ram[15876]) );
  DFF ram_reg_63__3_ ( .D(n20116), .CP(wclk), .Q(ram[15875]) );
  DFF ram_reg_63__2_ ( .D(n20115), .CP(wclk), .Q(ram[15874]) );
  DFF ram_reg_63__1_ ( .D(n20114), .CP(wclk), .Q(ram[15873]) );
  DFF ram_reg_63__0_ ( .D(n20113), .CP(wclk), .Q(ram[15872]) );
  DFF ram_reg_123__7_ ( .D(n19640), .CP(wclk), .Q(ram[15399]) );
  DFF ram_reg_123__6_ ( .D(n19639), .CP(wclk), .Q(ram[15398]) );
  DFF ram_reg_123__5_ ( .D(n19638), .CP(wclk), .Q(ram[15397]) );
  DFF ram_reg_123__4_ ( .D(n19637), .CP(wclk), .Q(ram[15396]) );
  DFF ram_reg_123__3_ ( .D(n19636), .CP(wclk), .Q(ram[15395]) );
  DFF ram_reg_123__2_ ( .D(n19635), .CP(wclk), .Q(ram[15394]) );
  DFF ram_reg_123__1_ ( .D(n19634), .CP(wclk), .Q(ram[15393]) );
  DFF ram_reg_123__0_ ( .D(n19633), .CP(wclk), .Q(ram[15392]) );
  DFF ram_reg_131__7_ ( .D(n19576), .CP(wclk), .Q(ram[15335]) );
  DFF ram_reg_131__6_ ( .D(n19575), .CP(wclk), .Q(ram[15334]) );
  DFF ram_reg_131__5_ ( .D(n19574), .CP(wclk), .Q(ram[15333]) );
  DFF ram_reg_131__4_ ( .D(n19573), .CP(wclk), .Q(ram[15332]) );
  DFF ram_reg_131__3_ ( .D(n19572), .CP(wclk), .Q(ram[15331]) );
  DFF ram_reg_131__2_ ( .D(n19571), .CP(wclk), .Q(ram[15330]) );
  DFF ram_reg_131__1_ ( .D(n19570), .CP(wclk), .Q(ram[15329]) );
  DFF ram_reg_131__0_ ( .D(n19569), .CP(wclk), .Q(ram[15328]) );
  DFF ram_reg_139__7_ ( .D(n19512), .CP(wclk), .Q(ram[15271]) );
  DFF ram_reg_139__6_ ( .D(n19511), .CP(wclk), .Q(ram[15270]) );
  DFF ram_reg_139__5_ ( .D(n19510), .CP(wclk), .Q(ram[15269]) );
  DFF ram_reg_139__4_ ( .D(n19509), .CP(wclk), .Q(ram[15268]) );
  DFF ram_reg_139__3_ ( .D(n19508), .CP(wclk), .Q(ram[15267]) );
  DFF ram_reg_139__2_ ( .D(n19507), .CP(wclk), .Q(ram[15266]) );
  DFF ram_reg_139__1_ ( .D(n19506), .CP(wclk), .Q(ram[15265]) );
  DFF ram_reg_139__0_ ( .D(n19505), .CP(wclk), .Q(ram[15264]) );
  DFF ram_reg_143__7_ ( .D(n19480), .CP(wclk), .Q(ram[15239]) );
  DFF ram_reg_143__6_ ( .D(n19479), .CP(wclk), .Q(ram[15238]) );
  DFF ram_reg_143__5_ ( .D(n19478), .CP(wclk), .Q(ram[15237]) );
  DFF ram_reg_143__4_ ( .D(n19477), .CP(wclk), .Q(ram[15236]) );
  DFF ram_reg_143__3_ ( .D(n19476), .CP(wclk), .Q(ram[15235]) );
  DFF ram_reg_143__2_ ( .D(n19475), .CP(wclk), .Q(ram[15234]) );
  DFF ram_reg_143__1_ ( .D(n19474), .CP(wclk), .Q(ram[15233]) );
  DFF ram_reg_143__0_ ( .D(n19473), .CP(wclk), .Q(ram[15232]) );
  DFF ram_reg_155__7_ ( .D(n19384), .CP(wclk), .Q(ram[15143]) );
  DFF ram_reg_155__6_ ( .D(n19383), .CP(wclk), .Q(ram[15142]) );
  DFF ram_reg_155__5_ ( .D(n19382), .CP(wclk), .Q(ram[15141]) );
  DFF ram_reg_155__4_ ( .D(n19381), .CP(wclk), .Q(ram[15140]) );
  DFF ram_reg_155__3_ ( .D(n19380), .CP(wclk), .Q(ram[15139]) );
  DFF ram_reg_155__2_ ( .D(n19379), .CP(wclk), .Q(ram[15138]) );
  DFF ram_reg_155__1_ ( .D(n19378), .CP(wclk), .Q(ram[15137]) );
  DFF ram_reg_155__0_ ( .D(n19377), .CP(wclk), .Q(ram[15136]) );
  DFF ram_reg_159__7_ ( .D(n19352), .CP(wclk), .Q(ram[15111]) );
  DFF ram_reg_159__6_ ( .D(n19351), .CP(wclk), .Q(ram[15110]) );
  DFF ram_reg_159__5_ ( .D(n19350), .CP(wclk), .Q(ram[15109]) );
  DFF ram_reg_159__4_ ( .D(n19349), .CP(wclk), .Q(ram[15108]) );
  DFF ram_reg_159__3_ ( .D(n19348), .CP(wclk), .Q(ram[15107]) );
  DFF ram_reg_159__2_ ( .D(n19347), .CP(wclk), .Q(ram[15106]) );
  DFF ram_reg_159__1_ ( .D(n19346), .CP(wclk), .Q(ram[15105]) );
  DFF ram_reg_159__0_ ( .D(n19345), .CP(wclk), .Q(ram[15104]) );
  DFF ram_reg_163__7_ ( .D(n19320), .CP(wclk), .Q(ram[15079]) );
  DFF ram_reg_163__6_ ( .D(n19319), .CP(wclk), .Q(ram[15078]) );
  DFF ram_reg_163__5_ ( .D(n19318), .CP(wclk), .Q(ram[15077]) );
  DFF ram_reg_163__4_ ( .D(n19317), .CP(wclk), .Q(ram[15076]) );
  DFF ram_reg_163__3_ ( .D(n19316), .CP(wclk), .Q(ram[15075]) );
  DFF ram_reg_163__2_ ( .D(n19315), .CP(wclk), .Q(ram[15074]) );
  DFF ram_reg_163__1_ ( .D(n19314), .CP(wclk), .Q(ram[15073]) );
  DFF ram_reg_163__0_ ( .D(n19313), .CP(wclk), .Q(ram[15072]) );
  DFF ram_reg_171__7_ ( .D(n19256), .CP(wclk), .Q(ram[15015]) );
  DFF ram_reg_171__6_ ( .D(n19255), .CP(wclk), .Q(ram[15014]) );
  DFF ram_reg_171__5_ ( .D(n19254), .CP(wclk), .Q(ram[15013]) );
  DFF ram_reg_171__4_ ( .D(n19253), .CP(wclk), .Q(ram[15012]) );
  DFF ram_reg_171__3_ ( .D(n19252), .CP(wclk), .Q(ram[15011]) );
  DFF ram_reg_171__2_ ( .D(n19251), .CP(wclk), .Q(ram[15010]) );
  DFF ram_reg_171__1_ ( .D(n19250), .CP(wclk), .Q(ram[15009]) );
  DFF ram_reg_171__0_ ( .D(n19249), .CP(wclk), .Q(ram[15008]) );
  DFF ram_reg_175__7_ ( .D(n19224), .CP(wclk), .Q(ram[14983]) );
  DFF ram_reg_175__6_ ( .D(n19223), .CP(wclk), .Q(ram[14982]) );
  DFF ram_reg_175__5_ ( .D(n19222), .CP(wclk), .Q(ram[14981]) );
  DFF ram_reg_175__4_ ( .D(n19221), .CP(wclk), .Q(ram[14980]) );
  DFF ram_reg_175__3_ ( .D(n19220), .CP(wclk), .Q(ram[14979]) );
  DFF ram_reg_175__2_ ( .D(n19219), .CP(wclk), .Q(ram[14978]) );
  DFF ram_reg_175__1_ ( .D(n19218), .CP(wclk), .Q(ram[14977]) );
  DFF ram_reg_175__0_ ( .D(n19217), .CP(wclk), .Q(ram[14976]) );
  DFF ram_reg_179__7_ ( .D(n19192), .CP(wclk), .Q(ram[14951]) );
  DFF ram_reg_179__6_ ( .D(n19191), .CP(wclk), .Q(ram[14950]) );
  DFF ram_reg_179__5_ ( .D(n19190), .CP(wclk), .Q(ram[14949]) );
  DFF ram_reg_179__4_ ( .D(n19189), .CP(wclk), .Q(ram[14948]) );
  DFF ram_reg_179__3_ ( .D(n19188), .CP(wclk), .Q(ram[14947]) );
  DFF ram_reg_179__2_ ( .D(n19187), .CP(wclk), .Q(ram[14946]) );
  DFF ram_reg_179__1_ ( .D(n19186), .CP(wclk), .Q(ram[14945]) );
  DFF ram_reg_179__0_ ( .D(n19185), .CP(wclk), .Q(ram[14944]) );
  DFF ram_reg_183__7_ ( .D(n19160), .CP(wclk), .Q(ram[14919]) );
  DFF ram_reg_183__6_ ( .D(n19159), .CP(wclk), .Q(ram[14918]) );
  DFF ram_reg_183__5_ ( .D(n19158), .CP(wclk), .Q(ram[14917]) );
  DFF ram_reg_183__4_ ( .D(n19157), .CP(wclk), .Q(ram[14916]) );
  DFF ram_reg_183__3_ ( .D(n19156), .CP(wclk), .Q(ram[14915]) );
  DFF ram_reg_183__2_ ( .D(n19155), .CP(wclk), .Q(ram[14914]) );
  DFF ram_reg_183__1_ ( .D(n19154), .CP(wclk), .Q(ram[14913]) );
  DFF ram_reg_183__0_ ( .D(n19153), .CP(wclk), .Q(ram[14912]) );
  DFF ram_reg_187__7_ ( .D(n19128), .CP(wclk), .Q(ram[14887]) );
  DFF ram_reg_187__6_ ( .D(n19127), .CP(wclk), .Q(ram[14886]) );
  DFF ram_reg_187__5_ ( .D(n19126), .CP(wclk), .Q(ram[14885]) );
  DFF ram_reg_187__4_ ( .D(n19125), .CP(wclk), .Q(ram[14884]) );
  DFF ram_reg_187__3_ ( .D(n19124), .CP(wclk), .Q(ram[14883]) );
  DFF ram_reg_187__2_ ( .D(n19123), .CP(wclk), .Q(ram[14882]) );
  DFF ram_reg_187__1_ ( .D(n19122), .CP(wclk), .Q(ram[14881]) );
  DFF ram_reg_187__0_ ( .D(n19121), .CP(wclk), .Q(ram[14880]) );
  DFF ram_reg_191__7_ ( .D(n19096), .CP(wclk), .Q(ram[14855]) );
  DFF ram_reg_191__6_ ( .D(n19095), .CP(wclk), .Q(ram[14854]) );
  DFF ram_reg_191__5_ ( .D(n19094), .CP(wclk), .Q(ram[14853]) );
  DFF ram_reg_191__4_ ( .D(n19093), .CP(wclk), .Q(ram[14852]) );
  DFF ram_reg_191__3_ ( .D(n19092), .CP(wclk), .Q(ram[14851]) );
  DFF ram_reg_191__2_ ( .D(n19091), .CP(wclk), .Q(ram[14850]) );
  DFF ram_reg_191__1_ ( .D(n19090), .CP(wclk), .Q(ram[14849]) );
  DFF ram_reg_191__0_ ( .D(n19089), .CP(wclk), .Q(ram[14848]) );
  DFF ram_reg_203__7_ ( .D(n19000), .CP(wclk), .Q(ram[14759]) );
  DFF ram_reg_203__6_ ( .D(n18999), .CP(wclk), .Q(ram[14758]) );
  DFF ram_reg_203__5_ ( .D(n18998), .CP(wclk), .Q(ram[14757]) );
  DFF ram_reg_203__4_ ( .D(n18997), .CP(wclk), .Q(ram[14756]) );
  DFF ram_reg_203__3_ ( .D(n18996), .CP(wclk), .Q(ram[14755]) );
  DFF ram_reg_203__2_ ( .D(n18995), .CP(wclk), .Q(ram[14754]) );
  DFF ram_reg_203__1_ ( .D(n18994), .CP(wclk), .Q(ram[14753]) );
  DFF ram_reg_203__0_ ( .D(n18993), .CP(wclk), .Q(ram[14752]) );
  DFF ram_reg_207__7_ ( .D(n18968), .CP(wclk), .Q(ram[14727]) );
  DFF ram_reg_207__6_ ( .D(n18967), .CP(wclk), .Q(ram[14726]) );
  DFF ram_reg_207__5_ ( .D(n18966), .CP(wclk), .Q(ram[14725]) );
  DFF ram_reg_207__4_ ( .D(n18965), .CP(wclk), .Q(ram[14724]) );
  DFF ram_reg_207__3_ ( .D(n18964), .CP(wclk), .Q(ram[14723]) );
  DFF ram_reg_207__2_ ( .D(n18963), .CP(wclk), .Q(ram[14722]) );
  DFF ram_reg_207__1_ ( .D(n18962), .CP(wclk), .Q(ram[14721]) );
  DFF ram_reg_207__0_ ( .D(n18961), .CP(wclk), .Q(ram[14720]) );
  DFF ram_reg_219__7_ ( .D(n18872), .CP(wclk), .Q(ram[14631]) );
  DFF ram_reg_219__6_ ( .D(n18871), .CP(wclk), .Q(ram[14630]) );
  DFF ram_reg_219__5_ ( .D(n18870), .CP(wclk), .Q(ram[14629]) );
  DFF ram_reg_219__4_ ( .D(n18869), .CP(wclk), .Q(ram[14628]) );
  DFF ram_reg_219__3_ ( .D(n18868), .CP(wclk), .Q(ram[14627]) );
  DFF ram_reg_219__2_ ( .D(n18867), .CP(wclk), .Q(ram[14626]) );
  DFF ram_reg_219__1_ ( .D(n18866), .CP(wclk), .Q(ram[14625]) );
  DFF ram_reg_219__0_ ( .D(n18865), .CP(wclk), .Q(ram[14624]) );
  DFF ram_reg_223__7_ ( .D(n18840), .CP(wclk), .Q(ram[14599]) );
  DFF ram_reg_223__6_ ( .D(n18839), .CP(wclk), .Q(ram[14598]) );
  DFF ram_reg_223__5_ ( .D(n18838), .CP(wclk), .Q(ram[14597]) );
  DFF ram_reg_223__4_ ( .D(n18837), .CP(wclk), .Q(ram[14596]) );
  DFF ram_reg_223__3_ ( .D(n18836), .CP(wclk), .Q(ram[14595]) );
  DFF ram_reg_223__2_ ( .D(n18835), .CP(wclk), .Q(ram[14594]) );
  DFF ram_reg_223__1_ ( .D(n18834), .CP(wclk), .Q(ram[14593]) );
  DFF ram_reg_223__0_ ( .D(n18833), .CP(wclk), .Q(ram[14592]) );
  DFF ram_reg_227__7_ ( .D(n18808), .CP(wclk), .Q(ram[14567]) );
  DFF ram_reg_227__6_ ( .D(n18807), .CP(wclk), .Q(ram[14566]) );
  DFF ram_reg_227__5_ ( .D(n18806), .CP(wclk), .Q(ram[14565]) );
  DFF ram_reg_227__4_ ( .D(n18805), .CP(wclk), .Q(ram[14564]) );
  DFF ram_reg_227__3_ ( .D(n18804), .CP(wclk), .Q(ram[14563]) );
  DFF ram_reg_227__2_ ( .D(n18803), .CP(wclk), .Q(ram[14562]) );
  DFF ram_reg_227__1_ ( .D(n18802), .CP(wclk), .Q(ram[14561]) );
  DFF ram_reg_227__0_ ( .D(n18801), .CP(wclk), .Q(ram[14560]) );
  DFF ram_reg_235__7_ ( .D(n18744), .CP(wclk), .Q(ram[14503]) );
  DFF ram_reg_235__6_ ( .D(n18743), .CP(wclk), .Q(ram[14502]) );
  DFF ram_reg_235__5_ ( .D(n18742), .CP(wclk), .Q(ram[14501]) );
  DFF ram_reg_235__4_ ( .D(n18741), .CP(wclk), .Q(ram[14500]) );
  DFF ram_reg_235__3_ ( .D(n18740), .CP(wclk), .Q(ram[14499]) );
  DFF ram_reg_235__2_ ( .D(n18739), .CP(wclk), .Q(ram[14498]) );
  DFF ram_reg_235__1_ ( .D(n18738), .CP(wclk), .Q(ram[14497]) );
  DFF ram_reg_235__0_ ( .D(n18737), .CP(wclk), .Q(ram[14496]) );
  DFF ram_reg_239__7_ ( .D(n18712), .CP(wclk), .Q(ram[14471]) );
  DFF ram_reg_239__6_ ( .D(n18711), .CP(wclk), .Q(ram[14470]) );
  DFF ram_reg_239__5_ ( .D(n18710), .CP(wclk), .Q(ram[14469]) );
  DFF ram_reg_239__4_ ( .D(n18709), .CP(wclk), .Q(ram[14468]) );
  DFF ram_reg_239__3_ ( .D(n18708), .CP(wclk), .Q(ram[14467]) );
  DFF ram_reg_239__2_ ( .D(n18707), .CP(wclk), .Q(ram[14466]) );
  DFF ram_reg_239__1_ ( .D(n18706), .CP(wclk), .Q(ram[14465]) );
  DFF ram_reg_239__0_ ( .D(n18705), .CP(wclk), .Q(ram[14464]) );
  DFF ram_reg_243__7_ ( .D(n18680), .CP(wclk), .Q(ram[14439]) );
  DFF ram_reg_243__6_ ( .D(n18679), .CP(wclk), .Q(ram[14438]) );
  DFF ram_reg_243__5_ ( .D(n18678), .CP(wclk), .Q(ram[14437]) );
  DFF ram_reg_243__4_ ( .D(n18677), .CP(wclk), .Q(ram[14436]) );
  DFF ram_reg_243__3_ ( .D(n18676), .CP(wclk), .Q(ram[14435]) );
  DFF ram_reg_243__2_ ( .D(n18675), .CP(wclk), .Q(ram[14434]) );
  DFF ram_reg_243__1_ ( .D(n18674), .CP(wclk), .Q(ram[14433]) );
  DFF ram_reg_243__0_ ( .D(n18673), .CP(wclk), .Q(ram[14432]) );
  DFF ram_reg_251__7_ ( .D(n18616), .CP(wclk), .Q(ram[14375]) );
  DFF ram_reg_251__6_ ( .D(n18615), .CP(wclk), .Q(ram[14374]) );
  DFF ram_reg_251__5_ ( .D(n18614), .CP(wclk), .Q(ram[14373]) );
  DFF ram_reg_251__4_ ( .D(n18613), .CP(wclk), .Q(ram[14372]) );
  DFF ram_reg_251__3_ ( .D(n18612), .CP(wclk), .Q(ram[14371]) );
  DFF ram_reg_251__2_ ( .D(n18611), .CP(wclk), .Q(ram[14370]) );
  DFF ram_reg_251__1_ ( .D(n18610), .CP(wclk), .Q(ram[14369]) );
  DFF ram_reg_251__0_ ( .D(n18609), .CP(wclk), .Q(ram[14368]) );
  DFF ram_reg_255__7_ ( .D(n18584), .CP(wclk), .Q(ram[14343]) );
  DFF ram_reg_255__6_ ( .D(n18583), .CP(wclk), .Q(ram[14342]) );
  DFF ram_reg_255__5_ ( .D(n18582), .CP(wclk), .Q(ram[14341]) );
  DFF ram_reg_255__4_ ( .D(n18581), .CP(wclk), .Q(ram[14340]) );
  DFF ram_reg_255__3_ ( .D(n18580), .CP(wclk), .Q(ram[14339]) );
  DFF ram_reg_255__2_ ( .D(n18579), .CP(wclk), .Q(ram[14338]) );
  DFF ram_reg_255__1_ ( .D(n18578), .CP(wclk), .Q(ram[14337]) );
  DFF ram_reg_255__0_ ( .D(n18577), .CP(wclk), .Q(ram[14336]) );
  DFF ram_reg_267__7_ ( .D(n18488), .CP(wclk), .Q(ram[14247]) );
  DFF ram_reg_267__6_ ( .D(n18487), .CP(wclk), .Q(ram[14246]) );
  DFF ram_reg_267__5_ ( .D(n18486), .CP(wclk), .Q(ram[14245]) );
  DFF ram_reg_267__4_ ( .D(n18485), .CP(wclk), .Q(ram[14244]) );
  DFF ram_reg_267__3_ ( .D(n18484), .CP(wclk), .Q(ram[14243]) );
  DFF ram_reg_267__2_ ( .D(n18483), .CP(wclk), .Q(ram[14242]) );
  DFF ram_reg_267__1_ ( .D(n18482), .CP(wclk), .Q(ram[14241]) );
  DFF ram_reg_267__0_ ( .D(n18481), .CP(wclk), .Q(ram[14240]) );
  DFF ram_reg_271__7_ ( .D(n18456), .CP(wclk), .Q(ram[14215]) );
  DFF ram_reg_271__6_ ( .D(n18455), .CP(wclk), .Q(ram[14214]) );
  DFF ram_reg_271__5_ ( .D(n18454), .CP(wclk), .Q(ram[14213]) );
  DFF ram_reg_271__4_ ( .D(n18453), .CP(wclk), .Q(ram[14212]) );
  DFF ram_reg_271__3_ ( .D(n18452), .CP(wclk), .Q(ram[14211]) );
  DFF ram_reg_271__2_ ( .D(n18451), .CP(wclk), .Q(ram[14210]) );
  DFF ram_reg_271__1_ ( .D(n18450), .CP(wclk), .Q(ram[14209]) );
  DFF ram_reg_271__0_ ( .D(n18449), .CP(wclk), .Q(ram[14208]) );
  DFF ram_reg_283__7_ ( .D(n18360), .CP(wclk), .Q(ram[14119]) );
  DFF ram_reg_283__6_ ( .D(n18359), .CP(wclk), .Q(ram[14118]) );
  DFF ram_reg_283__5_ ( .D(n18358), .CP(wclk), .Q(ram[14117]) );
  DFF ram_reg_283__4_ ( .D(n18357), .CP(wclk), .Q(ram[14116]) );
  DFF ram_reg_283__3_ ( .D(n18356), .CP(wclk), .Q(ram[14115]) );
  DFF ram_reg_283__2_ ( .D(n18355), .CP(wclk), .Q(ram[14114]) );
  DFF ram_reg_283__1_ ( .D(n18354), .CP(wclk), .Q(ram[14113]) );
  DFF ram_reg_283__0_ ( .D(n18353), .CP(wclk), .Q(ram[14112]) );
  DFF ram_reg_299__7_ ( .D(n18232), .CP(wclk), .Q(ram[13991]) );
  DFF ram_reg_299__6_ ( .D(n18231), .CP(wclk), .Q(ram[13990]) );
  DFF ram_reg_299__5_ ( .D(n18230), .CP(wclk), .Q(ram[13989]) );
  DFF ram_reg_299__4_ ( .D(n18229), .CP(wclk), .Q(ram[13988]) );
  DFF ram_reg_299__3_ ( .D(n18228), .CP(wclk), .Q(ram[13987]) );
  DFF ram_reg_299__2_ ( .D(n18227), .CP(wclk), .Q(ram[13986]) );
  DFF ram_reg_299__1_ ( .D(n18226), .CP(wclk), .Q(ram[13985]) );
  DFF ram_reg_299__0_ ( .D(n18225), .CP(wclk), .Q(ram[13984]) );
  DFF ram_reg_303__7_ ( .D(n18200), .CP(wclk), .Q(ram[13959]) );
  DFF ram_reg_303__6_ ( .D(n18199), .CP(wclk), .Q(ram[13958]) );
  DFF ram_reg_303__5_ ( .D(n18198), .CP(wclk), .Q(ram[13957]) );
  DFF ram_reg_303__4_ ( .D(n18197), .CP(wclk), .Q(ram[13956]) );
  DFF ram_reg_303__3_ ( .D(n18196), .CP(wclk), .Q(ram[13955]) );
  DFF ram_reg_303__2_ ( .D(n18195), .CP(wclk), .Q(ram[13954]) );
  DFF ram_reg_303__1_ ( .D(n18194), .CP(wclk), .Q(ram[13953]) );
  DFF ram_reg_303__0_ ( .D(n18193), .CP(wclk), .Q(ram[13952]) );
  DFF ram_reg_315__7_ ( .D(n18104), .CP(wclk), .Q(ram[13863]) );
  DFF ram_reg_315__6_ ( .D(n18103), .CP(wclk), .Q(ram[13862]) );
  DFF ram_reg_315__5_ ( .D(n18102), .CP(wclk), .Q(ram[13861]) );
  DFF ram_reg_315__4_ ( .D(n18101), .CP(wclk), .Q(ram[13860]) );
  DFF ram_reg_315__3_ ( .D(n18100), .CP(wclk), .Q(ram[13859]) );
  DFF ram_reg_315__2_ ( .D(n18099), .CP(wclk), .Q(ram[13858]) );
  DFF ram_reg_315__1_ ( .D(n18098), .CP(wclk), .Q(ram[13857]) );
  DFF ram_reg_315__0_ ( .D(n18097), .CP(wclk), .Q(ram[13856]) );
  DFF ram_reg_319__7_ ( .D(n18072), .CP(wclk), .Q(ram[13831]) );
  DFF ram_reg_319__6_ ( .D(n18071), .CP(wclk), .Q(ram[13830]) );
  DFF ram_reg_319__5_ ( .D(n18070), .CP(wclk), .Q(ram[13829]) );
  DFF ram_reg_319__4_ ( .D(n18069), .CP(wclk), .Q(ram[13828]) );
  DFF ram_reg_319__3_ ( .D(n18068), .CP(wclk), .Q(ram[13827]) );
  DFF ram_reg_319__2_ ( .D(n18067), .CP(wclk), .Q(ram[13826]) );
  DFF ram_reg_319__1_ ( .D(n18066), .CP(wclk), .Q(ram[13825]) );
  DFF ram_reg_319__0_ ( .D(n18065), .CP(wclk), .Q(ram[13824]) );
  DFF ram_reg_363__7_ ( .D(n17720), .CP(wclk), .Q(ram[13479]) );
  DFF ram_reg_363__6_ ( .D(n17719), .CP(wclk), .Q(ram[13478]) );
  DFF ram_reg_363__5_ ( .D(n17718), .CP(wclk), .Q(ram[13477]) );
  DFF ram_reg_363__4_ ( .D(n17717), .CP(wclk), .Q(ram[13476]) );
  DFF ram_reg_363__3_ ( .D(n17716), .CP(wclk), .Q(ram[13475]) );
  DFF ram_reg_363__2_ ( .D(n17715), .CP(wclk), .Q(ram[13474]) );
  DFF ram_reg_363__1_ ( .D(n17714), .CP(wclk), .Q(ram[13473]) );
  DFF ram_reg_363__0_ ( .D(n17713), .CP(wclk), .Q(ram[13472]) );
  DFF ram_reg_379__7_ ( .D(n17592), .CP(wclk), .Q(ram[13351]) );
  DFF ram_reg_379__6_ ( .D(n17591), .CP(wclk), .Q(ram[13350]) );
  DFF ram_reg_379__5_ ( .D(n17590), .CP(wclk), .Q(ram[13349]) );
  DFF ram_reg_379__4_ ( .D(n17589), .CP(wclk), .Q(ram[13348]) );
  DFF ram_reg_379__3_ ( .D(n17588), .CP(wclk), .Q(ram[13347]) );
  DFF ram_reg_379__2_ ( .D(n17587), .CP(wclk), .Q(ram[13346]) );
  DFF ram_reg_379__1_ ( .D(n17586), .CP(wclk), .Q(ram[13345]) );
  DFF ram_reg_379__0_ ( .D(n17585), .CP(wclk), .Q(ram[13344]) );
  DFF ram_reg_387__7_ ( .D(n17528), .CP(wclk), .Q(ram[13287]) );
  DFF ram_reg_387__6_ ( .D(n17527), .CP(wclk), .Q(ram[13286]) );
  DFF ram_reg_387__5_ ( .D(n17526), .CP(wclk), .Q(ram[13285]) );
  DFF ram_reg_387__4_ ( .D(n17525), .CP(wclk), .Q(ram[13284]) );
  DFF ram_reg_387__3_ ( .D(n17524), .CP(wclk), .Q(ram[13283]) );
  DFF ram_reg_387__2_ ( .D(n17523), .CP(wclk), .Q(ram[13282]) );
  DFF ram_reg_387__1_ ( .D(n17522), .CP(wclk), .Q(ram[13281]) );
  DFF ram_reg_387__0_ ( .D(n17521), .CP(wclk), .Q(ram[13280]) );
  DFF ram_reg_395__7_ ( .D(n17464), .CP(wclk), .Q(ram[13223]) );
  DFF ram_reg_395__6_ ( .D(n17463), .CP(wclk), .Q(ram[13222]) );
  DFF ram_reg_395__5_ ( .D(n17462), .CP(wclk), .Q(ram[13221]) );
  DFF ram_reg_395__4_ ( .D(n17461), .CP(wclk), .Q(ram[13220]) );
  DFF ram_reg_395__3_ ( .D(n17460), .CP(wclk), .Q(ram[13219]) );
  DFF ram_reg_395__2_ ( .D(n17459), .CP(wclk), .Q(ram[13218]) );
  DFF ram_reg_395__1_ ( .D(n17458), .CP(wclk), .Q(ram[13217]) );
  DFF ram_reg_395__0_ ( .D(n17457), .CP(wclk), .Q(ram[13216]) );
  DFF ram_reg_399__7_ ( .D(n17432), .CP(wclk), .Q(ram[13191]) );
  DFF ram_reg_399__6_ ( .D(n17431), .CP(wclk), .Q(ram[13190]) );
  DFF ram_reg_399__5_ ( .D(n17430), .CP(wclk), .Q(ram[13189]) );
  DFF ram_reg_399__4_ ( .D(n17429), .CP(wclk), .Q(ram[13188]) );
  DFF ram_reg_399__3_ ( .D(n17428), .CP(wclk), .Q(ram[13187]) );
  DFF ram_reg_399__2_ ( .D(n17427), .CP(wclk), .Q(ram[13186]) );
  DFF ram_reg_399__1_ ( .D(n17426), .CP(wclk), .Q(ram[13185]) );
  DFF ram_reg_399__0_ ( .D(n17425), .CP(wclk), .Q(ram[13184]) );
  DFF ram_reg_403__7_ ( .D(n17400), .CP(wclk), .Q(ram[13159]) );
  DFF ram_reg_403__6_ ( .D(n17399), .CP(wclk), .Q(ram[13158]) );
  DFF ram_reg_403__5_ ( .D(n17398), .CP(wclk), .Q(ram[13157]) );
  DFF ram_reg_403__4_ ( .D(n17397), .CP(wclk), .Q(ram[13156]) );
  DFF ram_reg_403__3_ ( .D(n17396), .CP(wclk), .Q(ram[13155]) );
  DFF ram_reg_403__2_ ( .D(n17395), .CP(wclk), .Q(ram[13154]) );
  DFF ram_reg_403__1_ ( .D(n17394), .CP(wclk), .Q(ram[13153]) );
  DFF ram_reg_403__0_ ( .D(n17393), .CP(wclk), .Q(ram[13152]) );
  DFF ram_reg_411__7_ ( .D(n17336), .CP(wclk), .Q(ram[13095]) );
  DFF ram_reg_411__6_ ( .D(n17335), .CP(wclk), .Q(ram[13094]) );
  DFF ram_reg_411__5_ ( .D(n17334), .CP(wclk), .Q(ram[13093]) );
  DFF ram_reg_411__4_ ( .D(n17333), .CP(wclk), .Q(ram[13092]) );
  DFF ram_reg_411__3_ ( .D(n17332), .CP(wclk), .Q(ram[13091]) );
  DFF ram_reg_411__2_ ( .D(n17331), .CP(wclk), .Q(ram[13090]) );
  DFF ram_reg_411__1_ ( .D(n17330), .CP(wclk), .Q(ram[13089]) );
  DFF ram_reg_411__0_ ( .D(n17329), .CP(wclk), .Q(ram[13088]) );
  DFF ram_reg_415__7_ ( .D(n17304), .CP(wclk), .Q(ram[13063]) );
  DFF ram_reg_415__6_ ( .D(n17303), .CP(wclk), .Q(ram[13062]) );
  DFF ram_reg_415__5_ ( .D(n17302), .CP(wclk), .Q(ram[13061]) );
  DFF ram_reg_415__4_ ( .D(n17301), .CP(wclk), .Q(ram[13060]) );
  DFF ram_reg_415__3_ ( .D(n17300), .CP(wclk), .Q(ram[13059]) );
  DFF ram_reg_415__2_ ( .D(n17299), .CP(wclk), .Q(ram[13058]) );
  DFF ram_reg_415__1_ ( .D(n17298), .CP(wclk), .Q(ram[13057]) );
  DFF ram_reg_415__0_ ( .D(n17297), .CP(wclk), .Q(ram[13056]) );
  DFF ram_reg_419__7_ ( .D(n17272), .CP(wclk), .Q(ram[13031]) );
  DFF ram_reg_419__6_ ( .D(n17271), .CP(wclk), .Q(ram[13030]) );
  DFF ram_reg_419__5_ ( .D(n17270), .CP(wclk), .Q(ram[13029]) );
  DFF ram_reg_419__4_ ( .D(n17269), .CP(wclk), .Q(ram[13028]) );
  DFF ram_reg_419__3_ ( .D(n17268), .CP(wclk), .Q(ram[13027]) );
  DFF ram_reg_419__2_ ( .D(n17267), .CP(wclk), .Q(ram[13026]) );
  DFF ram_reg_419__1_ ( .D(n17266), .CP(wclk), .Q(ram[13025]) );
  DFF ram_reg_419__0_ ( .D(n17265), .CP(wclk), .Q(ram[13024]) );
  DFF ram_reg_423__7_ ( .D(n17240), .CP(wclk), .Q(ram[12999]) );
  DFF ram_reg_423__6_ ( .D(n17239), .CP(wclk), .Q(ram[12998]) );
  DFF ram_reg_423__5_ ( .D(n17238), .CP(wclk), .Q(ram[12997]) );
  DFF ram_reg_423__4_ ( .D(n17237), .CP(wclk), .Q(ram[12996]) );
  DFF ram_reg_423__3_ ( .D(n17236), .CP(wclk), .Q(ram[12995]) );
  DFF ram_reg_423__2_ ( .D(n17235), .CP(wclk), .Q(ram[12994]) );
  DFF ram_reg_423__1_ ( .D(n17234), .CP(wclk), .Q(ram[12993]) );
  DFF ram_reg_423__0_ ( .D(n17233), .CP(wclk), .Q(ram[12992]) );
  DFF ram_reg_427__7_ ( .D(n17208), .CP(wclk), .Q(ram[12967]) );
  DFF ram_reg_427__6_ ( .D(n17207), .CP(wclk), .Q(ram[12966]) );
  DFF ram_reg_427__5_ ( .D(n17206), .CP(wclk), .Q(ram[12965]) );
  DFF ram_reg_427__4_ ( .D(n17205), .CP(wclk), .Q(ram[12964]) );
  DFF ram_reg_427__3_ ( .D(n17204), .CP(wclk), .Q(ram[12963]) );
  DFF ram_reg_427__2_ ( .D(n17203), .CP(wclk), .Q(ram[12962]) );
  DFF ram_reg_427__1_ ( .D(n17202), .CP(wclk), .Q(ram[12961]) );
  DFF ram_reg_427__0_ ( .D(n17201), .CP(wclk), .Q(ram[12960]) );
  DFF ram_reg_431__7_ ( .D(n17176), .CP(wclk), .Q(ram[12935]) );
  DFF ram_reg_431__6_ ( .D(n17175), .CP(wclk), .Q(ram[12934]) );
  DFF ram_reg_431__5_ ( .D(n17174), .CP(wclk), .Q(ram[12933]) );
  DFF ram_reg_431__4_ ( .D(n17173), .CP(wclk), .Q(ram[12932]) );
  DFF ram_reg_431__3_ ( .D(n17172), .CP(wclk), .Q(ram[12931]) );
  DFF ram_reg_431__2_ ( .D(n17171), .CP(wclk), .Q(ram[12930]) );
  DFF ram_reg_431__1_ ( .D(n17170), .CP(wclk), .Q(ram[12929]) );
  DFF ram_reg_431__0_ ( .D(n17169), .CP(wclk), .Q(ram[12928]) );
  DFF ram_reg_435__7_ ( .D(n17144), .CP(wclk), .Q(ram[12903]) );
  DFF ram_reg_435__6_ ( .D(n17143), .CP(wclk), .Q(ram[12902]) );
  DFF ram_reg_435__5_ ( .D(n17142), .CP(wclk), .Q(ram[12901]) );
  DFF ram_reg_435__4_ ( .D(n17141), .CP(wclk), .Q(ram[12900]) );
  DFF ram_reg_435__3_ ( .D(n17140), .CP(wclk), .Q(ram[12899]) );
  DFF ram_reg_435__2_ ( .D(n17139), .CP(wclk), .Q(ram[12898]) );
  DFF ram_reg_435__1_ ( .D(n17138), .CP(wclk), .Q(ram[12897]) );
  DFF ram_reg_435__0_ ( .D(n17137), .CP(wclk), .Q(ram[12896]) );
  DFF ram_reg_439__7_ ( .D(n17112), .CP(wclk), .Q(ram[12871]) );
  DFF ram_reg_439__6_ ( .D(n17111), .CP(wclk), .Q(ram[12870]) );
  DFF ram_reg_439__5_ ( .D(n17110), .CP(wclk), .Q(ram[12869]) );
  DFF ram_reg_439__4_ ( .D(n17109), .CP(wclk), .Q(ram[12868]) );
  DFF ram_reg_439__3_ ( .D(n17108), .CP(wclk), .Q(ram[12867]) );
  DFF ram_reg_439__2_ ( .D(n17107), .CP(wclk), .Q(ram[12866]) );
  DFF ram_reg_439__1_ ( .D(n17106), .CP(wclk), .Q(ram[12865]) );
  DFF ram_reg_439__0_ ( .D(n17105), .CP(wclk), .Q(ram[12864]) );
  DFF ram_reg_443__7_ ( .D(n17080), .CP(wclk), .Q(ram[12839]) );
  DFF ram_reg_443__6_ ( .D(n17079), .CP(wclk), .Q(ram[12838]) );
  DFF ram_reg_443__5_ ( .D(n17078), .CP(wclk), .Q(ram[12837]) );
  DFF ram_reg_443__4_ ( .D(n17077), .CP(wclk), .Q(ram[12836]) );
  DFF ram_reg_443__3_ ( .D(n17076), .CP(wclk), .Q(ram[12835]) );
  DFF ram_reg_443__2_ ( .D(n17075), .CP(wclk), .Q(ram[12834]) );
  DFF ram_reg_443__1_ ( .D(n17074), .CP(wclk), .Q(ram[12833]) );
  DFF ram_reg_443__0_ ( .D(n17073), .CP(wclk), .Q(ram[12832]) );
  DFF ram_reg_447__7_ ( .D(n17048), .CP(wclk), .Q(ram[12807]) );
  DFF ram_reg_447__6_ ( .D(n17047), .CP(wclk), .Q(ram[12806]) );
  DFF ram_reg_447__5_ ( .D(n17046), .CP(wclk), .Q(ram[12805]) );
  DFF ram_reg_447__4_ ( .D(n17045), .CP(wclk), .Q(ram[12804]) );
  DFF ram_reg_447__3_ ( .D(n17044), .CP(wclk), .Q(ram[12803]) );
  DFF ram_reg_447__2_ ( .D(n17043), .CP(wclk), .Q(ram[12802]) );
  DFF ram_reg_447__1_ ( .D(n17042), .CP(wclk), .Q(ram[12801]) );
  DFF ram_reg_447__0_ ( .D(n17041), .CP(wclk), .Q(ram[12800]) );
  DFF ram_reg_451__7_ ( .D(n17016), .CP(wclk), .Q(ram[12775]) );
  DFF ram_reg_451__6_ ( .D(n17015), .CP(wclk), .Q(ram[12774]) );
  DFF ram_reg_451__5_ ( .D(n17014), .CP(wclk), .Q(ram[12773]) );
  DFF ram_reg_451__4_ ( .D(n17013), .CP(wclk), .Q(ram[12772]) );
  DFF ram_reg_451__3_ ( .D(n17012), .CP(wclk), .Q(ram[12771]) );
  DFF ram_reg_451__2_ ( .D(n17011), .CP(wclk), .Q(ram[12770]) );
  DFF ram_reg_451__1_ ( .D(n17010), .CP(wclk), .Q(ram[12769]) );
  DFF ram_reg_451__0_ ( .D(n17009), .CP(wclk), .Q(ram[12768]) );
  DFF ram_reg_459__7_ ( .D(n16952), .CP(wclk), .Q(ram[12711]) );
  DFF ram_reg_459__6_ ( .D(n16951), .CP(wclk), .Q(ram[12710]) );
  DFF ram_reg_459__5_ ( .D(n16950), .CP(wclk), .Q(ram[12709]) );
  DFF ram_reg_459__4_ ( .D(n16949), .CP(wclk), .Q(ram[12708]) );
  DFF ram_reg_459__3_ ( .D(n16948), .CP(wclk), .Q(ram[12707]) );
  DFF ram_reg_459__2_ ( .D(n16947), .CP(wclk), .Q(ram[12706]) );
  DFF ram_reg_459__1_ ( .D(n16946), .CP(wclk), .Q(ram[12705]) );
  DFF ram_reg_459__0_ ( .D(n16945), .CP(wclk), .Q(ram[12704]) );
  DFF ram_reg_463__7_ ( .D(n16920), .CP(wclk), .Q(ram[12679]) );
  DFF ram_reg_463__6_ ( .D(n16919), .CP(wclk), .Q(ram[12678]) );
  DFF ram_reg_463__5_ ( .D(n16918), .CP(wclk), .Q(ram[12677]) );
  DFF ram_reg_463__4_ ( .D(n16917), .CP(wclk), .Q(ram[12676]) );
  DFF ram_reg_463__3_ ( .D(n16916), .CP(wclk), .Q(ram[12675]) );
  DFF ram_reg_463__2_ ( .D(n16915), .CP(wclk), .Q(ram[12674]) );
  DFF ram_reg_463__1_ ( .D(n16914), .CP(wclk), .Q(ram[12673]) );
  DFF ram_reg_463__0_ ( .D(n16913), .CP(wclk), .Q(ram[12672]) );
  DFF ram_reg_475__7_ ( .D(n16824), .CP(wclk), .Q(ram[12583]) );
  DFF ram_reg_475__6_ ( .D(n16823), .CP(wclk), .Q(ram[12582]) );
  DFF ram_reg_475__5_ ( .D(n16822), .CP(wclk), .Q(ram[12581]) );
  DFF ram_reg_475__4_ ( .D(n16821), .CP(wclk), .Q(ram[12580]) );
  DFF ram_reg_475__3_ ( .D(n16820), .CP(wclk), .Q(ram[12579]) );
  DFF ram_reg_475__2_ ( .D(n16819), .CP(wclk), .Q(ram[12578]) );
  DFF ram_reg_475__1_ ( .D(n16818), .CP(wclk), .Q(ram[12577]) );
  DFF ram_reg_475__0_ ( .D(n16817), .CP(wclk), .Q(ram[12576]) );
  DFF ram_reg_479__7_ ( .D(n16792), .CP(wclk), .Q(ram[12551]) );
  DFF ram_reg_479__6_ ( .D(n16791), .CP(wclk), .Q(ram[12550]) );
  DFF ram_reg_479__5_ ( .D(n16790), .CP(wclk), .Q(ram[12549]) );
  DFF ram_reg_479__4_ ( .D(n16789), .CP(wclk), .Q(ram[12548]) );
  DFF ram_reg_479__3_ ( .D(n16788), .CP(wclk), .Q(ram[12547]) );
  DFF ram_reg_479__2_ ( .D(n16787), .CP(wclk), .Q(ram[12546]) );
  DFF ram_reg_479__1_ ( .D(n16786), .CP(wclk), .Q(ram[12545]) );
  DFF ram_reg_479__0_ ( .D(n16785), .CP(wclk), .Q(ram[12544]) );
  DFF ram_reg_483__7_ ( .D(n16760), .CP(wclk), .Q(ram[12519]) );
  DFF ram_reg_483__6_ ( .D(n16759), .CP(wclk), .Q(ram[12518]) );
  DFF ram_reg_483__5_ ( .D(n16758), .CP(wclk), .Q(ram[12517]) );
  DFF ram_reg_483__4_ ( .D(n16757), .CP(wclk), .Q(ram[12516]) );
  DFF ram_reg_483__3_ ( .D(n16756), .CP(wclk), .Q(ram[12515]) );
  DFF ram_reg_483__2_ ( .D(n16755), .CP(wclk), .Q(ram[12514]) );
  DFF ram_reg_483__1_ ( .D(n16754), .CP(wclk), .Q(ram[12513]) );
  DFF ram_reg_483__0_ ( .D(n16753), .CP(wclk), .Q(ram[12512]) );
  DFF ram_reg_491__7_ ( .D(n16696), .CP(wclk), .Q(ram[12455]) );
  DFF ram_reg_491__6_ ( .D(n16695), .CP(wclk), .Q(ram[12454]) );
  DFF ram_reg_491__5_ ( .D(n16694), .CP(wclk), .Q(ram[12453]) );
  DFF ram_reg_491__4_ ( .D(n16693), .CP(wclk), .Q(ram[12452]) );
  DFF ram_reg_491__3_ ( .D(n16692), .CP(wclk), .Q(ram[12451]) );
  DFF ram_reg_491__2_ ( .D(n16691), .CP(wclk), .Q(ram[12450]) );
  DFF ram_reg_491__1_ ( .D(n16690), .CP(wclk), .Q(ram[12449]) );
  DFF ram_reg_491__0_ ( .D(n16689), .CP(wclk), .Q(ram[12448]) );
  DFF ram_reg_495__7_ ( .D(n16664), .CP(wclk), .Q(ram[12423]) );
  DFF ram_reg_495__6_ ( .D(n16663), .CP(wclk), .Q(ram[12422]) );
  DFF ram_reg_495__5_ ( .D(n16662), .CP(wclk), .Q(ram[12421]) );
  DFF ram_reg_495__4_ ( .D(n16661), .CP(wclk), .Q(ram[12420]) );
  DFF ram_reg_495__3_ ( .D(n16660), .CP(wclk), .Q(ram[12419]) );
  DFF ram_reg_495__2_ ( .D(n16659), .CP(wclk), .Q(ram[12418]) );
  DFF ram_reg_495__1_ ( .D(n16658), .CP(wclk), .Q(ram[12417]) );
  DFF ram_reg_495__0_ ( .D(n16657), .CP(wclk), .Q(ram[12416]) );
  DFF ram_reg_499__7_ ( .D(n16632), .CP(wclk), .Q(ram[12391]) );
  DFF ram_reg_499__6_ ( .D(n16631), .CP(wclk), .Q(ram[12390]) );
  DFF ram_reg_499__5_ ( .D(n16630), .CP(wclk), .Q(ram[12389]) );
  DFF ram_reg_499__4_ ( .D(n16629), .CP(wclk), .Q(ram[12388]) );
  DFF ram_reg_499__3_ ( .D(n16628), .CP(wclk), .Q(ram[12387]) );
  DFF ram_reg_499__2_ ( .D(n16627), .CP(wclk), .Q(ram[12386]) );
  DFF ram_reg_499__1_ ( .D(n16626), .CP(wclk), .Q(ram[12385]) );
  DFF ram_reg_499__0_ ( .D(n16625), .CP(wclk), .Q(ram[12384]) );
  DFF ram_reg_507__7_ ( .D(n16568), .CP(wclk), .Q(ram[12327]) );
  DFF ram_reg_507__6_ ( .D(n16567), .CP(wclk), .Q(ram[12326]) );
  DFF ram_reg_507__5_ ( .D(n16566), .CP(wclk), .Q(ram[12325]) );
  DFF ram_reg_507__4_ ( .D(n16565), .CP(wclk), .Q(ram[12324]) );
  DFF ram_reg_507__3_ ( .D(n16564), .CP(wclk), .Q(ram[12323]) );
  DFF ram_reg_507__2_ ( .D(n16563), .CP(wclk), .Q(ram[12322]) );
  DFF ram_reg_507__1_ ( .D(n16562), .CP(wclk), .Q(ram[12321]) );
  DFF ram_reg_507__0_ ( .D(n16561), .CP(wclk), .Q(ram[12320]) );
  DFF ram_reg_511__7_ ( .D(n16536), .CP(wclk), .Q(ram[12295]) );
  DFF ram_reg_511__6_ ( .D(n16535), .CP(wclk), .Q(ram[12294]) );
  DFF ram_reg_511__5_ ( .D(n16534), .CP(wclk), .Q(ram[12293]) );
  DFF ram_reg_511__4_ ( .D(n16533), .CP(wclk), .Q(ram[12292]) );
  DFF ram_reg_511__3_ ( .D(n16532), .CP(wclk), .Q(ram[12291]) );
  DFF ram_reg_511__2_ ( .D(n16531), .CP(wclk), .Q(ram[12290]) );
  DFF ram_reg_511__1_ ( .D(n16530), .CP(wclk), .Q(ram[12289]) );
  DFF ram_reg_511__0_ ( .D(n16529), .CP(wclk), .Q(ram[12288]) );
  DFF ram_reg_523__7_ ( .D(n16440), .CP(wclk), .Q(ram[12199]) );
  DFF ram_reg_523__6_ ( .D(n16439), .CP(wclk), .Q(ram[12198]) );
  DFF ram_reg_523__5_ ( .D(n16438), .CP(wclk), .Q(ram[12197]) );
  DFF ram_reg_523__4_ ( .D(n16437), .CP(wclk), .Q(ram[12196]) );
  DFF ram_reg_523__3_ ( .D(n16436), .CP(wclk), .Q(ram[12195]) );
  DFF ram_reg_523__2_ ( .D(n16435), .CP(wclk), .Q(ram[12194]) );
  DFF ram_reg_523__1_ ( .D(n16434), .CP(wclk), .Q(ram[12193]) );
  DFF ram_reg_523__0_ ( .D(n16433), .CP(wclk), .Q(ram[12192]) );
  DFF ram_reg_527__7_ ( .D(n16408), .CP(wclk), .Q(ram[12167]) );
  DFF ram_reg_527__6_ ( .D(n16407), .CP(wclk), .Q(ram[12166]) );
  DFF ram_reg_527__5_ ( .D(n16406), .CP(wclk), .Q(ram[12165]) );
  DFF ram_reg_527__4_ ( .D(n16405), .CP(wclk), .Q(ram[12164]) );
  DFF ram_reg_527__3_ ( .D(n16404), .CP(wclk), .Q(ram[12163]) );
  DFF ram_reg_527__2_ ( .D(n16403), .CP(wclk), .Q(ram[12162]) );
  DFF ram_reg_527__1_ ( .D(n16402), .CP(wclk), .Q(ram[12161]) );
  DFF ram_reg_527__0_ ( .D(n16401), .CP(wclk), .Q(ram[12160]) );
  DFF ram_reg_539__7_ ( .D(n16312), .CP(wclk), .Q(ram[12071]) );
  DFF ram_reg_539__6_ ( .D(n16311), .CP(wclk), .Q(ram[12070]) );
  DFF ram_reg_539__5_ ( .D(n16310), .CP(wclk), .Q(ram[12069]) );
  DFF ram_reg_539__4_ ( .D(n16309), .CP(wclk), .Q(ram[12068]) );
  DFF ram_reg_539__3_ ( .D(n16308), .CP(wclk), .Q(ram[12067]) );
  DFF ram_reg_539__2_ ( .D(n16307), .CP(wclk), .Q(ram[12066]) );
  DFF ram_reg_539__1_ ( .D(n16306), .CP(wclk), .Q(ram[12065]) );
  DFF ram_reg_539__0_ ( .D(n16305), .CP(wclk), .Q(ram[12064]) );
  DFF ram_reg_543__7_ ( .D(n16280), .CP(wclk), .Q(ram[12039]) );
  DFF ram_reg_543__6_ ( .D(n16279), .CP(wclk), .Q(ram[12038]) );
  DFF ram_reg_543__5_ ( .D(n16278), .CP(wclk), .Q(ram[12037]) );
  DFF ram_reg_543__4_ ( .D(n16277), .CP(wclk), .Q(ram[12036]) );
  DFF ram_reg_543__3_ ( .D(n16276), .CP(wclk), .Q(ram[12035]) );
  DFF ram_reg_543__2_ ( .D(n16275), .CP(wclk), .Q(ram[12034]) );
  DFF ram_reg_543__1_ ( .D(n16274), .CP(wclk), .Q(ram[12033]) );
  DFF ram_reg_543__0_ ( .D(n16273), .CP(wclk), .Q(ram[12032]) );
  DFF ram_reg_547__7_ ( .D(n16248), .CP(wclk), .Q(ram[12007]) );
  DFF ram_reg_547__6_ ( .D(n16247), .CP(wclk), .Q(ram[12006]) );
  DFF ram_reg_547__5_ ( .D(n16246), .CP(wclk), .Q(ram[12005]) );
  DFF ram_reg_547__4_ ( .D(n16245), .CP(wclk), .Q(ram[12004]) );
  DFF ram_reg_547__3_ ( .D(n16244), .CP(wclk), .Q(ram[12003]) );
  DFF ram_reg_547__2_ ( .D(n16243), .CP(wclk), .Q(ram[12002]) );
  DFF ram_reg_547__1_ ( .D(n16242), .CP(wclk), .Q(ram[12001]) );
  DFF ram_reg_547__0_ ( .D(n16241), .CP(wclk), .Q(ram[12000]) );
  DFF ram_reg_555__7_ ( .D(n16184), .CP(wclk), .Q(ram[11943]) );
  DFF ram_reg_555__6_ ( .D(n16183), .CP(wclk), .Q(ram[11942]) );
  DFF ram_reg_555__5_ ( .D(n16182), .CP(wclk), .Q(ram[11941]) );
  DFF ram_reg_555__4_ ( .D(n16181), .CP(wclk), .Q(ram[11940]) );
  DFF ram_reg_555__3_ ( .D(n16180), .CP(wclk), .Q(ram[11939]) );
  DFF ram_reg_555__2_ ( .D(n16179), .CP(wclk), .Q(ram[11938]) );
  DFF ram_reg_555__1_ ( .D(n16178), .CP(wclk), .Q(ram[11937]) );
  DFF ram_reg_555__0_ ( .D(n16177), .CP(wclk), .Q(ram[11936]) );
  DFF ram_reg_559__7_ ( .D(n16152), .CP(wclk), .Q(ram[11911]) );
  DFF ram_reg_559__6_ ( .D(n16151), .CP(wclk), .Q(ram[11910]) );
  DFF ram_reg_559__5_ ( .D(n16150), .CP(wclk), .Q(ram[11909]) );
  DFF ram_reg_559__4_ ( .D(n16149), .CP(wclk), .Q(ram[11908]) );
  DFF ram_reg_559__3_ ( .D(n16148), .CP(wclk), .Q(ram[11907]) );
  DFF ram_reg_559__2_ ( .D(n16147), .CP(wclk), .Q(ram[11906]) );
  DFF ram_reg_559__1_ ( .D(n16146), .CP(wclk), .Q(ram[11905]) );
  DFF ram_reg_559__0_ ( .D(n16145), .CP(wclk), .Q(ram[11904]) );
  DFF ram_reg_563__7_ ( .D(n16120), .CP(wclk), .Q(ram[11879]) );
  DFF ram_reg_563__6_ ( .D(n16119), .CP(wclk), .Q(ram[11878]) );
  DFF ram_reg_563__5_ ( .D(n16118), .CP(wclk), .Q(ram[11877]) );
  DFF ram_reg_563__4_ ( .D(n16117), .CP(wclk), .Q(ram[11876]) );
  DFF ram_reg_563__3_ ( .D(n16116), .CP(wclk), .Q(ram[11875]) );
  DFF ram_reg_563__2_ ( .D(n16115), .CP(wclk), .Q(ram[11874]) );
  DFF ram_reg_563__1_ ( .D(n16114), .CP(wclk), .Q(ram[11873]) );
  DFF ram_reg_563__0_ ( .D(n16113), .CP(wclk), .Q(ram[11872]) );
  DFF ram_reg_571__7_ ( .D(n16056), .CP(wclk), .Q(ram[11815]) );
  DFF ram_reg_571__6_ ( .D(n16055), .CP(wclk), .Q(ram[11814]) );
  DFF ram_reg_571__5_ ( .D(n16054), .CP(wclk), .Q(ram[11813]) );
  DFF ram_reg_571__4_ ( .D(n16053), .CP(wclk), .Q(ram[11812]) );
  DFF ram_reg_571__3_ ( .D(n16052), .CP(wclk), .Q(ram[11811]) );
  DFF ram_reg_571__2_ ( .D(n16051), .CP(wclk), .Q(ram[11810]) );
  DFF ram_reg_571__1_ ( .D(n16050), .CP(wclk), .Q(ram[11809]) );
  DFF ram_reg_571__0_ ( .D(n16049), .CP(wclk), .Q(ram[11808]) );
  DFF ram_reg_575__7_ ( .D(n16024), .CP(wclk), .Q(ram[11783]) );
  DFF ram_reg_575__6_ ( .D(n16023), .CP(wclk), .Q(ram[11782]) );
  DFF ram_reg_575__5_ ( .D(n16022), .CP(wclk), .Q(ram[11781]) );
  DFF ram_reg_575__4_ ( .D(n16021), .CP(wclk), .Q(ram[11780]) );
  DFF ram_reg_575__3_ ( .D(n16020), .CP(wclk), .Q(ram[11779]) );
  DFF ram_reg_575__2_ ( .D(n16019), .CP(wclk), .Q(ram[11778]) );
  DFF ram_reg_575__1_ ( .D(n16018), .CP(wclk), .Q(ram[11777]) );
  DFF ram_reg_575__0_ ( .D(n16017), .CP(wclk), .Q(ram[11776]) );
  DFF ram_reg_587__7_ ( .D(n15928), .CP(wclk), .Q(ram[11687]) );
  DFF ram_reg_587__6_ ( .D(n15927), .CP(wclk), .Q(ram[11686]) );
  DFF ram_reg_587__5_ ( .D(n15926), .CP(wclk), .Q(ram[11685]) );
  DFF ram_reg_587__4_ ( .D(n15925), .CP(wclk), .Q(ram[11684]) );
  DFF ram_reg_587__3_ ( .D(n15924), .CP(wclk), .Q(ram[11683]) );
  DFF ram_reg_587__2_ ( .D(n15923), .CP(wclk), .Q(ram[11682]) );
  DFF ram_reg_587__1_ ( .D(n15922), .CP(wclk), .Q(ram[11681]) );
  DFF ram_reg_587__0_ ( .D(n15921), .CP(wclk), .Q(ram[11680]) );
  DFF ram_reg_619__7_ ( .D(n15672), .CP(wclk), .Q(ram[11431]) );
  DFF ram_reg_619__6_ ( .D(n15671), .CP(wclk), .Q(ram[11430]) );
  DFF ram_reg_619__5_ ( .D(n15670), .CP(wclk), .Q(ram[11429]) );
  DFF ram_reg_619__4_ ( .D(n15669), .CP(wclk), .Q(ram[11428]) );
  DFF ram_reg_619__3_ ( .D(n15668), .CP(wclk), .Q(ram[11427]) );
  DFF ram_reg_619__2_ ( .D(n15667), .CP(wclk), .Q(ram[11426]) );
  DFF ram_reg_619__1_ ( .D(n15666), .CP(wclk), .Q(ram[11425]) );
  DFF ram_reg_619__0_ ( .D(n15665), .CP(wclk), .Q(ram[11424]) );
  DFF ram_reg_623__7_ ( .D(n15640), .CP(wclk), .Q(ram[11399]) );
  DFF ram_reg_623__6_ ( .D(n15639), .CP(wclk), .Q(ram[11398]) );
  DFF ram_reg_623__5_ ( .D(n15638), .CP(wclk), .Q(ram[11397]) );
  DFF ram_reg_623__4_ ( .D(n15637), .CP(wclk), .Q(ram[11396]) );
  DFF ram_reg_623__3_ ( .D(n15636), .CP(wclk), .Q(ram[11395]) );
  DFF ram_reg_623__2_ ( .D(n15635), .CP(wclk), .Q(ram[11394]) );
  DFF ram_reg_623__1_ ( .D(n15634), .CP(wclk), .Q(ram[11393]) );
  DFF ram_reg_623__0_ ( .D(n15633), .CP(wclk), .Q(ram[11392]) );
  DFF ram_reg_635__7_ ( .D(n15544), .CP(wclk), .Q(ram[11303]) );
  DFF ram_reg_635__6_ ( .D(n15543), .CP(wclk), .Q(ram[11302]) );
  DFF ram_reg_635__5_ ( .D(n15542), .CP(wclk), .Q(ram[11301]) );
  DFF ram_reg_635__4_ ( .D(n15541), .CP(wclk), .Q(ram[11300]) );
  DFF ram_reg_635__3_ ( .D(n15540), .CP(wclk), .Q(ram[11299]) );
  DFF ram_reg_635__2_ ( .D(n15539), .CP(wclk), .Q(ram[11298]) );
  DFF ram_reg_635__1_ ( .D(n15538), .CP(wclk), .Q(ram[11297]) );
  DFF ram_reg_635__0_ ( .D(n15537), .CP(wclk), .Q(ram[11296]) );
  DFF ram_reg_639__7_ ( .D(n15512), .CP(wclk), .Q(ram[11271]) );
  DFF ram_reg_639__6_ ( .D(n15511), .CP(wclk), .Q(ram[11270]) );
  DFF ram_reg_639__5_ ( .D(n15510), .CP(wclk), .Q(ram[11269]) );
  DFF ram_reg_639__4_ ( .D(n15509), .CP(wclk), .Q(ram[11268]) );
  DFF ram_reg_639__3_ ( .D(n15508), .CP(wclk), .Q(ram[11267]) );
  DFF ram_reg_639__2_ ( .D(n15507), .CP(wclk), .Q(ram[11266]) );
  DFF ram_reg_639__1_ ( .D(n15506), .CP(wclk), .Q(ram[11265]) );
  DFF ram_reg_639__0_ ( .D(n15505), .CP(wclk), .Q(ram[11264]) );
  DFF ram_reg_643__7_ ( .D(n15480), .CP(wclk), .Q(ram[11239]) );
  DFF ram_reg_643__6_ ( .D(n15479), .CP(wclk), .Q(ram[11238]) );
  DFF ram_reg_643__5_ ( .D(n15478), .CP(wclk), .Q(ram[11237]) );
  DFF ram_reg_643__4_ ( .D(n15477), .CP(wclk), .Q(ram[11236]) );
  DFF ram_reg_643__3_ ( .D(n15476), .CP(wclk), .Q(ram[11235]) );
  DFF ram_reg_643__2_ ( .D(n15475), .CP(wclk), .Q(ram[11234]) );
  DFF ram_reg_643__1_ ( .D(n15474), .CP(wclk), .Q(ram[11233]) );
  DFF ram_reg_643__0_ ( .D(n15473), .CP(wclk), .Q(ram[11232]) );
  DFF ram_reg_647__7_ ( .D(n15448), .CP(wclk), .Q(ram[11207]) );
  DFF ram_reg_647__6_ ( .D(n15447), .CP(wclk), .Q(ram[11206]) );
  DFF ram_reg_647__5_ ( .D(n15446), .CP(wclk), .Q(ram[11205]) );
  DFF ram_reg_647__4_ ( .D(n15445), .CP(wclk), .Q(ram[11204]) );
  DFF ram_reg_647__3_ ( .D(n15444), .CP(wclk), .Q(ram[11203]) );
  DFF ram_reg_647__2_ ( .D(n15443), .CP(wclk), .Q(ram[11202]) );
  DFF ram_reg_647__1_ ( .D(n15442), .CP(wclk), .Q(ram[11201]) );
  DFF ram_reg_647__0_ ( .D(n15441), .CP(wclk), .Q(ram[11200]) );
  DFF ram_reg_651__7_ ( .D(n15416), .CP(wclk), .Q(ram[11175]) );
  DFF ram_reg_651__6_ ( .D(n15415), .CP(wclk), .Q(ram[11174]) );
  DFF ram_reg_651__5_ ( .D(n15414), .CP(wclk), .Q(ram[11173]) );
  DFF ram_reg_651__4_ ( .D(n15413), .CP(wclk), .Q(ram[11172]) );
  DFF ram_reg_651__3_ ( .D(n15412), .CP(wclk), .Q(ram[11171]) );
  DFF ram_reg_651__2_ ( .D(n15411), .CP(wclk), .Q(ram[11170]) );
  DFF ram_reg_651__1_ ( .D(n15410), .CP(wclk), .Q(ram[11169]) );
  DFF ram_reg_651__0_ ( .D(n15409), .CP(wclk), .Q(ram[11168]) );
  DFF ram_reg_655__7_ ( .D(n15384), .CP(wclk), .Q(ram[11143]) );
  DFF ram_reg_655__6_ ( .D(n15383), .CP(wclk), .Q(ram[11142]) );
  DFF ram_reg_655__5_ ( .D(n15382), .CP(wclk), .Q(ram[11141]) );
  DFF ram_reg_655__4_ ( .D(n15381), .CP(wclk), .Q(ram[11140]) );
  DFF ram_reg_655__3_ ( .D(n15380), .CP(wclk), .Q(ram[11139]) );
  DFF ram_reg_655__2_ ( .D(n15379), .CP(wclk), .Q(ram[11138]) );
  DFF ram_reg_655__1_ ( .D(n15378), .CP(wclk), .Q(ram[11137]) );
  DFF ram_reg_655__0_ ( .D(n15377), .CP(wclk), .Q(ram[11136]) );
  DFF ram_reg_659__7_ ( .D(n15352), .CP(wclk), .Q(ram[11111]) );
  DFF ram_reg_659__6_ ( .D(n15351), .CP(wclk), .Q(ram[11110]) );
  DFF ram_reg_659__5_ ( .D(n15350), .CP(wclk), .Q(ram[11109]) );
  DFF ram_reg_659__4_ ( .D(n15349), .CP(wclk), .Q(ram[11108]) );
  DFF ram_reg_659__3_ ( .D(n15348), .CP(wclk), .Q(ram[11107]) );
  DFF ram_reg_659__2_ ( .D(n15347), .CP(wclk), .Q(ram[11106]) );
  DFF ram_reg_659__1_ ( .D(n15346), .CP(wclk), .Q(ram[11105]) );
  DFF ram_reg_659__0_ ( .D(n15345), .CP(wclk), .Q(ram[11104]) );
  DFF ram_reg_667__7_ ( .D(n15288), .CP(wclk), .Q(ram[11047]) );
  DFF ram_reg_667__6_ ( .D(n15287), .CP(wclk), .Q(ram[11046]) );
  DFF ram_reg_667__5_ ( .D(n15286), .CP(wclk), .Q(ram[11045]) );
  DFF ram_reg_667__4_ ( .D(n15285), .CP(wclk), .Q(ram[11044]) );
  DFF ram_reg_667__3_ ( .D(n15284), .CP(wclk), .Q(ram[11043]) );
  DFF ram_reg_667__2_ ( .D(n15283), .CP(wclk), .Q(ram[11042]) );
  DFF ram_reg_667__1_ ( .D(n15282), .CP(wclk), .Q(ram[11041]) );
  DFF ram_reg_667__0_ ( .D(n15281), .CP(wclk), .Q(ram[11040]) );
  DFF ram_reg_671__7_ ( .D(n15256), .CP(wclk), .Q(ram[11015]) );
  DFF ram_reg_671__6_ ( .D(n15255), .CP(wclk), .Q(ram[11014]) );
  DFF ram_reg_671__5_ ( .D(n15254), .CP(wclk), .Q(ram[11013]) );
  DFF ram_reg_671__4_ ( .D(n15253), .CP(wclk), .Q(ram[11012]) );
  DFF ram_reg_671__3_ ( .D(n15252), .CP(wclk), .Q(ram[11011]) );
  DFF ram_reg_671__2_ ( .D(n15251), .CP(wclk), .Q(ram[11010]) );
  DFF ram_reg_671__1_ ( .D(n15250), .CP(wclk), .Q(ram[11009]) );
  DFF ram_reg_671__0_ ( .D(n15249), .CP(wclk), .Q(ram[11008]) );
  DFF ram_reg_675__7_ ( .D(n15224), .CP(wclk), .Q(ram[10983]) );
  DFF ram_reg_675__6_ ( .D(n15223), .CP(wclk), .Q(ram[10982]) );
  DFF ram_reg_675__5_ ( .D(n15222), .CP(wclk), .Q(ram[10981]) );
  DFF ram_reg_675__4_ ( .D(n15221), .CP(wclk), .Q(ram[10980]) );
  DFF ram_reg_675__3_ ( .D(n15220), .CP(wclk), .Q(ram[10979]) );
  DFF ram_reg_675__2_ ( .D(n15219), .CP(wclk), .Q(ram[10978]) );
  DFF ram_reg_675__1_ ( .D(n15218), .CP(wclk), .Q(ram[10977]) );
  DFF ram_reg_675__0_ ( .D(n15217), .CP(wclk), .Q(ram[10976]) );
  DFF ram_reg_679__7_ ( .D(n15192), .CP(wclk), .Q(ram[10951]) );
  DFF ram_reg_679__6_ ( .D(n15191), .CP(wclk), .Q(ram[10950]) );
  DFF ram_reg_679__5_ ( .D(n15190), .CP(wclk), .Q(ram[10949]) );
  DFF ram_reg_679__4_ ( .D(n15189), .CP(wclk), .Q(ram[10948]) );
  DFF ram_reg_679__3_ ( .D(n15188), .CP(wclk), .Q(ram[10947]) );
  DFF ram_reg_679__2_ ( .D(n15187), .CP(wclk), .Q(ram[10946]) );
  DFF ram_reg_679__1_ ( .D(n15186), .CP(wclk), .Q(ram[10945]) );
  DFF ram_reg_679__0_ ( .D(n15185), .CP(wclk), .Q(ram[10944]) );
  DFF ram_reg_683__7_ ( .D(n15160), .CP(wclk), .Q(ram[10919]) );
  DFF ram_reg_683__6_ ( .D(n15159), .CP(wclk), .Q(ram[10918]) );
  DFF ram_reg_683__5_ ( .D(n15158), .CP(wclk), .Q(ram[10917]) );
  DFF ram_reg_683__4_ ( .D(n15157), .CP(wclk), .Q(ram[10916]) );
  DFF ram_reg_683__3_ ( .D(n15156), .CP(wclk), .Q(ram[10915]) );
  DFF ram_reg_683__2_ ( .D(n15155), .CP(wclk), .Q(ram[10914]) );
  DFF ram_reg_683__1_ ( .D(n15154), .CP(wclk), .Q(ram[10913]) );
  DFF ram_reg_683__0_ ( .D(n15153), .CP(wclk), .Q(ram[10912]) );
  DFF ram_reg_687__7_ ( .D(n15128), .CP(wclk), .Q(ram[10887]) );
  DFF ram_reg_687__6_ ( .D(n15127), .CP(wclk), .Q(ram[10886]) );
  DFF ram_reg_687__5_ ( .D(n15126), .CP(wclk), .Q(ram[10885]) );
  DFF ram_reg_687__4_ ( .D(n15125), .CP(wclk), .Q(ram[10884]) );
  DFF ram_reg_687__3_ ( .D(n15124), .CP(wclk), .Q(ram[10883]) );
  DFF ram_reg_687__2_ ( .D(n15123), .CP(wclk), .Q(ram[10882]) );
  DFF ram_reg_687__1_ ( .D(n15122), .CP(wclk), .Q(ram[10881]) );
  DFF ram_reg_687__0_ ( .D(n15121), .CP(wclk), .Q(ram[10880]) );
  DFF ram_reg_691__7_ ( .D(n15096), .CP(wclk), .Q(ram[10855]) );
  DFF ram_reg_691__6_ ( .D(n15095), .CP(wclk), .Q(ram[10854]) );
  DFF ram_reg_691__5_ ( .D(n15094), .CP(wclk), .Q(ram[10853]) );
  DFF ram_reg_691__4_ ( .D(n15093), .CP(wclk), .Q(ram[10852]) );
  DFF ram_reg_691__3_ ( .D(n15092), .CP(wclk), .Q(ram[10851]) );
  DFF ram_reg_691__2_ ( .D(n15091), .CP(wclk), .Q(ram[10850]) );
  DFF ram_reg_691__1_ ( .D(n15090), .CP(wclk), .Q(ram[10849]) );
  DFF ram_reg_691__0_ ( .D(n15089), .CP(wclk), .Q(ram[10848]) );
  DFF ram_reg_695__7_ ( .D(n15064), .CP(wclk), .Q(ram[10823]) );
  DFF ram_reg_695__6_ ( .D(n15063), .CP(wclk), .Q(ram[10822]) );
  DFF ram_reg_695__5_ ( .D(n15062), .CP(wclk), .Q(ram[10821]) );
  DFF ram_reg_695__4_ ( .D(n15061), .CP(wclk), .Q(ram[10820]) );
  DFF ram_reg_695__3_ ( .D(n15060), .CP(wclk), .Q(ram[10819]) );
  DFF ram_reg_695__2_ ( .D(n15059), .CP(wclk), .Q(ram[10818]) );
  DFF ram_reg_695__1_ ( .D(n15058), .CP(wclk), .Q(ram[10817]) );
  DFF ram_reg_695__0_ ( .D(n15057), .CP(wclk), .Q(ram[10816]) );
  DFF ram_reg_699__7_ ( .D(n15032), .CP(wclk), .Q(ram[10791]) );
  DFF ram_reg_699__6_ ( .D(n15031), .CP(wclk), .Q(ram[10790]) );
  DFF ram_reg_699__5_ ( .D(n15030), .CP(wclk), .Q(ram[10789]) );
  DFF ram_reg_699__4_ ( .D(n15029), .CP(wclk), .Q(ram[10788]) );
  DFF ram_reg_699__3_ ( .D(n15028), .CP(wclk), .Q(ram[10787]) );
  DFF ram_reg_699__2_ ( .D(n15027), .CP(wclk), .Q(ram[10786]) );
  DFF ram_reg_699__1_ ( .D(n15026), .CP(wclk), .Q(ram[10785]) );
  DFF ram_reg_699__0_ ( .D(n15025), .CP(wclk), .Q(ram[10784]) );
  DFF ram_reg_703__7_ ( .D(n15000), .CP(wclk), .Q(ram[10759]) );
  DFF ram_reg_703__6_ ( .D(n14999), .CP(wclk), .Q(ram[10758]) );
  DFF ram_reg_703__5_ ( .D(n14998), .CP(wclk), .Q(ram[10757]) );
  DFF ram_reg_703__4_ ( .D(n14997), .CP(wclk), .Q(ram[10756]) );
  DFF ram_reg_703__3_ ( .D(n14996), .CP(wclk), .Q(ram[10755]) );
  DFF ram_reg_703__2_ ( .D(n14995), .CP(wclk), .Q(ram[10754]) );
  DFF ram_reg_703__1_ ( .D(n14994), .CP(wclk), .Q(ram[10753]) );
  DFF ram_reg_703__0_ ( .D(n14993), .CP(wclk), .Q(ram[10752]) );
  DFF ram_reg_707__7_ ( .D(n14968), .CP(wclk), .Q(ram[10727]) );
  DFF ram_reg_707__6_ ( .D(n14967), .CP(wclk), .Q(ram[10726]) );
  DFF ram_reg_707__5_ ( .D(n14966), .CP(wclk), .Q(ram[10725]) );
  DFF ram_reg_707__4_ ( .D(n14965), .CP(wclk), .Q(ram[10724]) );
  DFF ram_reg_707__3_ ( .D(n14964), .CP(wclk), .Q(ram[10723]) );
  DFF ram_reg_707__2_ ( .D(n14963), .CP(wclk), .Q(ram[10722]) );
  DFF ram_reg_707__1_ ( .D(n14962), .CP(wclk), .Q(ram[10721]) );
  DFF ram_reg_707__0_ ( .D(n14961), .CP(wclk), .Q(ram[10720]) );
  DFF ram_reg_715__7_ ( .D(n14904), .CP(wclk), .Q(ram[10663]) );
  DFF ram_reg_715__6_ ( .D(n14903), .CP(wclk), .Q(ram[10662]) );
  DFF ram_reg_715__5_ ( .D(n14902), .CP(wclk), .Q(ram[10661]) );
  DFF ram_reg_715__4_ ( .D(n14901), .CP(wclk), .Q(ram[10660]) );
  DFF ram_reg_715__3_ ( .D(n14900), .CP(wclk), .Q(ram[10659]) );
  DFF ram_reg_715__2_ ( .D(n14899), .CP(wclk), .Q(ram[10658]) );
  DFF ram_reg_715__1_ ( .D(n14898), .CP(wclk), .Q(ram[10657]) );
  DFF ram_reg_715__0_ ( .D(n14897), .CP(wclk), .Q(ram[10656]) );
  DFF ram_reg_719__7_ ( .D(n14872), .CP(wclk), .Q(ram[10631]) );
  DFF ram_reg_719__6_ ( .D(n14871), .CP(wclk), .Q(ram[10630]) );
  DFF ram_reg_719__5_ ( .D(n14870), .CP(wclk), .Q(ram[10629]) );
  DFF ram_reg_719__4_ ( .D(n14869), .CP(wclk), .Q(ram[10628]) );
  DFF ram_reg_719__3_ ( .D(n14868), .CP(wclk), .Q(ram[10627]) );
  DFF ram_reg_719__2_ ( .D(n14867), .CP(wclk), .Q(ram[10626]) );
  DFF ram_reg_719__1_ ( .D(n14866), .CP(wclk), .Q(ram[10625]) );
  DFF ram_reg_719__0_ ( .D(n14865), .CP(wclk), .Q(ram[10624]) );
  DFF ram_reg_723__7_ ( .D(n14840), .CP(wclk), .Q(ram[10599]) );
  DFF ram_reg_723__6_ ( .D(n14839), .CP(wclk), .Q(ram[10598]) );
  DFF ram_reg_723__5_ ( .D(n14838), .CP(wclk), .Q(ram[10597]) );
  DFF ram_reg_723__4_ ( .D(n14837), .CP(wclk), .Q(ram[10596]) );
  DFF ram_reg_723__3_ ( .D(n14836), .CP(wclk), .Q(ram[10595]) );
  DFF ram_reg_723__2_ ( .D(n14835), .CP(wclk), .Q(ram[10594]) );
  DFF ram_reg_723__1_ ( .D(n14834), .CP(wclk), .Q(ram[10593]) );
  DFF ram_reg_723__0_ ( .D(n14833), .CP(wclk), .Q(ram[10592]) );
  DFF ram_reg_731__7_ ( .D(n14776), .CP(wclk), .Q(ram[10535]) );
  DFF ram_reg_731__6_ ( .D(n14775), .CP(wclk), .Q(ram[10534]) );
  DFF ram_reg_731__5_ ( .D(n14774), .CP(wclk), .Q(ram[10533]) );
  DFF ram_reg_731__4_ ( .D(n14773), .CP(wclk), .Q(ram[10532]) );
  DFF ram_reg_731__3_ ( .D(n14772), .CP(wclk), .Q(ram[10531]) );
  DFF ram_reg_731__2_ ( .D(n14771), .CP(wclk), .Q(ram[10530]) );
  DFF ram_reg_731__1_ ( .D(n14770), .CP(wclk), .Q(ram[10529]) );
  DFF ram_reg_731__0_ ( .D(n14769), .CP(wclk), .Q(ram[10528]) );
  DFF ram_reg_735__7_ ( .D(n14744), .CP(wclk), .Q(ram[10503]) );
  DFF ram_reg_735__6_ ( .D(n14743), .CP(wclk), .Q(ram[10502]) );
  DFF ram_reg_735__5_ ( .D(n14742), .CP(wclk), .Q(ram[10501]) );
  DFF ram_reg_735__4_ ( .D(n14741), .CP(wclk), .Q(ram[10500]) );
  DFF ram_reg_735__3_ ( .D(n14740), .CP(wclk), .Q(ram[10499]) );
  DFF ram_reg_735__2_ ( .D(n14739), .CP(wclk), .Q(ram[10498]) );
  DFF ram_reg_735__1_ ( .D(n14738), .CP(wclk), .Q(ram[10497]) );
  DFF ram_reg_735__0_ ( .D(n14737), .CP(wclk), .Q(ram[10496]) );
  DFF ram_reg_739__7_ ( .D(n14712), .CP(wclk), .Q(ram[10471]) );
  DFF ram_reg_739__6_ ( .D(n14711), .CP(wclk), .Q(ram[10470]) );
  DFF ram_reg_739__5_ ( .D(n14710), .CP(wclk), .Q(ram[10469]) );
  DFF ram_reg_739__4_ ( .D(n14709), .CP(wclk), .Q(ram[10468]) );
  DFF ram_reg_739__3_ ( .D(n14708), .CP(wclk), .Q(ram[10467]) );
  DFF ram_reg_739__2_ ( .D(n14707), .CP(wclk), .Q(ram[10466]) );
  DFF ram_reg_739__1_ ( .D(n14706), .CP(wclk), .Q(ram[10465]) );
  DFF ram_reg_739__0_ ( .D(n14705), .CP(wclk), .Q(ram[10464]) );
  DFF ram_reg_743__7_ ( .D(n14680), .CP(wclk), .Q(ram[10439]) );
  DFF ram_reg_743__6_ ( .D(n14679), .CP(wclk), .Q(ram[10438]) );
  DFF ram_reg_743__5_ ( .D(n14678), .CP(wclk), .Q(ram[10437]) );
  DFF ram_reg_743__4_ ( .D(n14677), .CP(wclk), .Q(ram[10436]) );
  DFF ram_reg_743__3_ ( .D(n14676), .CP(wclk), .Q(ram[10435]) );
  DFF ram_reg_743__2_ ( .D(n14675), .CP(wclk), .Q(ram[10434]) );
  DFF ram_reg_743__1_ ( .D(n14674), .CP(wclk), .Q(ram[10433]) );
  DFF ram_reg_743__0_ ( .D(n14673), .CP(wclk), .Q(ram[10432]) );
  DFF ram_reg_747__7_ ( .D(n14648), .CP(wclk), .Q(ram[10407]) );
  DFF ram_reg_747__6_ ( .D(n14647), .CP(wclk), .Q(ram[10406]) );
  DFF ram_reg_747__5_ ( .D(n14646), .CP(wclk), .Q(ram[10405]) );
  DFF ram_reg_747__4_ ( .D(n14645), .CP(wclk), .Q(ram[10404]) );
  DFF ram_reg_747__3_ ( .D(n14644), .CP(wclk), .Q(ram[10403]) );
  DFF ram_reg_747__2_ ( .D(n14643), .CP(wclk), .Q(ram[10402]) );
  DFF ram_reg_747__1_ ( .D(n14642), .CP(wclk), .Q(ram[10401]) );
  DFF ram_reg_747__0_ ( .D(n14641), .CP(wclk), .Q(ram[10400]) );
  DFF ram_reg_751__7_ ( .D(n14616), .CP(wclk), .Q(ram[10375]) );
  DFF ram_reg_751__6_ ( .D(n14615), .CP(wclk), .Q(ram[10374]) );
  DFF ram_reg_751__5_ ( .D(n14614), .CP(wclk), .Q(ram[10373]) );
  DFF ram_reg_751__4_ ( .D(n14613), .CP(wclk), .Q(ram[10372]) );
  DFF ram_reg_751__3_ ( .D(n14612), .CP(wclk), .Q(ram[10371]) );
  DFF ram_reg_751__2_ ( .D(n14611), .CP(wclk), .Q(ram[10370]) );
  DFF ram_reg_751__1_ ( .D(n14610), .CP(wclk), .Q(ram[10369]) );
  DFF ram_reg_751__0_ ( .D(n14609), .CP(wclk), .Q(ram[10368]) );
  DFF ram_reg_755__7_ ( .D(n14584), .CP(wclk), .Q(ram[10343]) );
  DFF ram_reg_755__6_ ( .D(n14583), .CP(wclk), .Q(ram[10342]) );
  DFF ram_reg_755__5_ ( .D(n14582), .CP(wclk), .Q(ram[10341]) );
  DFF ram_reg_755__4_ ( .D(n14581), .CP(wclk), .Q(ram[10340]) );
  DFF ram_reg_755__3_ ( .D(n14580), .CP(wclk), .Q(ram[10339]) );
  DFF ram_reg_755__2_ ( .D(n14579), .CP(wclk), .Q(ram[10338]) );
  DFF ram_reg_755__1_ ( .D(n14578), .CP(wclk), .Q(ram[10337]) );
  DFF ram_reg_755__0_ ( .D(n14577), .CP(wclk), .Q(ram[10336]) );
  DFF ram_reg_759__7_ ( .D(n14552), .CP(wclk), .Q(ram[10311]) );
  DFF ram_reg_759__6_ ( .D(n14551), .CP(wclk), .Q(ram[10310]) );
  DFF ram_reg_759__5_ ( .D(n14550), .CP(wclk), .Q(ram[10309]) );
  DFF ram_reg_759__4_ ( .D(n14549), .CP(wclk), .Q(ram[10308]) );
  DFF ram_reg_759__3_ ( .D(n14548), .CP(wclk), .Q(ram[10307]) );
  DFF ram_reg_759__2_ ( .D(n14547), .CP(wclk), .Q(ram[10306]) );
  DFF ram_reg_759__1_ ( .D(n14546), .CP(wclk), .Q(ram[10305]) );
  DFF ram_reg_759__0_ ( .D(n14545), .CP(wclk), .Q(ram[10304]) );
  DFF ram_reg_763__7_ ( .D(n14520), .CP(wclk), .Q(ram[10279]) );
  DFF ram_reg_763__6_ ( .D(n14519), .CP(wclk), .Q(ram[10278]) );
  DFF ram_reg_763__5_ ( .D(n14518), .CP(wclk), .Q(ram[10277]) );
  DFF ram_reg_763__4_ ( .D(n14517), .CP(wclk), .Q(ram[10276]) );
  DFF ram_reg_763__3_ ( .D(n14516), .CP(wclk), .Q(ram[10275]) );
  DFF ram_reg_763__2_ ( .D(n14515), .CP(wclk), .Q(ram[10274]) );
  DFF ram_reg_763__1_ ( .D(n14514), .CP(wclk), .Q(ram[10273]) );
  DFF ram_reg_763__0_ ( .D(n14513), .CP(wclk), .Q(ram[10272]) );
  DFF ram_reg_767__7_ ( .D(n14488), .CP(wclk), .Q(ram[10247]) );
  DFF ram_reg_767__6_ ( .D(n14487), .CP(wclk), .Q(ram[10246]) );
  DFF ram_reg_767__5_ ( .D(n14486), .CP(wclk), .Q(ram[10245]) );
  DFF ram_reg_767__4_ ( .D(n14485), .CP(wclk), .Q(ram[10244]) );
  DFF ram_reg_767__3_ ( .D(n14484), .CP(wclk), .Q(ram[10243]) );
  DFF ram_reg_767__2_ ( .D(n14483), .CP(wclk), .Q(ram[10242]) );
  DFF ram_reg_767__1_ ( .D(n14482), .CP(wclk), .Q(ram[10241]) );
  DFF ram_reg_767__0_ ( .D(n14481), .CP(wclk), .Q(ram[10240]) );
  DFF ram_reg_771__7_ ( .D(n14456), .CP(wclk), .Q(ram[10215]) );
  DFF ram_reg_771__6_ ( .D(n14455), .CP(wclk), .Q(ram[10214]) );
  DFF ram_reg_771__5_ ( .D(n14454), .CP(wclk), .Q(ram[10213]) );
  DFF ram_reg_771__4_ ( .D(n14453), .CP(wclk), .Q(ram[10212]) );
  DFF ram_reg_771__3_ ( .D(n14452), .CP(wclk), .Q(ram[10211]) );
  DFF ram_reg_771__2_ ( .D(n14451), .CP(wclk), .Q(ram[10210]) );
  DFF ram_reg_771__1_ ( .D(n14450), .CP(wclk), .Q(ram[10209]) );
  DFF ram_reg_771__0_ ( .D(n14449), .CP(wclk), .Q(ram[10208]) );
  DFF ram_reg_779__7_ ( .D(n14392), .CP(wclk), .Q(ram[10151]) );
  DFF ram_reg_779__6_ ( .D(n14391), .CP(wclk), .Q(ram[10150]) );
  DFF ram_reg_779__5_ ( .D(n14390), .CP(wclk), .Q(ram[10149]) );
  DFF ram_reg_779__4_ ( .D(n14389), .CP(wclk), .Q(ram[10148]) );
  DFF ram_reg_779__3_ ( .D(n14388), .CP(wclk), .Q(ram[10147]) );
  DFF ram_reg_779__2_ ( .D(n14387), .CP(wclk), .Q(ram[10146]) );
  DFF ram_reg_779__1_ ( .D(n14386), .CP(wclk), .Q(ram[10145]) );
  DFF ram_reg_779__0_ ( .D(n14385), .CP(wclk), .Q(ram[10144]) );
  DFF ram_reg_783__7_ ( .D(n14360), .CP(wclk), .Q(ram[10119]) );
  DFF ram_reg_783__6_ ( .D(n14359), .CP(wclk), .Q(ram[10118]) );
  DFF ram_reg_783__5_ ( .D(n14358), .CP(wclk), .Q(ram[10117]) );
  DFF ram_reg_783__4_ ( .D(n14357), .CP(wclk), .Q(ram[10116]) );
  DFF ram_reg_783__3_ ( .D(n14356), .CP(wclk), .Q(ram[10115]) );
  DFF ram_reg_783__2_ ( .D(n14355), .CP(wclk), .Q(ram[10114]) );
  DFF ram_reg_783__1_ ( .D(n14354), .CP(wclk), .Q(ram[10113]) );
  DFF ram_reg_783__0_ ( .D(n14353), .CP(wclk), .Q(ram[10112]) );
  DFF ram_reg_795__7_ ( .D(n14264), .CP(wclk), .Q(ram[10023]) );
  DFF ram_reg_795__6_ ( .D(n14263), .CP(wclk), .Q(ram[10022]) );
  DFF ram_reg_795__5_ ( .D(n14262), .CP(wclk), .Q(ram[10021]) );
  DFF ram_reg_795__4_ ( .D(n14261), .CP(wclk), .Q(ram[10020]) );
  DFF ram_reg_795__3_ ( .D(n14260), .CP(wclk), .Q(ram[10019]) );
  DFF ram_reg_795__2_ ( .D(n14259), .CP(wclk), .Q(ram[10018]) );
  DFF ram_reg_795__1_ ( .D(n14258), .CP(wclk), .Q(ram[10017]) );
  DFF ram_reg_795__0_ ( .D(n14257), .CP(wclk), .Q(ram[10016]) );
  DFF ram_reg_799__7_ ( .D(n14232), .CP(wclk), .Q(ram[9991]) );
  DFF ram_reg_799__6_ ( .D(n14231), .CP(wclk), .Q(ram[9990]) );
  DFF ram_reg_799__5_ ( .D(n14230), .CP(wclk), .Q(ram[9989]) );
  DFF ram_reg_799__4_ ( .D(n14229), .CP(wclk), .Q(ram[9988]) );
  DFF ram_reg_799__3_ ( .D(n14228), .CP(wclk), .Q(ram[9987]) );
  DFF ram_reg_799__2_ ( .D(n14227), .CP(wclk), .Q(ram[9986]) );
  DFF ram_reg_799__1_ ( .D(n14226), .CP(wclk), .Q(ram[9985]) );
  DFF ram_reg_799__0_ ( .D(n14225), .CP(wclk), .Q(ram[9984]) );
  DFF ram_reg_803__7_ ( .D(n14200), .CP(wclk), .Q(ram[9959]) );
  DFF ram_reg_803__6_ ( .D(n14199), .CP(wclk), .Q(ram[9958]) );
  DFF ram_reg_803__5_ ( .D(n14198), .CP(wclk), .Q(ram[9957]) );
  DFF ram_reg_803__4_ ( .D(n14197), .CP(wclk), .Q(ram[9956]) );
  DFF ram_reg_803__3_ ( .D(n14196), .CP(wclk), .Q(ram[9955]) );
  DFF ram_reg_803__2_ ( .D(n14195), .CP(wclk), .Q(ram[9954]) );
  DFF ram_reg_803__1_ ( .D(n14194), .CP(wclk), .Q(ram[9953]) );
  DFF ram_reg_803__0_ ( .D(n14193), .CP(wclk), .Q(ram[9952]) );
  DFF ram_reg_811__7_ ( .D(n14136), .CP(wclk), .Q(ram[9895]) );
  DFF ram_reg_811__6_ ( .D(n14135), .CP(wclk), .Q(ram[9894]) );
  DFF ram_reg_811__5_ ( .D(n14134), .CP(wclk), .Q(ram[9893]) );
  DFF ram_reg_811__4_ ( .D(n14133), .CP(wclk), .Q(ram[9892]) );
  DFF ram_reg_811__3_ ( .D(n14132), .CP(wclk), .Q(ram[9891]) );
  DFF ram_reg_811__2_ ( .D(n14131), .CP(wclk), .Q(ram[9890]) );
  DFF ram_reg_811__1_ ( .D(n14130), .CP(wclk), .Q(ram[9889]) );
  DFF ram_reg_811__0_ ( .D(n14129), .CP(wclk), .Q(ram[9888]) );
  DFF ram_reg_815__7_ ( .D(n14104), .CP(wclk), .Q(ram[9863]) );
  DFF ram_reg_815__6_ ( .D(n14103), .CP(wclk), .Q(ram[9862]) );
  DFF ram_reg_815__5_ ( .D(n14102), .CP(wclk), .Q(ram[9861]) );
  DFF ram_reg_815__4_ ( .D(n14101), .CP(wclk), .Q(ram[9860]) );
  DFF ram_reg_815__3_ ( .D(n14100), .CP(wclk), .Q(ram[9859]) );
  DFF ram_reg_815__2_ ( .D(n14099), .CP(wclk), .Q(ram[9858]) );
  DFF ram_reg_815__1_ ( .D(n14098), .CP(wclk), .Q(ram[9857]) );
  DFF ram_reg_815__0_ ( .D(n14097), .CP(wclk), .Q(ram[9856]) );
  DFF ram_reg_819__7_ ( .D(n14072), .CP(wclk), .Q(ram[9831]) );
  DFF ram_reg_819__6_ ( .D(n14071), .CP(wclk), .Q(ram[9830]) );
  DFF ram_reg_819__5_ ( .D(n14070), .CP(wclk), .Q(ram[9829]) );
  DFF ram_reg_819__4_ ( .D(n14069), .CP(wclk), .Q(ram[9828]) );
  DFF ram_reg_819__3_ ( .D(n14068), .CP(wclk), .Q(ram[9827]) );
  DFF ram_reg_819__2_ ( .D(n14067), .CP(wclk), .Q(ram[9826]) );
  DFF ram_reg_819__1_ ( .D(n14066), .CP(wclk), .Q(ram[9825]) );
  DFF ram_reg_819__0_ ( .D(n14065), .CP(wclk), .Q(ram[9824]) );
  DFF ram_reg_827__7_ ( .D(n14008), .CP(wclk), .Q(ram[9767]) );
  DFF ram_reg_827__6_ ( .D(n14007), .CP(wclk), .Q(ram[9766]) );
  DFF ram_reg_827__5_ ( .D(n14006), .CP(wclk), .Q(ram[9765]) );
  DFF ram_reg_827__4_ ( .D(n14005), .CP(wclk), .Q(ram[9764]) );
  DFF ram_reg_827__3_ ( .D(n14004), .CP(wclk), .Q(ram[9763]) );
  DFF ram_reg_827__2_ ( .D(n14003), .CP(wclk), .Q(ram[9762]) );
  DFF ram_reg_827__1_ ( .D(n14002), .CP(wclk), .Q(ram[9761]) );
  DFF ram_reg_827__0_ ( .D(n14001), .CP(wclk), .Q(ram[9760]) );
  DFF ram_reg_831__7_ ( .D(n13976), .CP(wclk), .Q(ram[9735]) );
  DFF ram_reg_831__6_ ( .D(n13975), .CP(wclk), .Q(ram[9734]) );
  DFF ram_reg_831__5_ ( .D(n13974), .CP(wclk), .Q(ram[9733]) );
  DFF ram_reg_831__4_ ( .D(n13973), .CP(wclk), .Q(ram[9732]) );
  DFF ram_reg_831__3_ ( .D(n13972), .CP(wclk), .Q(ram[9731]) );
  DFF ram_reg_831__2_ ( .D(n13971), .CP(wclk), .Q(ram[9730]) );
  DFF ram_reg_831__1_ ( .D(n13970), .CP(wclk), .Q(ram[9729]) );
  DFF ram_reg_831__0_ ( .D(n13969), .CP(wclk), .Q(ram[9728]) );
  DFF ram_reg_843__7_ ( .D(n13880), .CP(wclk), .Q(ram[9639]) );
  DFF ram_reg_843__6_ ( .D(n13879), .CP(wclk), .Q(ram[9638]) );
  DFF ram_reg_843__5_ ( .D(n13878), .CP(wclk), .Q(ram[9637]) );
  DFF ram_reg_843__4_ ( .D(n13877), .CP(wclk), .Q(ram[9636]) );
  DFF ram_reg_843__3_ ( .D(n13876), .CP(wclk), .Q(ram[9635]) );
  DFF ram_reg_843__2_ ( .D(n13875), .CP(wclk), .Q(ram[9634]) );
  DFF ram_reg_843__1_ ( .D(n13874), .CP(wclk), .Q(ram[9633]) );
  DFF ram_reg_843__0_ ( .D(n13873), .CP(wclk), .Q(ram[9632]) );
  DFF ram_reg_859__7_ ( .D(n13752), .CP(wclk), .Q(ram[9511]) );
  DFF ram_reg_859__6_ ( .D(n13751), .CP(wclk), .Q(ram[9510]) );
  DFF ram_reg_859__5_ ( .D(n13750), .CP(wclk), .Q(ram[9509]) );
  DFF ram_reg_859__4_ ( .D(n13749), .CP(wclk), .Q(ram[9508]) );
  DFF ram_reg_859__3_ ( .D(n13748), .CP(wclk), .Q(ram[9507]) );
  DFF ram_reg_859__2_ ( .D(n13747), .CP(wclk), .Q(ram[9506]) );
  DFF ram_reg_859__1_ ( .D(n13746), .CP(wclk), .Q(ram[9505]) );
  DFF ram_reg_859__0_ ( .D(n13745), .CP(wclk), .Q(ram[9504]) );
  DFF ram_reg_875__7_ ( .D(n13624), .CP(wclk), .Q(ram[9383]) );
  DFF ram_reg_875__6_ ( .D(n13623), .CP(wclk), .Q(ram[9382]) );
  DFF ram_reg_875__5_ ( .D(n13622), .CP(wclk), .Q(ram[9381]) );
  DFF ram_reg_875__4_ ( .D(n13621), .CP(wclk), .Q(ram[9380]) );
  DFF ram_reg_875__3_ ( .D(n13620), .CP(wclk), .Q(ram[9379]) );
  DFF ram_reg_875__2_ ( .D(n13619), .CP(wclk), .Q(ram[9378]) );
  DFF ram_reg_875__1_ ( .D(n13618), .CP(wclk), .Q(ram[9377]) );
  DFF ram_reg_875__0_ ( .D(n13617), .CP(wclk), .Q(ram[9376]) );
  DFF ram_reg_879__7_ ( .D(n13592), .CP(wclk), .Q(ram[9351]) );
  DFF ram_reg_879__6_ ( .D(n13591), .CP(wclk), .Q(ram[9350]) );
  DFF ram_reg_879__5_ ( .D(n13590), .CP(wclk), .Q(ram[9349]) );
  DFF ram_reg_879__4_ ( .D(n13589), .CP(wclk), .Q(ram[9348]) );
  DFF ram_reg_879__3_ ( .D(n13588), .CP(wclk), .Q(ram[9347]) );
  DFF ram_reg_879__2_ ( .D(n13587), .CP(wclk), .Q(ram[9346]) );
  DFF ram_reg_879__1_ ( .D(n13586), .CP(wclk), .Q(ram[9345]) );
  DFF ram_reg_879__0_ ( .D(n13585), .CP(wclk), .Q(ram[9344]) );
  DFF ram_reg_891__7_ ( .D(n13496), .CP(wclk), .Q(ram[9255]) );
  DFF ram_reg_891__6_ ( .D(n13495), .CP(wclk), .Q(ram[9254]) );
  DFF ram_reg_891__5_ ( .D(n13494), .CP(wclk), .Q(ram[9253]) );
  DFF ram_reg_891__4_ ( .D(n13493), .CP(wclk), .Q(ram[9252]) );
  DFF ram_reg_891__3_ ( .D(n13492), .CP(wclk), .Q(ram[9251]) );
  DFF ram_reg_891__2_ ( .D(n13491), .CP(wclk), .Q(ram[9250]) );
  DFF ram_reg_891__1_ ( .D(n13490), .CP(wclk), .Q(ram[9249]) );
  DFF ram_reg_891__0_ ( .D(n13489), .CP(wclk), .Q(ram[9248]) );
  DFF ram_reg_895__7_ ( .D(n13464), .CP(wclk), .Q(ram[9223]) );
  DFF ram_reg_895__6_ ( .D(n13463), .CP(wclk), .Q(ram[9222]) );
  DFF ram_reg_895__5_ ( .D(n13462), .CP(wclk), .Q(ram[9221]) );
  DFF ram_reg_895__4_ ( .D(n13461), .CP(wclk), .Q(ram[9220]) );
  DFF ram_reg_895__3_ ( .D(n13460), .CP(wclk), .Q(ram[9219]) );
  DFF ram_reg_895__2_ ( .D(n13459), .CP(wclk), .Q(ram[9218]) );
  DFF ram_reg_895__1_ ( .D(n13458), .CP(wclk), .Q(ram[9217]) );
  DFF ram_reg_895__0_ ( .D(n13457), .CP(wclk), .Q(ram[9216]) );
  DFF ram_reg_899__7_ ( .D(n13432), .CP(wclk), .Q(ram[9191]) );
  DFF ram_reg_899__6_ ( .D(n13431), .CP(wclk), .Q(ram[9190]) );
  DFF ram_reg_899__5_ ( .D(n13430), .CP(wclk), .Q(ram[9189]) );
  DFF ram_reg_899__4_ ( .D(n13429), .CP(wclk), .Q(ram[9188]) );
  DFF ram_reg_899__3_ ( .D(n13428), .CP(wclk), .Q(ram[9187]) );
  DFF ram_reg_899__2_ ( .D(n13427), .CP(wclk), .Q(ram[9186]) );
  DFF ram_reg_899__1_ ( .D(n13426), .CP(wclk), .Q(ram[9185]) );
  DFF ram_reg_899__0_ ( .D(n13425), .CP(wclk), .Q(ram[9184]) );
  DFF ram_reg_903__7_ ( .D(n13400), .CP(wclk), .Q(ram[9159]) );
  DFF ram_reg_903__6_ ( .D(n13399), .CP(wclk), .Q(ram[9158]) );
  DFF ram_reg_903__5_ ( .D(n13398), .CP(wclk), .Q(ram[9157]) );
  DFF ram_reg_903__4_ ( .D(n13397), .CP(wclk), .Q(ram[9156]) );
  DFF ram_reg_903__3_ ( .D(n13396), .CP(wclk), .Q(ram[9155]) );
  DFF ram_reg_903__2_ ( .D(n13395), .CP(wclk), .Q(ram[9154]) );
  DFF ram_reg_903__1_ ( .D(n13394), .CP(wclk), .Q(ram[9153]) );
  DFF ram_reg_903__0_ ( .D(n13393), .CP(wclk), .Q(ram[9152]) );
  DFF ram_reg_907__7_ ( .D(n13368), .CP(wclk), .Q(ram[9127]) );
  DFF ram_reg_907__6_ ( .D(n13367), .CP(wclk), .Q(ram[9126]) );
  DFF ram_reg_907__5_ ( .D(n13366), .CP(wclk), .Q(ram[9125]) );
  DFF ram_reg_907__4_ ( .D(n13365), .CP(wclk), .Q(ram[9124]) );
  DFF ram_reg_907__3_ ( .D(n13364), .CP(wclk), .Q(ram[9123]) );
  DFF ram_reg_907__2_ ( .D(n13363), .CP(wclk), .Q(ram[9122]) );
  DFF ram_reg_907__1_ ( .D(n13362), .CP(wclk), .Q(ram[9121]) );
  DFF ram_reg_907__0_ ( .D(n13361), .CP(wclk), .Q(ram[9120]) );
  DFF ram_reg_911__7_ ( .D(n13336), .CP(wclk), .Q(ram[9095]) );
  DFF ram_reg_911__6_ ( .D(n13335), .CP(wclk), .Q(ram[9094]) );
  DFF ram_reg_911__5_ ( .D(n13334), .CP(wclk), .Q(ram[9093]) );
  DFF ram_reg_911__4_ ( .D(n13333), .CP(wclk), .Q(ram[9092]) );
  DFF ram_reg_911__3_ ( .D(n13332), .CP(wclk), .Q(ram[9091]) );
  DFF ram_reg_911__2_ ( .D(n13331), .CP(wclk), .Q(ram[9090]) );
  DFF ram_reg_911__1_ ( .D(n13330), .CP(wclk), .Q(ram[9089]) );
  DFF ram_reg_911__0_ ( .D(n13329), .CP(wclk), .Q(ram[9088]) );
  DFF ram_reg_915__7_ ( .D(n13304), .CP(wclk), .Q(ram[9063]) );
  DFF ram_reg_915__6_ ( .D(n13303), .CP(wclk), .Q(ram[9062]) );
  DFF ram_reg_915__5_ ( .D(n13302), .CP(wclk), .Q(ram[9061]) );
  DFF ram_reg_915__4_ ( .D(n13301), .CP(wclk), .Q(ram[9060]) );
  DFF ram_reg_915__3_ ( .D(n13300), .CP(wclk), .Q(ram[9059]) );
  DFF ram_reg_915__2_ ( .D(n13299), .CP(wclk), .Q(ram[9058]) );
  DFF ram_reg_915__1_ ( .D(n13298), .CP(wclk), .Q(ram[9057]) );
  DFF ram_reg_915__0_ ( .D(n13297), .CP(wclk), .Q(ram[9056]) );
  DFF ram_reg_919__7_ ( .D(n13272), .CP(wclk), .Q(ram[9031]) );
  DFF ram_reg_919__6_ ( .D(n13271), .CP(wclk), .Q(ram[9030]) );
  DFF ram_reg_919__5_ ( .D(n13270), .CP(wclk), .Q(ram[9029]) );
  DFF ram_reg_919__4_ ( .D(n13269), .CP(wclk), .Q(ram[9028]) );
  DFF ram_reg_919__3_ ( .D(n13268), .CP(wclk), .Q(ram[9027]) );
  DFF ram_reg_919__2_ ( .D(n13267), .CP(wclk), .Q(ram[9026]) );
  DFF ram_reg_919__1_ ( .D(n13266), .CP(wclk), .Q(ram[9025]) );
  DFF ram_reg_919__0_ ( .D(n13265), .CP(wclk), .Q(ram[9024]) );
  DFF ram_reg_923__7_ ( .D(n13240), .CP(wclk), .Q(ram[8999]) );
  DFF ram_reg_923__6_ ( .D(n13239), .CP(wclk), .Q(ram[8998]) );
  DFF ram_reg_923__5_ ( .D(n13238), .CP(wclk), .Q(ram[8997]) );
  DFF ram_reg_923__4_ ( .D(n13237), .CP(wclk), .Q(ram[8996]) );
  DFF ram_reg_923__3_ ( .D(n13236), .CP(wclk), .Q(ram[8995]) );
  DFF ram_reg_923__2_ ( .D(n13235), .CP(wclk), .Q(ram[8994]) );
  DFF ram_reg_923__1_ ( .D(n13234), .CP(wclk), .Q(ram[8993]) );
  DFF ram_reg_923__0_ ( .D(n13233), .CP(wclk), .Q(ram[8992]) );
  DFF ram_reg_927__7_ ( .D(n13208), .CP(wclk), .Q(ram[8967]) );
  DFF ram_reg_927__6_ ( .D(n13207), .CP(wclk), .Q(ram[8966]) );
  DFF ram_reg_927__5_ ( .D(n13206), .CP(wclk), .Q(ram[8965]) );
  DFF ram_reg_927__4_ ( .D(n13205), .CP(wclk), .Q(ram[8964]) );
  DFF ram_reg_927__3_ ( .D(n13204), .CP(wclk), .Q(ram[8963]) );
  DFF ram_reg_927__2_ ( .D(n13203), .CP(wclk), .Q(ram[8962]) );
  DFF ram_reg_927__1_ ( .D(n13202), .CP(wclk), .Q(ram[8961]) );
  DFF ram_reg_927__0_ ( .D(n13201), .CP(wclk), .Q(ram[8960]) );
  DFF ram_reg_931__7_ ( .D(n13176), .CP(wclk), .Q(ram[8935]) );
  DFF ram_reg_931__6_ ( .D(n13175), .CP(wclk), .Q(ram[8934]) );
  DFF ram_reg_931__5_ ( .D(n13174), .CP(wclk), .Q(ram[8933]) );
  DFF ram_reg_931__4_ ( .D(n13173), .CP(wclk), .Q(ram[8932]) );
  DFF ram_reg_931__3_ ( .D(n13172), .CP(wclk), .Q(ram[8931]) );
  DFF ram_reg_931__2_ ( .D(n13171), .CP(wclk), .Q(ram[8930]) );
  DFF ram_reg_931__1_ ( .D(n13170), .CP(wclk), .Q(ram[8929]) );
  DFF ram_reg_931__0_ ( .D(n13169), .CP(wclk), .Q(ram[8928]) );
  DFF ram_reg_935__7_ ( .D(n13144), .CP(wclk), .Q(ram[8903]) );
  DFF ram_reg_935__6_ ( .D(n13143), .CP(wclk), .Q(ram[8902]) );
  DFF ram_reg_935__5_ ( .D(n13142), .CP(wclk), .Q(ram[8901]) );
  DFF ram_reg_935__4_ ( .D(n13141), .CP(wclk), .Q(ram[8900]) );
  DFF ram_reg_935__3_ ( .D(n13140), .CP(wclk), .Q(ram[8899]) );
  DFF ram_reg_935__2_ ( .D(n13139), .CP(wclk), .Q(ram[8898]) );
  DFF ram_reg_935__1_ ( .D(n13138), .CP(wclk), .Q(ram[8897]) );
  DFF ram_reg_935__0_ ( .D(n13137), .CP(wclk), .Q(ram[8896]) );
  DFF ram_reg_939__7_ ( .D(n13112), .CP(wclk), .Q(ram[8871]) );
  DFF ram_reg_939__6_ ( .D(n13111), .CP(wclk), .Q(ram[8870]) );
  DFF ram_reg_939__5_ ( .D(n13110), .CP(wclk), .Q(ram[8869]) );
  DFF ram_reg_939__4_ ( .D(n13109), .CP(wclk), .Q(ram[8868]) );
  DFF ram_reg_939__3_ ( .D(n13108), .CP(wclk), .Q(ram[8867]) );
  DFF ram_reg_939__2_ ( .D(n13107), .CP(wclk), .Q(ram[8866]) );
  DFF ram_reg_939__1_ ( .D(n13106), .CP(wclk), .Q(ram[8865]) );
  DFF ram_reg_939__0_ ( .D(n13105), .CP(wclk), .Q(ram[8864]) );
  DFF ram_reg_943__7_ ( .D(n13080), .CP(wclk), .Q(ram[8839]) );
  DFF ram_reg_943__6_ ( .D(n13079), .CP(wclk), .Q(ram[8838]) );
  DFF ram_reg_943__5_ ( .D(n13078), .CP(wclk), .Q(ram[8837]) );
  DFF ram_reg_943__4_ ( .D(n13077), .CP(wclk), .Q(ram[8836]) );
  DFF ram_reg_943__3_ ( .D(n13076), .CP(wclk), .Q(ram[8835]) );
  DFF ram_reg_943__2_ ( .D(n13075), .CP(wclk), .Q(ram[8834]) );
  DFF ram_reg_943__1_ ( .D(n13074), .CP(wclk), .Q(ram[8833]) );
  DFF ram_reg_943__0_ ( .D(n13073), .CP(wclk), .Q(ram[8832]) );
  DFF ram_reg_947__7_ ( .D(n13048), .CP(wclk), .Q(ram[8807]) );
  DFF ram_reg_947__6_ ( .D(n13047), .CP(wclk), .Q(ram[8806]) );
  DFF ram_reg_947__5_ ( .D(n13046), .CP(wclk), .Q(ram[8805]) );
  DFF ram_reg_947__4_ ( .D(n13045), .CP(wclk), .Q(ram[8804]) );
  DFF ram_reg_947__3_ ( .D(n13044), .CP(wclk), .Q(ram[8803]) );
  DFF ram_reg_947__2_ ( .D(n13043), .CP(wclk), .Q(ram[8802]) );
  DFF ram_reg_947__1_ ( .D(n13042), .CP(wclk), .Q(ram[8801]) );
  DFF ram_reg_947__0_ ( .D(n13041), .CP(wclk), .Q(ram[8800]) );
  DFF ram_reg_951__7_ ( .D(n13016), .CP(wclk), .Q(ram[8775]) );
  DFF ram_reg_951__6_ ( .D(n13015), .CP(wclk), .Q(ram[8774]) );
  DFF ram_reg_951__5_ ( .D(n13014), .CP(wclk), .Q(ram[8773]) );
  DFF ram_reg_951__4_ ( .D(n13013), .CP(wclk), .Q(ram[8772]) );
  DFF ram_reg_951__3_ ( .D(n13012), .CP(wclk), .Q(ram[8771]) );
  DFF ram_reg_951__2_ ( .D(n13011), .CP(wclk), .Q(ram[8770]) );
  DFF ram_reg_951__1_ ( .D(n13010), .CP(wclk), .Q(ram[8769]) );
  DFF ram_reg_951__0_ ( .D(n13009), .CP(wclk), .Q(ram[8768]) );
  DFF ram_reg_955__7_ ( .D(n12984), .CP(wclk), .Q(ram[8743]) );
  DFF ram_reg_955__6_ ( .D(n12983), .CP(wclk), .Q(ram[8742]) );
  DFF ram_reg_955__5_ ( .D(n12982), .CP(wclk), .Q(ram[8741]) );
  DFF ram_reg_955__4_ ( .D(n12981), .CP(wclk), .Q(ram[8740]) );
  DFF ram_reg_955__3_ ( .D(n12980), .CP(wclk), .Q(ram[8739]) );
  DFF ram_reg_955__2_ ( .D(n12979), .CP(wclk), .Q(ram[8738]) );
  DFF ram_reg_955__1_ ( .D(n12978), .CP(wclk), .Q(ram[8737]) );
  DFF ram_reg_955__0_ ( .D(n12977), .CP(wclk), .Q(ram[8736]) );
  DFF ram_reg_959__7_ ( .D(n12952), .CP(wclk), .Q(ram[8711]) );
  DFF ram_reg_959__6_ ( .D(n12951), .CP(wclk), .Q(ram[8710]) );
  DFF ram_reg_959__5_ ( .D(n12950), .CP(wclk), .Q(ram[8709]) );
  DFF ram_reg_959__4_ ( .D(n12949), .CP(wclk), .Q(ram[8708]) );
  DFF ram_reg_959__3_ ( .D(n12948), .CP(wclk), .Q(ram[8707]) );
  DFF ram_reg_959__2_ ( .D(n12947), .CP(wclk), .Q(ram[8706]) );
  DFF ram_reg_959__1_ ( .D(n12946), .CP(wclk), .Q(ram[8705]) );
  DFF ram_reg_959__0_ ( .D(n12945), .CP(wclk), .Q(ram[8704]) );
  DFF ram_reg_963__7_ ( .D(n12920), .CP(wclk), .Q(ram[8679]) );
  DFF ram_reg_963__6_ ( .D(n12919), .CP(wclk), .Q(ram[8678]) );
  DFF ram_reg_963__5_ ( .D(n12918), .CP(wclk), .Q(ram[8677]) );
  DFF ram_reg_963__4_ ( .D(n12917), .CP(wclk), .Q(ram[8676]) );
  DFF ram_reg_963__3_ ( .D(n12916), .CP(wclk), .Q(ram[8675]) );
  DFF ram_reg_963__2_ ( .D(n12915), .CP(wclk), .Q(ram[8674]) );
  DFF ram_reg_963__1_ ( .D(n12914), .CP(wclk), .Q(ram[8673]) );
  DFF ram_reg_963__0_ ( .D(n12913), .CP(wclk), .Q(ram[8672]) );
  DFF ram_reg_971__7_ ( .D(n12856), .CP(wclk), .Q(ram[8615]) );
  DFF ram_reg_971__6_ ( .D(n12855), .CP(wclk), .Q(ram[8614]) );
  DFF ram_reg_971__5_ ( .D(n12854), .CP(wclk), .Q(ram[8613]) );
  DFF ram_reg_971__4_ ( .D(n12853), .CP(wclk), .Q(ram[8612]) );
  DFF ram_reg_971__3_ ( .D(n12852), .CP(wclk), .Q(ram[8611]) );
  DFF ram_reg_971__2_ ( .D(n12851), .CP(wclk), .Q(ram[8610]) );
  DFF ram_reg_971__1_ ( .D(n12850), .CP(wclk), .Q(ram[8609]) );
  DFF ram_reg_971__0_ ( .D(n12849), .CP(wclk), .Q(ram[8608]) );
  DFF ram_reg_975__7_ ( .D(n12824), .CP(wclk), .Q(ram[8583]) );
  DFF ram_reg_975__6_ ( .D(n12823), .CP(wclk), .Q(ram[8582]) );
  DFF ram_reg_975__5_ ( .D(n12822), .CP(wclk), .Q(ram[8581]) );
  DFF ram_reg_975__4_ ( .D(n12821), .CP(wclk), .Q(ram[8580]) );
  DFF ram_reg_975__3_ ( .D(n12820), .CP(wclk), .Q(ram[8579]) );
  DFF ram_reg_975__2_ ( .D(n12819), .CP(wclk), .Q(ram[8578]) );
  DFF ram_reg_975__1_ ( .D(n12818), .CP(wclk), .Q(ram[8577]) );
  DFF ram_reg_975__0_ ( .D(n12817), .CP(wclk), .Q(ram[8576]) );
  DFF ram_reg_979__7_ ( .D(n12792), .CP(wclk), .Q(ram[8551]) );
  DFF ram_reg_979__6_ ( .D(n12791), .CP(wclk), .Q(ram[8550]) );
  DFF ram_reg_979__5_ ( .D(n12790), .CP(wclk), .Q(ram[8549]) );
  DFF ram_reg_979__4_ ( .D(n12789), .CP(wclk), .Q(ram[8548]) );
  DFF ram_reg_979__3_ ( .D(n12788), .CP(wclk), .Q(ram[8547]) );
  DFF ram_reg_979__2_ ( .D(n12787), .CP(wclk), .Q(ram[8546]) );
  DFF ram_reg_979__1_ ( .D(n12786), .CP(wclk), .Q(ram[8545]) );
  DFF ram_reg_979__0_ ( .D(n12785), .CP(wclk), .Q(ram[8544]) );
  DFF ram_reg_987__7_ ( .D(n12728), .CP(wclk), .Q(ram[8487]) );
  DFF ram_reg_987__6_ ( .D(n12727), .CP(wclk), .Q(ram[8486]) );
  DFF ram_reg_987__5_ ( .D(n12726), .CP(wclk), .Q(ram[8485]) );
  DFF ram_reg_987__4_ ( .D(n12725), .CP(wclk), .Q(ram[8484]) );
  DFF ram_reg_987__3_ ( .D(n12724), .CP(wclk), .Q(ram[8483]) );
  DFF ram_reg_987__2_ ( .D(n12723), .CP(wclk), .Q(ram[8482]) );
  DFF ram_reg_987__1_ ( .D(n12722), .CP(wclk), .Q(ram[8481]) );
  DFF ram_reg_987__0_ ( .D(n12721), .CP(wclk), .Q(ram[8480]) );
  DFF ram_reg_991__7_ ( .D(n12696), .CP(wclk), .Q(ram[8455]) );
  DFF ram_reg_991__6_ ( .D(n12695), .CP(wclk), .Q(ram[8454]) );
  DFF ram_reg_991__5_ ( .D(n12694), .CP(wclk), .Q(ram[8453]) );
  DFF ram_reg_991__4_ ( .D(n12693), .CP(wclk), .Q(ram[8452]) );
  DFF ram_reg_991__3_ ( .D(n12692), .CP(wclk), .Q(ram[8451]) );
  DFF ram_reg_991__2_ ( .D(n12691), .CP(wclk), .Q(ram[8450]) );
  DFF ram_reg_991__1_ ( .D(n12690), .CP(wclk), .Q(ram[8449]) );
  DFF ram_reg_991__0_ ( .D(n12689), .CP(wclk), .Q(ram[8448]) );
  DFF ram_reg_995__7_ ( .D(n12664), .CP(wclk), .Q(ram[8423]) );
  DFF ram_reg_995__6_ ( .D(n12663), .CP(wclk), .Q(ram[8422]) );
  DFF ram_reg_995__5_ ( .D(n12662), .CP(wclk), .Q(ram[8421]) );
  DFF ram_reg_995__4_ ( .D(n12661), .CP(wclk), .Q(ram[8420]) );
  DFF ram_reg_995__3_ ( .D(n12660), .CP(wclk), .Q(ram[8419]) );
  DFF ram_reg_995__2_ ( .D(n12659), .CP(wclk), .Q(ram[8418]) );
  DFF ram_reg_995__1_ ( .D(n12658), .CP(wclk), .Q(ram[8417]) );
  DFF ram_reg_995__0_ ( .D(n12657), .CP(wclk), .Q(ram[8416]) );
  DFF ram_reg_999__7_ ( .D(n12632), .CP(wclk), .Q(ram[8391]) );
  DFF ram_reg_999__6_ ( .D(n12631), .CP(wclk), .Q(ram[8390]) );
  DFF ram_reg_999__5_ ( .D(n12630), .CP(wclk), .Q(ram[8389]) );
  DFF ram_reg_999__4_ ( .D(n12629), .CP(wclk), .Q(ram[8388]) );
  DFF ram_reg_999__3_ ( .D(n12628), .CP(wclk), .Q(ram[8387]) );
  DFF ram_reg_999__2_ ( .D(n12627), .CP(wclk), .Q(ram[8386]) );
  DFF ram_reg_999__1_ ( .D(n12626), .CP(wclk), .Q(ram[8385]) );
  DFF ram_reg_999__0_ ( .D(n12625), .CP(wclk), .Q(ram[8384]) );
  DFF ram_reg_1003__7_ ( .D(n12600), .CP(wclk), .Q(ram[8359]) );
  DFF ram_reg_1003__6_ ( .D(n12599), .CP(wclk), .Q(ram[8358]) );
  DFF ram_reg_1003__5_ ( .D(n12598), .CP(wclk), .Q(ram[8357]) );
  DFF ram_reg_1003__4_ ( .D(n12597), .CP(wclk), .Q(ram[8356]) );
  DFF ram_reg_1003__3_ ( .D(n12596), .CP(wclk), .Q(ram[8355]) );
  DFF ram_reg_1003__2_ ( .D(n12595), .CP(wclk), .Q(ram[8354]) );
  DFF ram_reg_1003__1_ ( .D(n12594), .CP(wclk), .Q(ram[8353]) );
  DFF ram_reg_1003__0_ ( .D(n12593), .CP(wclk), .Q(ram[8352]) );
  DFF ram_reg_1007__7_ ( .D(n12568), .CP(wclk), .Q(ram[8327]) );
  DFF ram_reg_1007__6_ ( .D(n12567), .CP(wclk), .Q(ram[8326]) );
  DFF ram_reg_1007__5_ ( .D(n12566), .CP(wclk), .Q(ram[8325]) );
  DFF ram_reg_1007__4_ ( .D(n12565), .CP(wclk), .Q(ram[8324]) );
  DFF ram_reg_1007__3_ ( .D(n12564), .CP(wclk), .Q(ram[8323]) );
  DFF ram_reg_1007__2_ ( .D(n12563), .CP(wclk), .Q(ram[8322]) );
  DFF ram_reg_1007__1_ ( .D(n12562), .CP(wclk), .Q(ram[8321]) );
  DFF ram_reg_1007__0_ ( .D(n12561), .CP(wclk), .Q(ram[8320]) );
  DFF ram_reg_1011__7_ ( .D(n12536), .CP(wclk), .Q(ram[8295]) );
  DFF ram_reg_1011__6_ ( .D(n12535), .CP(wclk), .Q(ram[8294]) );
  DFF ram_reg_1011__5_ ( .D(n12534), .CP(wclk), .Q(ram[8293]) );
  DFF ram_reg_1011__4_ ( .D(n12533), .CP(wclk), .Q(ram[8292]) );
  DFF ram_reg_1011__3_ ( .D(n12532), .CP(wclk), .Q(ram[8291]) );
  DFF ram_reg_1011__2_ ( .D(n12531), .CP(wclk), .Q(ram[8290]) );
  DFF ram_reg_1011__1_ ( .D(n12530), .CP(wclk), .Q(ram[8289]) );
  DFF ram_reg_1011__0_ ( .D(n12529), .CP(wclk), .Q(ram[8288]) );
  DFF ram_reg_1015__7_ ( .D(n12504), .CP(wclk), .Q(ram[8263]) );
  DFF ram_reg_1015__6_ ( .D(n12503), .CP(wclk), .Q(ram[8262]) );
  DFF ram_reg_1015__5_ ( .D(n12502), .CP(wclk), .Q(ram[8261]) );
  DFF ram_reg_1015__4_ ( .D(n12501), .CP(wclk), .Q(ram[8260]) );
  DFF ram_reg_1015__3_ ( .D(n12500), .CP(wclk), .Q(ram[8259]) );
  DFF ram_reg_1015__2_ ( .D(n12499), .CP(wclk), .Q(ram[8258]) );
  DFF ram_reg_1015__1_ ( .D(n12498), .CP(wclk), .Q(ram[8257]) );
  DFF ram_reg_1015__0_ ( .D(n12497), .CP(wclk), .Q(ram[8256]) );
  DFF ram_reg_1019__7_ ( .D(n12472), .CP(wclk), .Q(ram[8231]) );
  DFF ram_reg_1019__6_ ( .D(n12471), .CP(wclk), .Q(ram[8230]) );
  DFF ram_reg_1019__5_ ( .D(n12470), .CP(wclk), .Q(ram[8229]) );
  DFF ram_reg_1019__4_ ( .D(n12469), .CP(wclk), .Q(ram[8228]) );
  DFF ram_reg_1019__3_ ( .D(n12468), .CP(wclk), .Q(ram[8227]) );
  DFF ram_reg_1019__2_ ( .D(n12467), .CP(wclk), .Q(ram[8226]) );
  DFF ram_reg_1019__1_ ( .D(n12466), .CP(wclk), .Q(ram[8225]) );
  DFF ram_reg_1019__0_ ( .D(n12465), .CP(wclk), .Q(ram[8224]) );
  DFF ram_reg_1023__7_ ( .D(n12440), .CP(wclk), .Q(ram[8199]) );
  DFF ram_reg_1023__6_ ( .D(n12439), .CP(wclk), .Q(ram[8198]) );
  DFF ram_reg_1023__5_ ( .D(n12438), .CP(wclk), .Q(ram[8197]) );
  DFF ram_reg_1023__4_ ( .D(n12437), .CP(wclk), .Q(ram[8196]) );
  DFF ram_reg_1023__3_ ( .D(n12436), .CP(wclk), .Q(ram[8195]) );
  DFF ram_reg_1023__2_ ( .D(n12435), .CP(wclk), .Q(ram[8194]) );
  DFF ram_reg_1023__1_ ( .D(n12434), .CP(wclk), .Q(ram[8193]) );
  DFF ram_reg_1023__0_ ( .D(n12433), .CP(wclk), .Q(ram[8192]) );
  DFF ram_reg_1035__7_ ( .D(n12344), .CP(wclk), .Q(ram[8103]) );
  DFF ram_reg_1035__6_ ( .D(n12343), .CP(wclk), .Q(ram[8102]) );
  DFF ram_reg_1035__5_ ( .D(n12342), .CP(wclk), .Q(ram[8101]) );
  DFF ram_reg_1035__4_ ( .D(n12341), .CP(wclk), .Q(ram[8100]) );
  DFF ram_reg_1035__3_ ( .D(n12340), .CP(wclk), .Q(ram[8099]) );
  DFF ram_reg_1035__2_ ( .D(n12339), .CP(wclk), .Q(ram[8098]) );
  DFF ram_reg_1035__1_ ( .D(n12338), .CP(wclk), .Q(ram[8097]) );
  DFF ram_reg_1035__0_ ( .D(n12337), .CP(wclk), .Q(ram[8096]) );
  DFF ram_reg_1039__7_ ( .D(n12312), .CP(wclk), .Q(ram[8071]) );
  DFF ram_reg_1039__6_ ( .D(n12311), .CP(wclk), .Q(ram[8070]) );
  DFF ram_reg_1039__5_ ( .D(n12310), .CP(wclk), .Q(ram[8069]) );
  DFF ram_reg_1039__4_ ( .D(n12309), .CP(wclk), .Q(ram[8068]) );
  DFF ram_reg_1039__3_ ( .D(n12308), .CP(wclk), .Q(ram[8067]) );
  DFF ram_reg_1039__2_ ( .D(n12307), .CP(wclk), .Q(ram[8066]) );
  DFF ram_reg_1039__1_ ( .D(n12306), .CP(wclk), .Q(ram[8065]) );
  DFF ram_reg_1039__0_ ( .D(n12305), .CP(wclk), .Q(ram[8064]) );
  DFF ram_reg_1051__7_ ( .D(n12216), .CP(wclk), .Q(ram[7975]) );
  DFF ram_reg_1051__6_ ( .D(n12215), .CP(wclk), .Q(ram[7974]) );
  DFF ram_reg_1051__5_ ( .D(n12214), .CP(wclk), .Q(ram[7973]) );
  DFF ram_reg_1051__4_ ( .D(n12213), .CP(wclk), .Q(ram[7972]) );
  DFF ram_reg_1051__3_ ( .D(n12212), .CP(wclk), .Q(ram[7971]) );
  DFF ram_reg_1051__2_ ( .D(n12211), .CP(wclk), .Q(ram[7970]) );
  DFF ram_reg_1051__1_ ( .D(n12210), .CP(wclk), .Q(ram[7969]) );
  DFF ram_reg_1051__0_ ( .D(n12209), .CP(wclk), .Q(ram[7968]) );
  DFF ram_reg_1059__7_ ( .D(n12152), .CP(wclk), .Q(ram[7911]) );
  DFF ram_reg_1059__6_ ( .D(n12151), .CP(wclk), .Q(ram[7910]) );
  DFF ram_reg_1059__5_ ( .D(n12150), .CP(wclk), .Q(ram[7909]) );
  DFF ram_reg_1059__4_ ( .D(n12149), .CP(wclk), .Q(ram[7908]) );
  DFF ram_reg_1059__3_ ( .D(n12148), .CP(wclk), .Q(ram[7907]) );
  DFF ram_reg_1059__2_ ( .D(n12147), .CP(wclk), .Q(ram[7906]) );
  DFF ram_reg_1059__1_ ( .D(n12146), .CP(wclk), .Q(ram[7905]) );
  DFF ram_reg_1059__0_ ( .D(n12145), .CP(wclk), .Q(ram[7904]) );
  DFF ram_reg_1067__7_ ( .D(n12088), .CP(wclk), .Q(ram[7847]) );
  DFF ram_reg_1067__6_ ( .D(n12087), .CP(wclk), .Q(ram[7846]) );
  DFF ram_reg_1067__5_ ( .D(n12086), .CP(wclk), .Q(ram[7845]) );
  DFF ram_reg_1067__4_ ( .D(n12085), .CP(wclk), .Q(ram[7844]) );
  DFF ram_reg_1067__3_ ( .D(n12084), .CP(wclk), .Q(ram[7843]) );
  DFF ram_reg_1067__2_ ( .D(n12083), .CP(wclk), .Q(ram[7842]) );
  DFF ram_reg_1067__1_ ( .D(n12082), .CP(wclk), .Q(ram[7841]) );
  DFF ram_reg_1067__0_ ( .D(n12081), .CP(wclk), .Q(ram[7840]) );
  DFF ram_reg_1071__7_ ( .D(n12056), .CP(wclk), .Q(ram[7815]) );
  DFF ram_reg_1071__6_ ( .D(n12055), .CP(wclk), .Q(ram[7814]) );
  DFF ram_reg_1071__5_ ( .D(n12054), .CP(wclk), .Q(ram[7813]) );
  DFF ram_reg_1071__4_ ( .D(n12053), .CP(wclk), .Q(ram[7812]) );
  DFF ram_reg_1071__3_ ( .D(n12052), .CP(wclk), .Q(ram[7811]) );
  DFF ram_reg_1071__2_ ( .D(n12051), .CP(wclk), .Q(ram[7810]) );
  DFF ram_reg_1071__1_ ( .D(n12050), .CP(wclk), .Q(ram[7809]) );
  DFF ram_reg_1071__0_ ( .D(n12049), .CP(wclk), .Q(ram[7808]) );
  DFF ram_reg_1075__7_ ( .D(n12024), .CP(wclk), .Q(ram[7783]) );
  DFF ram_reg_1075__6_ ( .D(n12023), .CP(wclk), .Q(ram[7782]) );
  DFF ram_reg_1075__5_ ( .D(n12022), .CP(wclk), .Q(ram[7781]) );
  DFF ram_reg_1075__4_ ( .D(n12021), .CP(wclk), .Q(ram[7780]) );
  DFF ram_reg_1075__3_ ( .D(n12020), .CP(wclk), .Q(ram[7779]) );
  DFF ram_reg_1075__2_ ( .D(n12019), .CP(wclk), .Q(ram[7778]) );
  DFF ram_reg_1075__1_ ( .D(n12018), .CP(wclk), .Q(ram[7777]) );
  DFF ram_reg_1075__0_ ( .D(n12017), .CP(wclk), .Q(ram[7776]) );
  DFF ram_reg_1083__7_ ( .D(n11960), .CP(wclk), .Q(ram[7719]) );
  DFF ram_reg_1083__6_ ( .D(n11959), .CP(wclk), .Q(ram[7718]) );
  DFF ram_reg_1083__5_ ( .D(n11958), .CP(wclk), .Q(ram[7717]) );
  DFF ram_reg_1083__4_ ( .D(n11957), .CP(wclk), .Q(ram[7716]) );
  DFF ram_reg_1083__3_ ( .D(n11956), .CP(wclk), .Q(ram[7715]) );
  DFF ram_reg_1083__2_ ( .D(n11955), .CP(wclk), .Q(ram[7714]) );
  DFF ram_reg_1083__1_ ( .D(n11954), .CP(wclk), .Q(ram[7713]) );
  DFF ram_reg_1083__0_ ( .D(n11953), .CP(wclk), .Q(ram[7712]) );
  DFF ram_reg_1087__7_ ( .D(n11928), .CP(wclk), .Q(ram[7687]) );
  DFF ram_reg_1087__6_ ( .D(n11927), .CP(wclk), .Q(ram[7686]) );
  DFF ram_reg_1087__5_ ( .D(n11926), .CP(wclk), .Q(ram[7685]) );
  DFF ram_reg_1087__4_ ( .D(n11925), .CP(wclk), .Q(ram[7684]) );
  DFF ram_reg_1087__3_ ( .D(n11924), .CP(wclk), .Q(ram[7683]) );
  DFF ram_reg_1087__2_ ( .D(n11923), .CP(wclk), .Q(ram[7682]) );
  DFF ram_reg_1087__1_ ( .D(n11922), .CP(wclk), .Q(ram[7681]) );
  DFF ram_reg_1087__0_ ( .D(n11921), .CP(wclk), .Q(ram[7680]) );
  DFF ram_reg_1131__7_ ( .D(n11576), .CP(wclk), .Q(ram[7335]) );
  DFF ram_reg_1131__6_ ( .D(n11575), .CP(wclk), .Q(ram[7334]) );
  DFF ram_reg_1131__5_ ( .D(n11574), .CP(wclk), .Q(ram[7333]) );
  DFF ram_reg_1131__4_ ( .D(n11573), .CP(wclk), .Q(ram[7332]) );
  DFF ram_reg_1131__3_ ( .D(n11572), .CP(wclk), .Q(ram[7331]) );
  DFF ram_reg_1131__2_ ( .D(n11571), .CP(wclk), .Q(ram[7330]) );
  DFF ram_reg_1131__1_ ( .D(n11570), .CP(wclk), .Q(ram[7329]) );
  DFF ram_reg_1131__0_ ( .D(n11569), .CP(wclk), .Q(ram[7328]) );
  DFF ram_reg_1147__7_ ( .D(n11448), .CP(wclk), .Q(ram[7207]) );
  DFF ram_reg_1147__6_ ( .D(n11447), .CP(wclk), .Q(ram[7206]) );
  DFF ram_reg_1147__5_ ( .D(n11446), .CP(wclk), .Q(ram[7205]) );
  DFF ram_reg_1147__4_ ( .D(n11445), .CP(wclk), .Q(ram[7204]) );
  DFF ram_reg_1147__3_ ( .D(n11444), .CP(wclk), .Q(ram[7203]) );
  DFF ram_reg_1147__2_ ( .D(n11443), .CP(wclk), .Q(ram[7202]) );
  DFF ram_reg_1147__1_ ( .D(n11442), .CP(wclk), .Q(ram[7201]) );
  DFF ram_reg_1147__0_ ( .D(n11441), .CP(wclk), .Q(ram[7200]) );
  DFF ram_reg_1151__7_ ( .D(n11416), .CP(wclk), .Q(ram[7175]) );
  DFF ram_reg_1151__6_ ( .D(n11415), .CP(wclk), .Q(ram[7174]) );
  DFF ram_reg_1151__5_ ( .D(n11414), .CP(wclk), .Q(ram[7173]) );
  DFF ram_reg_1151__4_ ( .D(n11413), .CP(wclk), .Q(ram[7172]) );
  DFF ram_reg_1151__3_ ( .D(n11412), .CP(wclk), .Q(ram[7171]) );
  DFF ram_reg_1151__2_ ( .D(n11411), .CP(wclk), .Q(ram[7170]) );
  DFF ram_reg_1151__1_ ( .D(n11410), .CP(wclk), .Q(ram[7169]) );
  DFF ram_reg_1151__0_ ( .D(n11409), .CP(wclk), .Q(ram[7168]) );
  DFF ram_reg_1155__7_ ( .D(n11384), .CP(wclk), .Q(ram[7143]) );
  DFF ram_reg_1155__6_ ( .D(n11383), .CP(wclk), .Q(ram[7142]) );
  DFF ram_reg_1155__5_ ( .D(n11382), .CP(wclk), .Q(ram[7141]) );
  DFF ram_reg_1155__4_ ( .D(n11381), .CP(wclk), .Q(ram[7140]) );
  DFF ram_reg_1155__3_ ( .D(n11380), .CP(wclk), .Q(ram[7139]) );
  DFF ram_reg_1155__2_ ( .D(n11379), .CP(wclk), .Q(ram[7138]) );
  DFF ram_reg_1155__1_ ( .D(n11378), .CP(wclk), .Q(ram[7137]) );
  DFF ram_reg_1155__0_ ( .D(n11377), .CP(wclk), .Q(ram[7136]) );
  DFF ram_reg_1163__7_ ( .D(n11320), .CP(wclk), .Q(ram[7079]) );
  DFF ram_reg_1163__6_ ( .D(n11319), .CP(wclk), .Q(ram[7078]) );
  DFF ram_reg_1163__5_ ( .D(n11318), .CP(wclk), .Q(ram[7077]) );
  DFF ram_reg_1163__4_ ( .D(n11317), .CP(wclk), .Q(ram[7076]) );
  DFF ram_reg_1163__3_ ( .D(n11316), .CP(wclk), .Q(ram[7075]) );
  DFF ram_reg_1163__2_ ( .D(n11315), .CP(wclk), .Q(ram[7074]) );
  DFF ram_reg_1163__1_ ( .D(n11314), .CP(wclk), .Q(ram[7073]) );
  DFF ram_reg_1163__0_ ( .D(n11313), .CP(wclk), .Q(ram[7072]) );
  DFF ram_reg_1167__7_ ( .D(n11288), .CP(wclk), .Q(ram[7047]) );
  DFF ram_reg_1167__6_ ( .D(n11287), .CP(wclk), .Q(ram[7046]) );
  DFF ram_reg_1167__5_ ( .D(n11286), .CP(wclk), .Q(ram[7045]) );
  DFF ram_reg_1167__4_ ( .D(n11285), .CP(wclk), .Q(ram[7044]) );
  DFF ram_reg_1167__3_ ( .D(n11284), .CP(wclk), .Q(ram[7043]) );
  DFF ram_reg_1167__2_ ( .D(n11283), .CP(wclk), .Q(ram[7042]) );
  DFF ram_reg_1167__1_ ( .D(n11282), .CP(wclk), .Q(ram[7041]) );
  DFF ram_reg_1167__0_ ( .D(n11281), .CP(wclk), .Q(ram[7040]) );
  DFF ram_reg_1171__7_ ( .D(n11256), .CP(wclk), .Q(ram[7015]) );
  DFF ram_reg_1171__6_ ( .D(n11255), .CP(wclk), .Q(ram[7014]) );
  DFF ram_reg_1171__5_ ( .D(n11254), .CP(wclk), .Q(ram[7013]) );
  DFF ram_reg_1171__4_ ( .D(n11253), .CP(wclk), .Q(ram[7012]) );
  DFF ram_reg_1171__3_ ( .D(n11252), .CP(wclk), .Q(ram[7011]) );
  DFF ram_reg_1171__2_ ( .D(n11251), .CP(wclk), .Q(ram[7010]) );
  DFF ram_reg_1171__1_ ( .D(n11250), .CP(wclk), .Q(ram[7009]) );
  DFF ram_reg_1171__0_ ( .D(n11249), .CP(wclk), .Q(ram[7008]) );
  DFF ram_reg_1179__7_ ( .D(n11192), .CP(wclk), .Q(ram[6951]) );
  DFF ram_reg_1179__6_ ( .D(n11191), .CP(wclk), .Q(ram[6950]) );
  DFF ram_reg_1179__5_ ( .D(n11190), .CP(wclk), .Q(ram[6949]) );
  DFF ram_reg_1179__4_ ( .D(n11189), .CP(wclk), .Q(ram[6948]) );
  DFF ram_reg_1179__3_ ( .D(n11188), .CP(wclk), .Q(ram[6947]) );
  DFF ram_reg_1179__2_ ( .D(n11187), .CP(wclk), .Q(ram[6946]) );
  DFF ram_reg_1179__1_ ( .D(n11186), .CP(wclk), .Q(ram[6945]) );
  DFF ram_reg_1179__0_ ( .D(n11185), .CP(wclk), .Q(ram[6944]) );
  DFF ram_reg_1183__7_ ( .D(n11160), .CP(wclk), .Q(ram[6919]) );
  DFF ram_reg_1183__6_ ( .D(n11159), .CP(wclk), .Q(ram[6918]) );
  DFF ram_reg_1183__5_ ( .D(n11158), .CP(wclk), .Q(ram[6917]) );
  DFF ram_reg_1183__4_ ( .D(n11157), .CP(wclk), .Q(ram[6916]) );
  DFF ram_reg_1183__3_ ( .D(n11156), .CP(wclk), .Q(ram[6915]) );
  DFF ram_reg_1183__2_ ( .D(n11155), .CP(wclk), .Q(ram[6914]) );
  DFF ram_reg_1183__1_ ( .D(n11154), .CP(wclk), .Q(ram[6913]) );
  DFF ram_reg_1183__0_ ( .D(n11153), .CP(wclk), .Q(ram[6912]) );
  DFF ram_reg_1187__7_ ( .D(n11128), .CP(wclk), .Q(ram[6887]) );
  DFF ram_reg_1187__6_ ( .D(n11127), .CP(wclk), .Q(ram[6886]) );
  DFF ram_reg_1187__5_ ( .D(n11126), .CP(wclk), .Q(ram[6885]) );
  DFF ram_reg_1187__4_ ( .D(n11125), .CP(wclk), .Q(ram[6884]) );
  DFF ram_reg_1187__3_ ( .D(n11124), .CP(wclk), .Q(ram[6883]) );
  DFF ram_reg_1187__2_ ( .D(n11123), .CP(wclk), .Q(ram[6882]) );
  DFF ram_reg_1187__1_ ( .D(n11122), .CP(wclk), .Q(ram[6881]) );
  DFF ram_reg_1187__0_ ( .D(n11121), .CP(wclk), .Q(ram[6880]) );
  DFF ram_reg_1191__7_ ( .D(n11096), .CP(wclk), .Q(ram[6855]) );
  DFF ram_reg_1191__6_ ( .D(n11095), .CP(wclk), .Q(ram[6854]) );
  DFF ram_reg_1191__5_ ( .D(n11094), .CP(wclk), .Q(ram[6853]) );
  DFF ram_reg_1191__4_ ( .D(n11093), .CP(wclk), .Q(ram[6852]) );
  DFF ram_reg_1191__3_ ( .D(n11092), .CP(wclk), .Q(ram[6851]) );
  DFF ram_reg_1191__2_ ( .D(n11091), .CP(wclk), .Q(ram[6850]) );
  DFF ram_reg_1191__1_ ( .D(n11090), .CP(wclk), .Q(ram[6849]) );
  DFF ram_reg_1191__0_ ( .D(n11089), .CP(wclk), .Q(ram[6848]) );
  DFF ram_reg_1195__7_ ( .D(n11064), .CP(wclk), .Q(ram[6823]) );
  DFF ram_reg_1195__6_ ( .D(n11063), .CP(wclk), .Q(ram[6822]) );
  DFF ram_reg_1195__5_ ( .D(n11062), .CP(wclk), .Q(ram[6821]) );
  DFF ram_reg_1195__4_ ( .D(n11061), .CP(wclk), .Q(ram[6820]) );
  DFF ram_reg_1195__3_ ( .D(n11060), .CP(wclk), .Q(ram[6819]) );
  DFF ram_reg_1195__2_ ( .D(n11059), .CP(wclk), .Q(ram[6818]) );
  DFF ram_reg_1195__1_ ( .D(n11058), .CP(wclk), .Q(ram[6817]) );
  DFF ram_reg_1195__0_ ( .D(n11057), .CP(wclk), .Q(ram[6816]) );
  DFF ram_reg_1199__7_ ( .D(n11032), .CP(wclk), .Q(ram[6791]) );
  DFF ram_reg_1199__6_ ( .D(n11031), .CP(wclk), .Q(ram[6790]) );
  DFF ram_reg_1199__5_ ( .D(n11030), .CP(wclk), .Q(ram[6789]) );
  DFF ram_reg_1199__4_ ( .D(n11029), .CP(wclk), .Q(ram[6788]) );
  DFF ram_reg_1199__3_ ( .D(n11028), .CP(wclk), .Q(ram[6787]) );
  DFF ram_reg_1199__2_ ( .D(n11027), .CP(wclk), .Q(ram[6786]) );
  DFF ram_reg_1199__1_ ( .D(n11026), .CP(wclk), .Q(ram[6785]) );
  DFF ram_reg_1199__0_ ( .D(n11025), .CP(wclk), .Q(ram[6784]) );
  DFF ram_reg_1203__7_ ( .D(n11000), .CP(wclk), .Q(ram[6759]) );
  DFF ram_reg_1203__6_ ( .D(n10999), .CP(wclk), .Q(ram[6758]) );
  DFF ram_reg_1203__5_ ( .D(n10998), .CP(wclk), .Q(ram[6757]) );
  DFF ram_reg_1203__4_ ( .D(n10997), .CP(wclk), .Q(ram[6756]) );
  DFF ram_reg_1203__3_ ( .D(n10996), .CP(wclk), .Q(ram[6755]) );
  DFF ram_reg_1203__2_ ( .D(n10995), .CP(wclk), .Q(ram[6754]) );
  DFF ram_reg_1203__1_ ( .D(n10994), .CP(wclk), .Q(ram[6753]) );
  DFF ram_reg_1203__0_ ( .D(n10993), .CP(wclk), .Q(ram[6752]) );
  DFF ram_reg_1207__7_ ( .D(n10968), .CP(wclk), .Q(ram[6727]) );
  DFF ram_reg_1207__6_ ( .D(n10967), .CP(wclk), .Q(ram[6726]) );
  DFF ram_reg_1207__5_ ( .D(n10966), .CP(wclk), .Q(ram[6725]) );
  DFF ram_reg_1207__4_ ( .D(n10965), .CP(wclk), .Q(ram[6724]) );
  DFF ram_reg_1207__3_ ( .D(n10964), .CP(wclk), .Q(ram[6723]) );
  DFF ram_reg_1207__2_ ( .D(n10963), .CP(wclk), .Q(ram[6722]) );
  DFF ram_reg_1207__1_ ( .D(n10962), .CP(wclk), .Q(ram[6721]) );
  DFF ram_reg_1207__0_ ( .D(n10961), .CP(wclk), .Q(ram[6720]) );
  DFF ram_reg_1211__7_ ( .D(n10936), .CP(wclk), .Q(ram[6695]) );
  DFF ram_reg_1211__6_ ( .D(n10935), .CP(wclk), .Q(ram[6694]) );
  DFF ram_reg_1211__5_ ( .D(n10934), .CP(wclk), .Q(ram[6693]) );
  DFF ram_reg_1211__4_ ( .D(n10933), .CP(wclk), .Q(ram[6692]) );
  DFF ram_reg_1211__3_ ( .D(n10932), .CP(wclk), .Q(ram[6691]) );
  DFF ram_reg_1211__2_ ( .D(n10931), .CP(wclk), .Q(ram[6690]) );
  DFF ram_reg_1211__1_ ( .D(n10930), .CP(wclk), .Q(ram[6689]) );
  DFF ram_reg_1211__0_ ( .D(n10929), .CP(wclk), .Q(ram[6688]) );
  DFF ram_reg_1215__7_ ( .D(n10904), .CP(wclk), .Q(ram[6663]) );
  DFF ram_reg_1215__6_ ( .D(n10903), .CP(wclk), .Q(ram[6662]) );
  DFF ram_reg_1215__5_ ( .D(n10902), .CP(wclk), .Q(ram[6661]) );
  DFF ram_reg_1215__4_ ( .D(n10901), .CP(wclk), .Q(ram[6660]) );
  DFF ram_reg_1215__3_ ( .D(n10900), .CP(wclk), .Q(ram[6659]) );
  DFF ram_reg_1215__2_ ( .D(n10899), .CP(wclk), .Q(ram[6658]) );
  DFF ram_reg_1215__1_ ( .D(n10898), .CP(wclk), .Q(ram[6657]) );
  DFF ram_reg_1215__0_ ( .D(n10897), .CP(wclk), .Q(ram[6656]) );
  DFF ram_reg_1219__7_ ( .D(n10872), .CP(wclk), .Q(ram[6631]) );
  DFF ram_reg_1219__6_ ( .D(n10871), .CP(wclk), .Q(ram[6630]) );
  DFF ram_reg_1219__5_ ( .D(n10870), .CP(wclk), .Q(ram[6629]) );
  DFF ram_reg_1219__4_ ( .D(n10869), .CP(wclk), .Q(ram[6628]) );
  DFF ram_reg_1219__3_ ( .D(n10868), .CP(wclk), .Q(ram[6627]) );
  DFF ram_reg_1219__2_ ( .D(n10867), .CP(wclk), .Q(ram[6626]) );
  DFF ram_reg_1219__1_ ( .D(n10866), .CP(wclk), .Q(ram[6625]) );
  DFF ram_reg_1219__0_ ( .D(n10865), .CP(wclk), .Q(ram[6624]) );
  DFF ram_reg_1227__7_ ( .D(n10808), .CP(wclk), .Q(ram[6567]) );
  DFF ram_reg_1227__6_ ( .D(n10807), .CP(wclk), .Q(ram[6566]) );
  DFF ram_reg_1227__5_ ( .D(n10806), .CP(wclk), .Q(ram[6565]) );
  DFF ram_reg_1227__4_ ( .D(n10805), .CP(wclk), .Q(ram[6564]) );
  DFF ram_reg_1227__3_ ( .D(n10804), .CP(wclk), .Q(ram[6563]) );
  DFF ram_reg_1227__2_ ( .D(n10803), .CP(wclk), .Q(ram[6562]) );
  DFF ram_reg_1227__1_ ( .D(n10802), .CP(wclk), .Q(ram[6561]) );
  DFF ram_reg_1227__0_ ( .D(n10801), .CP(wclk), .Q(ram[6560]) );
  DFF ram_reg_1231__7_ ( .D(n10776), .CP(wclk), .Q(ram[6535]) );
  DFF ram_reg_1231__6_ ( .D(n10775), .CP(wclk), .Q(ram[6534]) );
  DFF ram_reg_1231__5_ ( .D(n10774), .CP(wclk), .Q(ram[6533]) );
  DFF ram_reg_1231__4_ ( .D(n10773), .CP(wclk), .Q(ram[6532]) );
  DFF ram_reg_1231__3_ ( .D(n10772), .CP(wclk), .Q(ram[6531]) );
  DFF ram_reg_1231__2_ ( .D(n10771), .CP(wclk), .Q(ram[6530]) );
  DFF ram_reg_1231__1_ ( .D(n10770), .CP(wclk), .Q(ram[6529]) );
  DFF ram_reg_1231__0_ ( .D(n10769), .CP(wclk), .Q(ram[6528]) );
  DFF ram_reg_1243__7_ ( .D(n10680), .CP(wclk), .Q(ram[6439]) );
  DFF ram_reg_1243__6_ ( .D(n10679), .CP(wclk), .Q(ram[6438]) );
  DFF ram_reg_1243__5_ ( .D(n10678), .CP(wclk), .Q(ram[6437]) );
  DFF ram_reg_1243__4_ ( .D(n10677), .CP(wclk), .Q(ram[6436]) );
  DFF ram_reg_1243__3_ ( .D(n10676), .CP(wclk), .Q(ram[6435]) );
  DFF ram_reg_1243__2_ ( .D(n10675), .CP(wclk), .Q(ram[6434]) );
  DFF ram_reg_1243__1_ ( .D(n10674), .CP(wclk), .Q(ram[6433]) );
  DFF ram_reg_1243__0_ ( .D(n10673), .CP(wclk), .Q(ram[6432]) );
  DFF ram_reg_1247__7_ ( .D(n10648), .CP(wclk), .Q(ram[6407]) );
  DFF ram_reg_1247__6_ ( .D(n10647), .CP(wclk), .Q(ram[6406]) );
  DFF ram_reg_1247__5_ ( .D(n10646), .CP(wclk), .Q(ram[6405]) );
  DFF ram_reg_1247__4_ ( .D(n10645), .CP(wclk), .Q(ram[6404]) );
  DFF ram_reg_1247__3_ ( .D(n10644), .CP(wclk), .Q(ram[6403]) );
  DFF ram_reg_1247__2_ ( .D(n10643), .CP(wclk), .Q(ram[6402]) );
  DFF ram_reg_1247__1_ ( .D(n10642), .CP(wclk), .Q(ram[6401]) );
  DFF ram_reg_1247__0_ ( .D(n10641), .CP(wclk), .Q(ram[6400]) );
  DFF ram_reg_1251__7_ ( .D(n10616), .CP(wclk), .Q(ram[6375]) );
  DFF ram_reg_1251__6_ ( .D(n10615), .CP(wclk), .Q(ram[6374]) );
  DFF ram_reg_1251__5_ ( .D(n10614), .CP(wclk), .Q(ram[6373]) );
  DFF ram_reg_1251__4_ ( .D(n10613), .CP(wclk), .Q(ram[6372]) );
  DFF ram_reg_1251__3_ ( .D(n10612), .CP(wclk), .Q(ram[6371]) );
  DFF ram_reg_1251__2_ ( .D(n10611), .CP(wclk), .Q(ram[6370]) );
  DFF ram_reg_1251__1_ ( .D(n10610), .CP(wclk), .Q(ram[6369]) );
  DFF ram_reg_1251__0_ ( .D(n10609), .CP(wclk), .Q(ram[6368]) );
  DFF ram_reg_1259__7_ ( .D(n10552), .CP(wclk), .Q(ram[6311]) );
  DFF ram_reg_1259__6_ ( .D(n10551), .CP(wclk), .Q(ram[6310]) );
  DFF ram_reg_1259__5_ ( .D(n10550), .CP(wclk), .Q(ram[6309]) );
  DFF ram_reg_1259__4_ ( .D(n10549), .CP(wclk), .Q(ram[6308]) );
  DFF ram_reg_1259__3_ ( .D(n10548), .CP(wclk), .Q(ram[6307]) );
  DFF ram_reg_1259__2_ ( .D(n10547), .CP(wclk), .Q(ram[6306]) );
  DFF ram_reg_1259__1_ ( .D(n10546), .CP(wclk), .Q(ram[6305]) );
  DFF ram_reg_1259__0_ ( .D(n10545), .CP(wclk), .Q(ram[6304]) );
  DFF ram_reg_1263__7_ ( .D(n10520), .CP(wclk), .Q(ram[6279]) );
  DFF ram_reg_1263__6_ ( .D(n10519), .CP(wclk), .Q(ram[6278]) );
  DFF ram_reg_1263__5_ ( .D(n10518), .CP(wclk), .Q(ram[6277]) );
  DFF ram_reg_1263__4_ ( .D(n10517), .CP(wclk), .Q(ram[6276]) );
  DFF ram_reg_1263__3_ ( .D(n10516), .CP(wclk), .Q(ram[6275]) );
  DFF ram_reg_1263__2_ ( .D(n10515), .CP(wclk), .Q(ram[6274]) );
  DFF ram_reg_1263__1_ ( .D(n10514), .CP(wclk), .Q(ram[6273]) );
  DFF ram_reg_1263__0_ ( .D(n10513), .CP(wclk), .Q(ram[6272]) );
  DFF ram_reg_1267__7_ ( .D(n10488), .CP(wclk), .Q(ram[6247]) );
  DFF ram_reg_1267__6_ ( .D(n10487), .CP(wclk), .Q(ram[6246]) );
  DFF ram_reg_1267__5_ ( .D(n10486), .CP(wclk), .Q(ram[6245]) );
  DFF ram_reg_1267__4_ ( .D(n10485), .CP(wclk), .Q(ram[6244]) );
  DFF ram_reg_1267__3_ ( .D(n10484), .CP(wclk), .Q(ram[6243]) );
  DFF ram_reg_1267__2_ ( .D(n10483), .CP(wclk), .Q(ram[6242]) );
  DFF ram_reg_1267__1_ ( .D(n10482), .CP(wclk), .Q(ram[6241]) );
  DFF ram_reg_1267__0_ ( .D(n10481), .CP(wclk), .Q(ram[6240]) );
  DFF ram_reg_1271__7_ ( .D(n10456), .CP(wclk), .Q(ram[6215]) );
  DFF ram_reg_1271__6_ ( .D(n10455), .CP(wclk), .Q(ram[6214]) );
  DFF ram_reg_1271__5_ ( .D(n10454), .CP(wclk), .Q(ram[6213]) );
  DFF ram_reg_1271__4_ ( .D(n10453), .CP(wclk), .Q(ram[6212]) );
  DFF ram_reg_1271__3_ ( .D(n10452), .CP(wclk), .Q(ram[6211]) );
  DFF ram_reg_1271__2_ ( .D(n10451), .CP(wclk), .Q(ram[6210]) );
  DFF ram_reg_1271__1_ ( .D(n10450), .CP(wclk), .Q(ram[6209]) );
  DFF ram_reg_1271__0_ ( .D(n10449), .CP(wclk), .Q(ram[6208]) );
  DFF ram_reg_1275__7_ ( .D(n10424), .CP(wclk), .Q(ram[6183]) );
  DFF ram_reg_1275__6_ ( .D(n10423), .CP(wclk), .Q(ram[6182]) );
  DFF ram_reg_1275__5_ ( .D(n10422), .CP(wclk), .Q(ram[6181]) );
  DFF ram_reg_1275__4_ ( .D(n10421), .CP(wclk), .Q(ram[6180]) );
  DFF ram_reg_1275__3_ ( .D(n10420), .CP(wclk), .Q(ram[6179]) );
  DFF ram_reg_1275__2_ ( .D(n10419), .CP(wclk), .Q(ram[6178]) );
  DFF ram_reg_1275__1_ ( .D(n10418), .CP(wclk), .Q(ram[6177]) );
  DFF ram_reg_1275__0_ ( .D(n10417), .CP(wclk), .Q(ram[6176]) );
  DFF ram_reg_1279__7_ ( .D(n10392), .CP(wclk), .Q(ram[6151]) );
  DFF ram_reg_1279__6_ ( .D(n10391), .CP(wclk), .Q(ram[6150]) );
  DFF ram_reg_1279__5_ ( .D(n10390), .CP(wclk), .Q(ram[6149]) );
  DFF ram_reg_1279__4_ ( .D(n10389), .CP(wclk), .Q(ram[6148]) );
  DFF ram_reg_1279__3_ ( .D(n10388), .CP(wclk), .Q(ram[6147]) );
  DFF ram_reg_1279__2_ ( .D(n10387), .CP(wclk), .Q(ram[6146]) );
  DFF ram_reg_1279__1_ ( .D(n10386), .CP(wclk), .Q(ram[6145]) );
  DFF ram_reg_1279__0_ ( .D(n10385), .CP(wclk), .Q(ram[6144]) );
  DFF ram_reg_1283__7_ ( .D(n10360), .CP(wclk), .Q(ram[6119]) );
  DFF ram_reg_1283__6_ ( .D(n10359), .CP(wclk), .Q(ram[6118]) );
  DFF ram_reg_1283__5_ ( .D(n10358), .CP(wclk), .Q(ram[6117]) );
  DFF ram_reg_1283__4_ ( .D(n10357), .CP(wclk), .Q(ram[6116]) );
  DFF ram_reg_1283__3_ ( .D(n10356), .CP(wclk), .Q(ram[6115]) );
  DFF ram_reg_1283__2_ ( .D(n10355), .CP(wclk), .Q(ram[6114]) );
  DFF ram_reg_1283__1_ ( .D(n10354), .CP(wclk), .Q(ram[6113]) );
  DFF ram_reg_1283__0_ ( .D(n10353), .CP(wclk), .Q(ram[6112]) );
  DFF ram_reg_1291__7_ ( .D(n10296), .CP(wclk), .Q(ram[6055]) );
  DFF ram_reg_1291__6_ ( .D(n10295), .CP(wclk), .Q(ram[6054]) );
  DFF ram_reg_1291__5_ ( .D(n10294), .CP(wclk), .Q(ram[6053]) );
  DFF ram_reg_1291__4_ ( .D(n10293), .CP(wclk), .Q(ram[6052]) );
  DFF ram_reg_1291__3_ ( .D(n10292), .CP(wclk), .Q(ram[6051]) );
  DFF ram_reg_1291__2_ ( .D(n10291), .CP(wclk), .Q(ram[6050]) );
  DFF ram_reg_1291__1_ ( .D(n10290), .CP(wclk), .Q(ram[6049]) );
  DFF ram_reg_1291__0_ ( .D(n10289), .CP(wclk), .Q(ram[6048]) );
  DFF ram_reg_1295__7_ ( .D(n10264), .CP(wclk), .Q(ram[6023]) );
  DFF ram_reg_1295__6_ ( .D(n10263), .CP(wclk), .Q(ram[6022]) );
  DFF ram_reg_1295__5_ ( .D(n10262), .CP(wclk), .Q(ram[6021]) );
  DFF ram_reg_1295__4_ ( .D(n10261), .CP(wclk), .Q(ram[6020]) );
  DFF ram_reg_1295__3_ ( .D(n10260), .CP(wclk), .Q(ram[6019]) );
  DFF ram_reg_1295__2_ ( .D(n10259), .CP(wclk), .Q(ram[6018]) );
  DFF ram_reg_1295__1_ ( .D(n10258), .CP(wclk), .Q(ram[6017]) );
  DFF ram_reg_1295__0_ ( .D(n10257), .CP(wclk), .Q(ram[6016]) );
  DFF ram_reg_1299__7_ ( .D(n10232), .CP(wclk), .Q(ram[5991]) );
  DFF ram_reg_1299__6_ ( .D(n10231), .CP(wclk), .Q(ram[5990]) );
  DFF ram_reg_1299__5_ ( .D(n10230), .CP(wclk), .Q(ram[5989]) );
  DFF ram_reg_1299__4_ ( .D(n10229), .CP(wclk), .Q(ram[5988]) );
  DFF ram_reg_1299__3_ ( .D(n10228), .CP(wclk), .Q(ram[5987]) );
  DFF ram_reg_1299__2_ ( .D(n10227), .CP(wclk), .Q(ram[5986]) );
  DFF ram_reg_1299__1_ ( .D(n10226), .CP(wclk), .Q(ram[5985]) );
  DFF ram_reg_1299__0_ ( .D(n10225), .CP(wclk), .Q(ram[5984]) );
  DFF ram_reg_1307__7_ ( .D(n10168), .CP(wclk), .Q(ram[5927]) );
  DFF ram_reg_1307__6_ ( .D(n10167), .CP(wclk), .Q(ram[5926]) );
  DFF ram_reg_1307__5_ ( .D(n10166), .CP(wclk), .Q(ram[5925]) );
  DFF ram_reg_1307__4_ ( .D(n10165), .CP(wclk), .Q(ram[5924]) );
  DFF ram_reg_1307__3_ ( .D(n10164), .CP(wclk), .Q(ram[5923]) );
  DFF ram_reg_1307__2_ ( .D(n10163), .CP(wclk), .Q(ram[5922]) );
  DFF ram_reg_1307__1_ ( .D(n10162), .CP(wclk), .Q(ram[5921]) );
  DFF ram_reg_1307__0_ ( .D(n10161), .CP(wclk), .Q(ram[5920]) );
  DFF ram_reg_1311__7_ ( .D(n10136), .CP(wclk), .Q(ram[5895]) );
  DFF ram_reg_1311__6_ ( .D(n10135), .CP(wclk), .Q(ram[5894]) );
  DFF ram_reg_1311__5_ ( .D(n10134), .CP(wclk), .Q(ram[5893]) );
  DFF ram_reg_1311__4_ ( .D(n10133), .CP(wclk), .Q(ram[5892]) );
  DFF ram_reg_1311__3_ ( .D(n10132), .CP(wclk), .Q(ram[5891]) );
  DFF ram_reg_1311__2_ ( .D(n10131), .CP(wclk), .Q(ram[5890]) );
  DFF ram_reg_1311__1_ ( .D(n10130), .CP(wclk), .Q(ram[5889]) );
  DFF ram_reg_1311__0_ ( .D(n10129), .CP(wclk), .Q(ram[5888]) );
  DFF ram_reg_1315__7_ ( .D(n10104), .CP(wclk), .Q(ram[5863]) );
  DFF ram_reg_1315__6_ ( .D(n10103), .CP(wclk), .Q(ram[5862]) );
  DFF ram_reg_1315__5_ ( .D(n10102), .CP(wclk), .Q(ram[5861]) );
  DFF ram_reg_1315__4_ ( .D(n10101), .CP(wclk), .Q(ram[5860]) );
  DFF ram_reg_1315__3_ ( .D(n10100), .CP(wclk), .Q(ram[5859]) );
  DFF ram_reg_1315__2_ ( .D(n10099), .CP(wclk), .Q(ram[5858]) );
  DFF ram_reg_1315__1_ ( .D(n10098), .CP(wclk), .Q(ram[5857]) );
  DFF ram_reg_1315__0_ ( .D(n10097), .CP(wclk), .Q(ram[5856]) );
  DFF ram_reg_1323__7_ ( .D(n10040), .CP(wclk), .Q(ram[5799]) );
  DFF ram_reg_1323__6_ ( .D(n10039), .CP(wclk), .Q(ram[5798]) );
  DFF ram_reg_1323__5_ ( .D(n10038), .CP(wclk), .Q(ram[5797]) );
  DFF ram_reg_1323__4_ ( .D(n10037), .CP(wclk), .Q(ram[5796]) );
  DFF ram_reg_1323__3_ ( .D(n10036), .CP(wclk), .Q(ram[5795]) );
  DFF ram_reg_1323__2_ ( .D(n10035), .CP(wclk), .Q(ram[5794]) );
  DFF ram_reg_1323__1_ ( .D(n10034), .CP(wclk), .Q(ram[5793]) );
  DFF ram_reg_1323__0_ ( .D(n10033), .CP(wclk), .Q(ram[5792]) );
  DFF ram_reg_1327__7_ ( .D(n10008), .CP(wclk), .Q(ram[5767]) );
  DFF ram_reg_1327__6_ ( .D(n10007), .CP(wclk), .Q(ram[5766]) );
  DFF ram_reg_1327__5_ ( .D(n10006), .CP(wclk), .Q(ram[5765]) );
  DFF ram_reg_1327__4_ ( .D(n10005), .CP(wclk), .Q(ram[5764]) );
  DFF ram_reg_1327__3_ ( .D(n10004), .CP(wclk), .Q(ram[5763]) );
  DFF ram_reg_1327__2_ ( .D(n10003), .CP(wclk), .Q(ram[5762]) );
  DFF ram_reg_1327__1_ ( .D(n10002), .CP(wclk), .Q(ram[5761]) );
  DFF ram_reg_1327__0_ ( .D(n10001), .CP(wclk), .Q(ram[5760]) );
  DFF ram_reg_1331__7_ ( .D(n9976), .CP(wclk), .Q(ram[5735]) );
  DFF ram_reg_1331__6_ ( .D(n9975), .CP(wclk), .Q(ram[5734]) );
  DFF ram_reg_1331__5_ ( .D(n9974), .CP(wclk), .Q(ram[5733]) );
  DFF ram_reg_1331__4_ ( .D(n9973), .CP(wclk), .Q(ram[5732]) );
  DFF ram_reg_1331__3_ ( .D(n9972), .CP(wclk), .Q(ram[5731]) );
  DFF ram_reg_1331__2_ ( .D(n9971), .CP(wclk), .Q(ram[5730]) );
  DFF ram_reg_1331__1_ ( .D(n9970), .CP(wclk), .Q(ram[5729]) );
  DFF ram_reg_1331__0_ ( .D(n9969), .CP(wclk), .Q(ram[5728]) );
  DFF ram_reg_1335__7_ ( .D(n9944), .CP(wclk), .Q(ram[5703]) );
  DFF ram_reg_1335__6_ ( .D(n9943), .CP(wclk), .Q(ram[5702]) );
  DFF ram_reg_1335__5_ ( .D(n9942), .CP(wclk), .Q(ram[5701]) );
  DFF ram_reg_1335__4_ ( .D(n9941), .CP(wclk), .Q(ram[5700]) );
  DFF ram_reg_1335__3_ ( .D(n9940), .CP(wclk), .Q(ram[5699]) );
  DFF ram_reg_1335__2_ ( .D(n9939), .CP(wclk), .Q(ram[5698]) );
  DFF ram_reg_1335__1_ ( .D(n9938), .CP(wclk), .Q(ram[5697]) );
  DFF ram_reg_1335__0_ ( .D(n9937), .CP(wclk), .Q(ram[5696]) );
  DFF ram_reg_1339__7_ ( .D(n9912), .CP(wclk), .Q(ram[5671]) );
  DFF ram_reg_1339__6_ ( .D(n9911), .CP(wclk), .Q(ram[5670]) );
  DFF ram_reg_1339__5_ ( .D(n9910), .CP(wclk), .Q(ram[5669]) );
  DFF ram_reg_1339__4_ ( .D(n9909), .CP(wclk), .Q(ram[5668]) );
  DFF ram_reg_1339__3_ ( .D(n9908), .CP(wclk), .Q(ram[5667]) );
  DFF ram_reg_1339__2_ ( .D(n9907), .CP(wclk), .Q(ram[5666]) );
  DFF ram_reg_1339__1_ ( .D(n9906), .CP(wclk), .Q(ram[5665]) );
  DFF ram_reg_1339__0_ ( .D(n9905), .CP(wclk), .Q(ram[5664]) );
  DFF ram_reg_1343__7_ ( .D(n9880), .CP(wclk), .Q(ram[5639]) );
  DFF ram_reg_1343__6_ ( .D(n9879), .CP(wclk), .Q(ram[5638]) );
  DFF ram_reg_1343__5_ ( .D(n9878), .CP(wclk), .Q(ram[5637]) );
  DFF ram_reg_1343__4_ ( .D(n9877), .CP(wclk), .Q(ram[5636]) );
  DFF ram_reg_1343__3_ ( .D(n9876), .CP(wclk), .Q(ram[5635]) );
  DFF ram_reg_1343__2_ ( .D(n9875), .CP(wclk), .Q(ram[5634]) );
  DFF ram_reg_1343__1_ ( .D(n9874), .CP(wclk), .Q(ram[5633]) );
  DFF ram_reg_1343__0_ ( .D(n9873), .CP(wclk), .Q(ram[5632]) );
  DFF ram_reg_1355__7_ ( .D(n9784), .CP(wclk), .Q(ram[5543]) );
  DFF ram_reg_1355__6_ ( .D(n9783), .CP(wclk), .Q(ram[5542]) );
  DFF ram_reg_1355__5_ ( .D(n9782), .CP(wclk), .Q(ram[5541]) );
  DFF ram_reg_1355__4_ ( .D(n9781), .CP(wclk), .Q(ram[5540]) );
  DFF ram_reg_1355__3_ ( .D(n9780), .CP(wclk), .Q(ram[5539]) );
  DFF ram_reg_1355__2_ ( .D(n9779), .CP(wclk), .Q(ram[5538]) );
  DFF ram_reg_1355__1_ ( .D(n9778), .CP(wclk), .Q(ram[5537]) );
  DFF ram_reg_1355__0_ ( .D(n9777), .CP(wclk), .Q(ram[5536]) );
  DFF ram_reg_1359__7_ ( .D(n9752), .CP(wclk), .Q(ram[5511]) );
  DFF ram_reg_1359__6_ ( .D(n9751), .CP(wclk), .Q(ram[5510]) );
  DFF ram_reg_1359__5_ ( .D(n9750), .CP(wclk), .Q(ram[5509]) );
  DFF ram_reg_1359__4_ ( .D(n9749), .CP(wclk), .Q(ram[5508]) );
  DFF ram_reg_1359__3_ ( .D(n9748), .CP(wclk), .Q(ram[5507]) );
  DFF ram_reg_1359__2_ ( .D(n9747), .CP(wclk), .Q(ram[5506]) );
  DFF ram_reg_1359__1_ ( .D(n9746), .CP(wclk), .Q(ram[5505]) );
  DFF ram_reg_1359__0_ ( .D(n9745), .CP(wclk), .Q(ram[5504]) );
  DFF ram_reg_1371__7_ ( .D(n9656), .CP(wclk), .Q(ram[5415]) );
  DFF ram_reg_1371__6_ ( .D(n9655), .CP(wclk), .Q(ram[5414]) );
  DFF ram_reg_1371__5_ ( .D(n9654), .CP(wclk), .Q(ram[5413]) );
  DFF ram_reg_1371__4_ ( .D(n9653), .CP(wclk), .Q(ram[5412]) );
  DFF ram_reg_1371__3_ ( .D(n9652), .CP(wclk), .Q(ram[5411]) );
  DFF ram_reg_1371__2_ ( .D(n9651), .CP(wclk), .Q(ram[5410]) );
  DFF ram_reg_1371__1_ ( .D(n9650), .CP(wclk), .Q(ram[5409]) );
  DFF ram_reg_1371__0_ ( .D(n9649), .CP(wclk), .Q(ram[5408]) );
  DFF ram_reg_1387__7_ ( .D(n9528), .CP(wclk), .Q(ram[5287]) );
  DFF ram_reg_1387__6_ ( .D(n9527), .CP(wclk), .Q(ram[5286]) );
  DFF ram_reg_1387__5_ ( .D(n9526), .CP(wclk), .Q(ram[5285]) );
  DFF ram_reg_1387__4_ ( .D(n9525), .CP(wclk), .Q(ram[5284]) );
  DFF ram_reg_1387__3_ ( .D(n9524), .CP(wclk), .Q(ram[5283]) );
  DFF ram_reg_1387__2_ ( .D(n9523), .CP(wclk), .Q(ram[5282]) );
  DFF ram_reg_1387__1_ ( .D(n9522), .CP(wclk), .Q(ram[5281]) );
  DFF ram_reg_1387__0_ ( .D(n9521), .CP(wclk), .Q(ram[5280]) );
  DFF ram_reg_1391__7_ ( .D(n9496), .CP(wclk), .Q(ram[5255]) );
  DFF ram_reg_1391__6_ ( .D(n9495), .CP(wclk), .Q(ram[5254]) );
  DFF ram_reg_1391__5_ ( .D(n9494), .CP(wclk), .Q(ram[5253]) );
  DFF ram_reg_1391__4_ ( .D(n9493), .CP(wclk), .Q(ram[5252]) );
  DFF ram_reg_1391__3_ ( .D(n9492), .CP(wclk), .Q(ram[5251]) );
  DFF ram_reg_1391__2_ ( .D(n9491), .CP(wclk), .Q(ram[5250]) );
  DFF ram_reg_1391__1_ ( .D(n9490), .CP(wclk), .Q(ram[5249]) );
  DFF ram_reg_1391__0_ ( .D(n9489), .CP(wclk), .Q(ram[5248]) );
  DFF ram_reg_1395__7_ ( .D(n9464), .CP(wclk), .Q(ram[5223]) );
  DFF ram_reg_1395__6_ ( .D(n9463), .CP(wclk), .Q(ram[5222]) );
  DFF ram_reg_1395__5_ ( .D(n9462), .CP(wclk), .Q(ram[5221]) );
  DFF ram_reg_1395__4_ ( .D(n9461), .CP(wclk), .Q(ram[5220]) );
  DFF ram_reg_1395__3_ ( .D(n9460), .CP(wclk), .Q(ram[5219]) );
  DFF ram_reg_1395__2_ ( .D(n9459), .CP(wclk), .Q(ram[5218]) );
  DFF ram_reg_1395__1_ ( .D(n9458), .CP(wclk), .Q(ram[5217]) );
  DFF ram_reg_1395__0_ ( .D(n9457), .CP(wclk), .Q(ram[5216]) );
  DFF ram_reg_1403__7_ ( .D(n9400), .CP(wclk), .Q(ram[5159]) );
  DFF ram_reg_1403__6_ ( .D(n9399), .CP(wclk), .Q(ram[5158]) );
  DFF ram_reg_1403__5_ ( .D(n9398), .CP(wclk), .Q(ram[5157]) );
  DFF ram_reg_1403__4_ ( .D(n9397), .CP(wclk), .Q(ram[5156]) );
  DFF ram_reg_1403__3_ ( .D(n9396), .CP(wclk), .Q(ram[5155]) );
  DFF ram_reg_1403__2_ ( .D(n9395), .CP(wclk), .Q(ram[5154]) );
  DFF ram_reg_1403__1_ ( .D(n9394), .CP(wclk), .Q(ram[5153]) );
  DFF ram_reg_1403__0_ ( .D(n9393), .CP(wclk), .Q(ram[5152]) );
  DFF ram_reg_1407__7_ ( .D(n9368), .CP(wclk), .Q(ram[5127]) );
  DFF ram_reg_1407__6_ ( .D(n9367), .CP(wclk), .Q(ram[5126]) );
  DFF ram_reg_1407__5_ ( .D(n9366), .CP(wclk), .Q(ram[5125]) );
  DFF ram_reg_1407__4_ ( .D(n9365), .CP(wclk), .Q(ram[5124]) );
  DFF ram_reg_1407__3_ ( .D(n9364), .CP(wclk), .Q(ram[5123]) );
  DFF ram_reg_1407__2_ ( .D(n9363), .CP(wclk), .Q(ram[5122]) );
  DFF ram_reg_1407__1_ ( .D(n9362), .CP(wclk), .Q(ram[5121]) );
  DFF ram_reg_1407__0_ ( .D(n9361), .CP(wclk), .Q(ram[5120]) );
  DFF ram_reg_1411__7_ ( .D(n9336), .CP(wclk), .Q(ram[5095]) );
  DFF ram_reg_1411__6_ ( .D(n9335), .CP(wclk), .Q(ram[5094]) );
  DFF ram_reg_1411__5_ ( .D(n9334), .CP(wclk), .Q(ram[5093]) );
  DFF ram_reg_1411__4_ ( .D(n9333), .CP(wclk), .Q(ram[5092]) );
  DFF ram_reg_1411__3_ ( .D(n9332), .CP(wclk), .Q(ram[5091]) );
  DFF ram_reg_1411__2_ ( .D(n9331), .CP(wclk), .Q(ram[5090]) );
  DFF ram_reg_1411__1_ ( .D(n9330), .CP(wclk), .Q(ram[5089]) );
  DFF ram_reg_1411__0_ ( .D(n9329), .CP(wclk), .Q(ram[5088]) );
  DFF ram_reg_1415__7_ ( .D(n9304), .CP(wclk), .Q(ram[5063]) );
  DFF ram_reg_1415__6_ ( .D(n9303), .CP(wclk), .Q(ram[5062]) );
  DFF ram_reg_1415__5_ ( .D(n9302), .CP(wclk), .Q(ram[5061]) );
  DFF ram_reg_1415__4_ ( .D(n9301), .CP(wclk), .Q(ram[5060]) );
  DFF ram_reg_1415__3_ ( .D(n9300), .CP(wclk), .Q(ram[5059]) );
  DFF ram_reg_1415__2_ ( .D(n9299), .CP(wclk), .Q(ram[5058]) );
  DFF ram_reg_1415__1_ ( .D(n9298), .CP(wclk), .Q(ram[5057]) );
  DFF ram_reg_1415__0_ ( .D(n9297), .CP(wclk), .Q(ram[5056]) );
  DFF ram_reg_1419__7_ ( .D(n9272), .CP(wclk), .Q(ram[5031]) );
  DFF ram_reg_1419__6_ ( .D(n9271), .CP(wclk), .Q(ram[5030]) );
  DFF ram_reg_1419__5_ ( .D(n9270), .CP(wclk), .Q(ram[5029]) );
  DFF ram_reg_1419__4_ ( .D(n9269), .CP(wclk), .Q(ram[5028]) );
  DFF ram_reg_1419__3_ ( .D(n9268), .CP(wclk), .Q(ram[5027]) );
  DFF ram_reg_1419__2_ ( .D(n9267), .CP(wclk), .Q(ram[5026]) );
  DFF ram_reg_1419__1_ ( .D(n9266), .CP(wclk), .Q(ram[5025]) );
  DFF ram_reg_1419__0_ ( .D(n9265), .CP(wclk), .Q(ram[5024]) );
  DFF ram_reg_1423__7_ ( .D(n9240), .CP(wclk), .Q(ram[4999]) );
  DFF ram_reg_1423__6_ ( .D(n9239), .CP(wclk), .Q(ram[4998]) );
  DFF ram_reg_1423__5_ ( .D(n9238), .CP(wclk), .Q(ram[4997]) );
  DFF ram_reg_1423__4_ ( .D(n9237), .CP(wclk), .Q(ram[4996]) );
  DFF ram_reg_1423__3_ ( .D(n9236), .CP(wclk), .Q(ram[4995]) );
  DFF ram_reg_1423__2_ ( .D(n9235), .CP(wclk), .Q(ram[4994]) );
  DFF ram_reg_1423__1_ ( .D(n9234), .CP(wclk), .Q(ram[4993]) );
  DFF ram_reg_1423__0_ ( .D(n9233), .CP(wclk), .Q(ram[4992]) );
  DFF ram_reg_1427__7_ ( .D(n9208), .CP(wclk), .Q(ram[4967]) );
  DFF ram_reg_1427__6_ ( .D(n9207), .CP(wclk), .Q(ram[4966]) );
  DFF ram_reg_1427__5_ ( .D(n9206), .CP(wclk), .Q(ram[4965]) );
  DFF ram_reg_1427__4_ ( .D(n9205), .CP(wclk), .Q(ram[4964]) );
  DFF ram_reg_1427__3_ ( .D(n9204), .CP(wclk), .Q(ram[4963]) );
  DFF ram_reg_1427__2_ ( .D(n9203), .CP(wclk), .Q(ram[4962]) );
  DFF ram_reg_1427__1_ ( .D(n9202), .CP(wclk), .Q(ram[4961]) );
  DFF ram_reg_1427__0_ ( .D(n9201), .CP(wclk), .Q(ram[4960]) );
  DFF ram_reg_1431__7_ ( .D(n9176), .CP(wclk), .Q(ram[4935]) );
  DFF ram_reg_1431__6_ ( .D(n9175), .CP(wclk), .Q(ram[4934]) );
  DFF ram_reg_1431__5_ ( .D(n9174), .CP(wclk), .Q(ram[4933]) );
  DFF ram_reg_1431__4_ ( .D(n9173), .CP(wclk), .Q(ram[4932]) );
  DFF ram_reg_1431__3_ ( .D(n9172), .CP(wclk), .Q(ram[4931]) );
  DFF ram_reg_1431__2_ ( .D(n9171), .CP(wclk), .Q(ram[4930]) );
  DFF ram_reg_1431__1_ ( .D(n9170), .CP(wclk), .Q(ram[4929]) );
  DFF ram_reg_1431__0_ ( .D(n9169), .CP(wclk), .Q(ram[4928]) );
  DFF ram_reg_1435__7_ ( .D(n9144), .CP(wclk), .Q(ram[4903]) );
  DFF ram_reg_1435__6_ ( .D(n9143), .CP(wclk), .Q(ram[4902]) );
  DFF ram_reg_1435__5_ ( .D(n9142), .CP(wclk), .Q(ram[4901]) );
  DFF ram_reg_1435__4_ ( .D(n9141), .CP(wclk), .Q(ram[4900]) );
  DFF ram_reg_1435__3_ ( .D(n9140), .CP(wclk), .Q(ram[4899]) );
  DFF ram_reg_1435__2_ ( .D(n9139), .CP(wclk), .Q(ram[4898]) );
  DFF ram_reg_1435__1_ ( .D(n9138), .CP(wclk), .Q(ram[4897]) );
  DFF ram_reg_1435__0_ ( .D(n9137), .CP(wclk), .Q(ram[4896]) );
  DFF ram_reg_1439__7_ ( .D(n9112), .CP(wclk), .Q(ram[4871]) );
  DFF ram_reg_1439__6_ ( .D(n9111), .CP(wclk), .Q(ram[4870]) );
  DFF ram_reg_1439__5_ ( .D(n9110), .CP(wclk), .Q(ram[4869]) );
  DFF ram_reg_1439__4_ ( .D(n9109), .CP(wclk), .Q(ram[4868]) );
  DFF ram_reg_1439__3_ ( .D(n9108), .CP(wclk), .Q(ram[4867]) );
  DFF ram_reg_1439__2_ ( .D(n9107), .CP(wclk), .Q(ram[4866]) );
  DFF ram_reg_1439__1_ ( .D(n9106), .CP(wclk), .Q(ram[4865]) );
  DFF ram_reg_1439__0_ ( .D(n9105), .CP(wclk), .Q(ram[4864]) );
  DFF ram_reg_1443__7_ ( .D(n9080), .CP(wclk), .Q(ram[4839]) );
  DFF ram_reg_1443__6_ ( .D(n9079), .CP(wclk), .Q(ram[4838]) );
  DFF ram_reg_1443__5_ ( .D(n9078), .CP(wclk), .Q(ram[4837]) );
  DFF ram_reg_1443__4_ ( .D(n9077), .CP(wclk), .Q(ram[4836]) );
  DFF ram_reg_1443__3_ ( .D(n9076), .CP(wclk), .Q(ram[4835]) );
  DFF ram_reg_1443__2_ ( .D(n9075), .CP(wclk), .Q(ram[4834]) );
  DFF ram_reg_1443__1_ ( .D(n9074), .CP(wclk), .Q(ram[4833]) );
  DFF ram_reg_1443__0_ ( .D(n9073), .CP(wclk), .Q(ram[4832]) );
  DFF ram_reg_1447__7_ ( .D(n9048), .CP(wclk), .Q(ram[4807]) );
  DFF ram_reg_1447__6_ ( .D(n9047), .CP(wclk), .Q(ram[4806]) );
  DFF ram_reg_1447__5_ ( .D(n9046), .CP(wclk), .Q(ram[4805]) );
  DFF ram_reg_1447__4_ ( .D(n9045), .CP(wclk), .Q(ram[4804]) );
  DFF ram_reg_1447__3_ ( .D(n9044), .CP(wclk), .Q(ram[4803]) );
  DFF ram_reg_1447__2_ ( .D(n9043), .CP(wclk), .Q(ram[4802]) );
  DFF ram_reg_1447__1_ ( .D(n9042), .CP(wclk), .Q(ram[4801]) );
  DFF ram_reg_1447__0_ ( .D(n9041), .CP(wclk), .Q(ram[4800]) );
  DFF ram_reg_1451__7_ ( .D(n9016), .CP(wclk), .Q(ram[4775]) );
  DFF ram_reg_1451__6_ ( .D(n9015), .CP(wclk), .Q(ram[4774]) );
  DFF ram_reg_1451__5_ ( .D(n9014), .CP(wclk), .Q(ram[4773]) );
  DFF ram_reg_1451__4_ ( .D(n9013), .CP(wclk), .Q(ram[4772]) );
  DFF ram_reg_1451__3_ ( .D(n9012), .CP(wclk), .Q(ram[4771]) );
  DFF ram_reg_1451__2_ ( .D(n9011), .CP(wclk), .Q(ram[4770]) );
  DFF ram_reg_1451__1_ ( .D(n9010), .CP(wclk), .Q(ram[4769]) );
  DFF ram_reg_1451__0_ ( .D(n9009), .CP(wclk), .Q(ram[4768]) );
  DFF ram_reg_1455__7_ ( .D(n8984), .CP(wclk), .Q(ram[4743]) );
  DFF ram_reg_1455__6_ ( .D(n8983), .CP(wclk), .Q(ram[4742]) );
  DFF ram_reg_1455__5_ ( .D(n8982), .CP(wclk), .Q(ram[4741]) );
  DFF ram_reg_1455__4_ ( .D(n8981), .CP(wclk), .Q(ram[4740]) );
  DFF ram_reg_1455__3_ ( .D(n8980), .CP(wclk), .Q(ram[4739]) );
  DFF ram_reg_1455__2_ ( .D(n8979), .CP(wclk), .Q(ram[4738]) );
  DFF ram_reg_1455__1_ ( .D(n8978), .CP(wclk), .Q(ram[4737]) );
  DFF ram_reg_1455__0_ ( .D(n8977), .CP(wclk), .Q(ram[4736]) );
  DFF ram_reg_1459__7_ ( .D(n8952), .CP(wclk), .Q(ram[4711]) );
  DFF ram_reg_1459__6_ ( .D(n8951), .CP(wclk), .Q(ram[4710]) );
  DFF ram_reg_1459__5_ ( .D(n8950), .CP(wclk), .Q(ram[4709]) );
  DFF ram_reg_1459__4_ ( .D(n8949), .CP(wclk), .Q(ram[4708]) );
  DFF ram_reg_1459__3_ ( .D(n8948), .CP(wclk), .Q(ram[4707]) );
  DFF ram_reg_1459__2_ ( .D(n8947), .CP(wclk), .Q(ram[4706]) );
  DFF ram_reg_1459__1_ ( .D(n8946), .CP(wclk), .Q(ram[4705]) );
  DFF ram_reg_1459__0_ ( .D(n8945), .CP(wclk), .Q(ram[4704]) );
  DFF ram_reg_1463__7_ ( .D(n8920), .CP(wclk), .Q(ram[4679]) );
  DFF ram_reg_1463__6_ ( .D(n8919), .CP(wclk), .Q(ram[4678]) );
  DFF ram_reg_1463__5_ ( .D(n8918), .CP(wclk), .Q(ram[4677]) );
  DFF ram_reg_1463__4_ ( .D(n8917), .CP(wclk), .Q(ram[4676]) );
  DFF ram_reg_1463__3_ ( .D(n8916), .CP(wclk), .Q(ram[4675]) );
  DFF ram_reg_1463__2_ ( .D(n8915), .CP(wclk), .Q(ram[4674]) );
  DFF ram_reg_1463__1_ ( .D(n8914), .CP(wclk), .Q(ram[4673]) );
  DFF ram_reg_1463__0_ ( .D(n8913), .CP(wclk), .Q(ram[4672]) );
  DFF ram_reg_1467__7_ ( .D(n8888), .CP(wclk), .Q(ram[4647]) );
  DFF ram_reg_1467__6_ ( .D(n8887), .CP(wclk), .Q(ram[4646]) );
  DFF ram_reg_1467__5_ ( .D(n8886), .CP(wclk), .Q(ram[4645]) );
  DFF ram_reg_1467__4_ ( .D(n8885), .CP(wclk), .Q(ram[4644]) );
  DFF ram_reg_1467__3_ ( .D(n8884), .CP(wclk), .Q(ram[4643]) );
  DFF ram_reg_1467__2_ ( .D(n8883), .CP(wclk), .Q(ram[4642]) );
  DFF ram_reg_1467__1_ ( .D(n8882), .CP(wclk), .Q(ram[4641]) );
  DFF ram_reg_1467__0_ ( .D(n8881), .CP(wclk), .Q(ram[4640]) );
  DFF ram_reg_1471__7_ ( .D(n8856), .CP(wclk), .Q(ram[4615]) );
  DFF ram_reg_1471__6_ ( .D(n8855), .CP(wclk), .Q(ram[4614]) );
  DFF ram_reg_1471__5_ ( .D(n8854), .CP(wclk), .Q(ram[4613]) );
  DFF ram_reg_1471__4_ ( .D(n8853), .CP(wclk), .Q(ram[4612]) );
  DFF ram_reg_1471__3_ ( .D(n8852), .CP(wclk), .Q(ram[4611]) );
  DFF ram_reg_1471__2_ ( .D(n8851), .CP(wclk), .Q(ram[4610]) );
  DFF ram_reg_1471__1_ ( .D(n8850), .CP(wclk), .Q(ram[4609]) );
  DFF ram_reg_1471__0_ ( .D(n8849), .CP(wclk), .Q(ram[4608]) );
  DFF ram_reg_1475__7_ ( .D(n8824), .CP(wclk), .Q(ram[4583]) );
  DFF ram_reg_1475__6_ ( .D(n8823), .CP(wclk), .Q(ram[4582]) );
  DFF ram_reg_1475__5_ ( .D(n8822), .CP(wclk), .Q(ram[4581]) );
  DFF ram_reg_1475__4_ ( .D(n8821), .CP(wclk), .Q(ram[4580]) );
  DFF ram_reg_1475__3_ ( .D(n8820), .CP(wclk), .Q(ram[4579]) );
  DFF ram_reg_1475__2_ ( .D(n8819), .CP(wclk), .Q(ram[4578]) );
  DFF ram_reg_1475__1_ ( .D(n8818), .CP(wclk), .Q(ram[4577]) );
  DFF ram_reg_1475__0_ ( .D(n8817), .CP(wclk), .Q(ram[4576]) );
  DFF ram_reg_1479__7_ ( .D(n8792), .CP(wclk), .Q(ram[4551]) );
  DFF ram_reg_1479__6_ ( .D(n8791), .CP(wclk), .Q(ram[4550]) );
  DFF ram_reg_1479__5_ ( .D(n8790), .CP(wclk), .Q(ram[4549]) );
  DFF ram_reg_1479__4_ ( .D(n8789), .CP(wclk), .Q(ram[4548]) );
  DFF ram_reg_1479__3_ ( .D(n8788), .CP(wclk), .Q(ram[4547]) );
  DFF ram_reg_1479__2_ ( .D(n8787), .CP(wclk), .Q(ram[4546]) );
  DFF ram_reg_1479__1_ ( .D(n8786), .CP(wclk), .Q(ram[4545]) );
  DFF ram_reg_1479__0_ ( .D(n8785), .CP(wclk), .Q(ram[4544]) );
  DFF ram_reg_1483__7_ ( .D(n8760), .CP(wclk), .Q(ram[4519]) );
  DFF ram_reg_1483__6_ ( .D(n8759), .CP(wclk), .Q(ram[4518]) );
  DFF ram_reg_1483__5_ ( .D(n8758), .CP(wclk), .Q(ram[4517]) );
  DFF ram_reg_1483__4_ ( .D(n8757), .CP(wclk), .Q(ram[4516]) );
  DFF ram_reg_1483__3_ ( .D(n8756), .CP(wclk), .Q(ram[4515]) );
  DFF ram_reg_1483__2_ ( .D(n8755), .CP(wclk), .Q(ram[4514]) );
  DFF ram_reg_1483__1_ ( .D(n8754), .CP(wclk), .Q(ram[4513]) );
  DFF ram_reg_1483__0_ ( .D(n8753), .CP(wclk), .Q(ram[4512]) );
  DFF ram_reg_1487__7_ ( .D(n8728), .CP(wclk), .Q(ram[4487]) );
  DFF ram_reg_1487__6_ ( .D(n8727), .CP(wclk), .Q(ram[4486]) );
  DFF ram_reg_1487__5_ ( .D(n8726), .CP(wclk), .Q(ram[4485]) );
  DFF ram_reg_1487__4_ ( .D(n8725), .CP(wclk), .Q(ram[4484]) );
  DFF ram_reg_1487__3_ ( .D(n8724), .CP(wclk), .Q(ram[4483]) );
  DFF ram_reg_1487__2_ ( .D(n8723), .CP(wclk), .Q(ram[4482]) );
  DFF ram_reg_1487__1_ ( .D(n8722), .CP(wclk), .Q(ram[4481]) );
  DFF ram_reg_1487__0_ ( .D(n8721), .CP(wclk), .Q(ram[4480]) );
  DFF ram_reg_1491__7_ ( .D(n8696), .CP(wclk), .Q(ram[4455]) );
  DFF ram_reg_1491__6_ ( .D(n8695), .CP(wclk), .Q(ram[4454]) );
  DFF ram_reg_1491__5_ ( .D(n8694), .CP(wclk), .Q(ram[4453]) );
  DFF ram_reg_1491__4_ ( .D(n8693), .CP(wclk), .Q(ram[4452]) );
  DFF ram_reg_1491__3_ ( .D(n8692), .CP(wclk), .Q(ram[4451]) );
  DFF ram_reg_1491__2_ ( .D(n8691), .CP(wclk), .Q(ram[4450]) );
  DFF ram_reg_1491__1_ ( .D(n8690), .CP(wclk), .Q(ram[4449]) );
  DFF ram_reg_1491__0_ ( .D(n8689), .CP(wclk), .Q(ram[4448]) );
  DFF ram_reg_1499__7_ ( .D(n8632), .CP(wclk), .Q(ram[4391]) );
  DFF ram_reg_1499__6_ ( .D(n8631), .CP(wclk), .Q(ram[4390]) );
  DFF ram_reg_1499__5_ ( .D(n8630), .CP(wclk), .Q(ram[4389]) );
  DFF ram_reg_1499__4_ ( .D(n8629), .CP(wclk), .Q(ram[4388]) );
  DFF ram_reg_1499__3_ ( .D(n8628), .CP(wclk), .Q(ram[4387]) );
  DFF ram_reg_1499__2_ ( .D(n8627), .CP(wclk), .Q(ram[4386]) );
  DFF ram_reg_1499__1_ ( .D(n8626), .CP(wclk), .Q(ram[4385]) );
  DFF ram_reg_1499__0_ ( .D(n8625), .CP(wclk), .Q(ram[4384]) );
  DFF ram_reg_1503__7_ ( .D(n8600), .CP(wclk), .Q(ram[4359]) );
  DFF ram_reg_1503__6_ ( .D(n8599), .CP(wclk), .Q(ram[4358]) );
  DFF ram_reg_1503__5_ ( .D(n8598), .CP(wclk), .Q(ram[4357]) );
  DFF ram_reg_1503__4_ ( .D(n8597), .CP(wclk), .Q(ram[4356]) );
  DFF ram_reg_1503__3_ ( .D(n8596), .CP(wclk), .Q(ram[4355]) );
  DFF ram_reg_1503__2_ ( .D(n8595), .CP(wclk), .Q(ram[4354]) );
  DFF ram_reg_1503__1_ ( .D(n8594), .CP(wclk), .Q(ram[4353]) );
  DFF ram_reg_1503__0_ ( .D(n8593), .CP(wclk), .Q(ram[4352]) );
  DFF ram_reg_1507__7_ ( .D(n8568), .CP(wclk), .Q(ram[4327]) );
  DFF ram_reg_1507__6_ ( .D(n8567), .CP(wclk), .Q(ram[4326]) );
  DFF ram_reg_1507__5_ ( .D(n8566), .CP(wclk), .Q(ram[4325]) );
  DFF ram_reg_1507__4_ ( .D(n8565), .CP(wclk), .Q(ram[4324]) );
  DFF ram_reg_1507__3_ ( .D(n8564), .CP(wclk), .Q(ram[4323]) );
  DFF ram_reg_1507__2_ ( .D(n8563), .CP(wclk), .Q(ram[4322]) );
  DFF ram_reg_1507__1_ ( .D(n8562), .CP(wclk), .Q(ram[4321]) );
  DFF ram_reg_1507__0_ ( .D(n8561), .CP(wclk), .Q(ram[4320]) );
  DFF ram_reg_1511__7_ ( .D(n8536), .CP(wclk), .Q(ram[4295]) );
  DFF ram_reg_1511__6_ ( .D(n8535), .CP(wclk), .Q(ram[4294]) );
  DFF ram_reg_1511__5_ ( .D(n8534), .CP(wclk), .Q(ram[4293]) );
  DFF ram_reg_1511__4_ ( .D(n8533), .CP(wclk), .Q(ram[4292]) );
  DFF ram_reg_1511__3_ ( .D(n8532), .CP(wclk), .Q(ram[4291]) );
  DFF ram_reg_1511__2_ ( .D(n8531), .CP(wclk), .Q(ram[4290]) );
  DFF ram_reg_1511__1_ ( .D(n8530), .CP(wclk), .Q(ram[4289]) );
  DFF ram_reg_1511__0_ ( .D(n8529), .CP(wclk), .Q(ram[4288]) );
  DFF ram_reg_1515__7_ ( .D(n8504), .CP(wclk), .Q(ram[4263]) );
  DFF ram_reg_1515__6_ ( .D(n8503), .CP(wclk), .Q(ram[4262]) );
  DFF ram_reg_1515__5_ ( .D(n8502), .CP(wclk), .Q(ram[4261]) );
  DFF ram_reg_1515__4_ ( .D(n8501), .CP(wclk), .Q(ram[4260]) );
  DFF ram_reg_1515__3_ ( .D(n8500), .CP(wclk), .Q(ram[4259]) );
  DFF ram_reg_1515__2_ ( .D(n8499), .CP(wclk), .Q(ram[4258]) );
  DFF ram_reg_1515__1_ ( .D(n8498), .CP(wclk), .Q(ram[4257]) );
  DFF ram_reg_1515__0_ ( .D(n8497), .CP(wclk), .Q(ram[4256]) );
  DFF ram_reg_1519__7_ ( .D(n8472), .CP(wclk), .Q(ram[4231]) );
  DFF ram_reg_1519__6_ ( .D(n8471), .CP(wclk), .Q(ram[4230]) );
  DFF ram_reg_1519__5_ ( .D(n8470), .CP(wclk), .Q(ram[4229]) );
  DFF ram_reg_1519__4_ ( .D(n8469), .CP(wclk), .Q(ram[4228]) );
  DFF ram_reg_1519__3_ ( .D(n8468), .CP(wclk), .Q(ram[4227]) );
  DFF ram_reg_1519__2_ ( .D(n8467), .CP(wclk), .Q(ram[4226]) );
  DFF ram_reg_1519__1_ ( .D(n8466), .CP(wclk), .Q(ram[4225]) );
  DFF ram_reg_1519__0_ ( .D(n8465), .CP(wclk), .Q(ram[4224]) );
  DFF ram_reg_1523__7_ ( .D(n8440), .CP(wclk), .Q(ram[4199]) );
  DFF ram_reg_1523__6_ ( .D(n8439), .CP(wclk), .Q(ram[4198]) );
  DFF ram_reg_1523__5_ ( .D(n8438), .CP(wclk), .Q(ram[4197]) );
  DFF ram_reg_1523__4_ ( .D(n8437), .CP(wclk), .Q(ram[4196]) );
  DFF ram_reg_1523__3_ ( .D(n8436), .CP(wclk), .Q(ram[4195]) );
  DFF ram_reg_1523__2_ ( .D(n8435), .CP(wclk), .Q(ram[4194]) );
  DFF ram_reg_1523__1_ ( .D(n8434), .CP(wclk), .Q(ram[4193]) );
  DFF ram_reg_1523__0_ ( .D(n8433), .CP(wclk), .Q(ram[4192]) );
  DFF ram_reg_1527__7_ ( .D(n8408), .CP(wclk), .Q(ram[4167]) );
  DFF ram_reg_1527__6_ ( .D(n8407), .CP(wclk), .Q(ram[4166]) );
  DFF ram_reg_1527__5_ ( .D(n8406), .CP(wclk), .Q(ram[4165]) );
  DFF ram_reg_1527__4_ ( .D(n8405), .CP(wclk), .Q(ram[4164]) );
  DFF ram_reg_1527__3_ ( .D(n8404), .CP(wclk), .Q(ram[4163]) );
  DFF ram_reg_1527__2_ ( .D(n8403), .CP(wclk), .Q(ram[4162]) );
  DFF ram_reg_1527__1_ ( .D(n8402), .CP(wclk), .Q(ram[4161]) );
  DFF ram_reg_1527__0_ ( .D(n8401), .CP(wclk), .Q(ram[4160]) );
  DFF ram_reg_1531__7_ ( .D(n8376), .CP(wclk), .Q(ram[4135]) );
  DFF ram_reg_1531__6_ ( .D(n8375), .CP(wclk), .Q(ram[4134]) );
  DFF ram_reg_1531__5_ ( .D(n8374), .CP(wclk), .Q(ram[4133]) );
  DFF ram_reg_1531__4_ ( .D(n8373), .CP(wclk), .Q(ram[4132]) );
  DFF ram_reg_1531__3_ ( .D(n8372), .CP(wclk), .Q(ram[4131]) );
  DFF ram_reg_1531__2_ ( .D(n8371), .CP(wclk), .Q(ram[4130]) );
  DFF ram_reg_1531__1_ ( .D(n8370), .CP(wclk), .Q(ram[4129]) );
  DFF ram_reg_1531__0_ ( .D(n8369), .CP(wclk), .Q(ram[4128]) );
  DFF ram_reg_1535__7_ ( .D(n8344), .CP(wclk), .Q(ram[4103]) );
  DFF ram_reg_1535__6_ ( .D(n8343), .CP(wclk), .Q(ram[4102]) );
  DFF ram_reg_1535__5_ ( .D(n8342), .CP(wclk), .Q(ram[4101]) );
  DFF ram_reg_1535__4_ ( .D(n8341), .CP(wclk), .Q(ram[4100]) );
  DFF ram_reg_1535__3_ ( .D(n8340), .CP(wclk), .Q(ram[4099]) );
  DFF ram_reg_1535__2_ ( .D(n8339), .CP(wclk), .Q(ram[4098]) );
  DFF ram_reg_1535__1_ ( .D(n8338), .CP(wclk), .Q(ram[4097]) );
  DFF ram_reg_1535__0_ ( .D(n8337), .CP(wclk), .Q(ram[4096]) );
  DFF ram_reg_1547__7_ ( .D(n8248), .CP(wclk), .Q(ram[4007]) );
  DFF ram_reg_1547__6_ ( .D(n8247), .CP(wclk), .Q(ram[4006]) );
  DFF ram_reg_1547__5_ ( .D(n8246), .CP(wclk), .Q(ram[4005]) );
  DFF ram_reg_1547__4_ ( .D(n8245), .CP(wclk), .Q(ram[4004]) );
  DFF ram_reg_1547__3_ ( .D(n8244), .CP(wclk), .Q(ram[4003]) );
  DFF ram_reg_1547__2_ ( .D(n8243), .CP(wclk), .Q(ram[4002]) );
  DFF ram_reg_1547__1_ ( .D(n8242), .CP(wclk), .Q(ram[4001]) );
  DFF ram_reg_1547__0_ ( .D(n8241), .CP(wclk), .Q(ram[4000]) );
  DFF ram_reg_1551__7_ ( .D(n8216), .CP(wclk), .Q(ram[3975]) );
  DFF ram_reg_1551__6_ ( .D(n8215), .CP(wclk), .Q(ram[3974]) );
  DFF ram_reg_1551__5_ ( .D(n8214), .CP(wclk), .Q(ram[3973]) );
  DFF ram_reg_1551__4_ ( .D(n8213), .CP(wclk), .Q(ram[3972]) );
  DFF ram_reg_1551__3_ ( .D(n8212), .CP(wclk), .Q(ram[3971]) );
  DFF ram_reg_1551__2_ ( .D(n8211), .CP(wclk), .Q(ram[3970]) );
  DFF ram_reg_1551__1_ ( .D(n8210), .CP(wclk), .Q(ram[3969]) );
  DFF ram_reg_1551__0_ ( .D(n8209), .CP(wclk), .Q(ram[3968]) );
  DFF ram_reg_1563__7_ ( .D(n8120), .CP(wclk), .Q(ram[3879]) );
  DFF ram_reg_1563__6_ ( .D(n8119), .CP(wclk), .Q(ram[3878]) );
  DFF ram_reg_1563__5_ ( .D(n8118), .CP(wclk), .Q(ram[3877]) );
  DFF ram_reg_1563__4_ ( .D(n8117), .CP(wclk), .Q(ram[3876]) );
  DFF ram_reg_1563__3_ ( .D(n8116), .CP(wclk), .Q(ram[3875]) );
  DFF ram_reg_1563__2_ ( .D(n8115), .CP(wclk), .Q(ram[3874]) );
  DFF ram_reg_1563__1_ ( .D(n8114), .CP(wclk), .Q(ram[3873]) );
  DFF ram_reg_1563__0_ ( .D(n8113), .CP(wclk), .Q(ram[3872]) );
  DFF ram_reg_1571__7_ ( .D(n8056), .CP(wclk), .Q(ram[3815]) );
  DFF ram_reg_1571__6_ ( .D(n8055), .CP(wclk), .Q(ram[3814]) );
  DFF ram_reg_1571__5_ ( .D(n8054), .CP(wclk), .Q(ram[3813]) );
  DFF ram_reg_1571__4_ ( .D(n8053), .CP(wclk), .Q(ram[3812]) );
  DFF ram_reg_1571__3_ ( .D(n8052), .CP(wclk), .Q(ram[3811]) );
  DFF ram_reg_1571__2_ ( .D(n8051), .CP(wclk), .Q(ram[3810]) );
  DFF ram_reg_1571__1_ ( .D(n8050), .CP(wclk), .Q(ram[3809]) );
  DFF ram_reg_1571__0_ ( .D(n8049), .CP(wclk), .Q(ram[3808]) );
  DFF ram_reg_1579__7_ ( .D(n7992), .CP(wclk), .Q(ram[3751]) );
  DFF ram_reg_1579__6_ ( .D(n7991), .CP(wclk), .Q(ram[3750]) );
  DFF ram_reg_1579__5_ ( .D(n7990), .CP(wclk), .Q(ram[3749]) );
  DFF ram_reg_1579__4_ ( .D(n7989), .CP(wclk), .Q(ram[3748]) );
  DFF ram_reg_1579__3_ ( .D(n7988), .CP(wclk), .Q(ram[3747]) );
  DFF ram_reg_1579__2_ ( .D(n7987), .CP(wclk), .Q(ram[3746]) );
  DFF ram_reg_1579__1_ ( .D(n7986), .CP(wclk), .Q(ram[3745]) );
  DFF ram_reg_1579__0_ ( .D(n7985), .CP(wclk), .Q(ram[3744]) );
  DFF ram_reg_1583__7_ ( .D(n7960), .CP(wclk), .Q(ram[3719]) );
  DFF ram_reg_1583__6_ ( .D(n7959), .CP(wclk), .Q(ram[3718]) );
  DFF ram_reg_1583__5_ ( .D(n7958), .CP(wclk), .Q(ram[3717]) );
  DFF ram_reg_1583__4_ ( .D(n7957), .CP(wclk), .Q(ram[3716]) );
  DFF ram_reg_1583__3_ ( .D(n7956), .CP(wclk), .Q(ram[3715]) );
  DFF ram_reg_1583__2_ ( .D(n7955), .CP(wclk), .Q(ram[3714]) );
  DFF ram_reg_1583__1_ ( .D(n7954), .CP(wclk), .Q(ram[3713]) );
  DFF ram_reg_1583__0_ ( .D(n7953), .CP(wclk), .Q(ram[3712]) );
  DFF ram_reg_1587__7_ ( .D(n7928), .CP(wclk), .Q(ram[3687]) );
  DFF ram_reg_1587__6_ ( .D(n7927), .CP(wclk), .Q(ram[3686]) );
  DFF ram_reg_1587__5_ ( .D(n7926), .CP(wclk), .Q(ram[3685]) );
  DFF ram_reg_1587__4_ ( .D(n7925), .CP(wclk), .Q(ram[3684]) );
  DFF ram_reg_1587__3_ ( .D(n7924), .CP(wclk), .Q(ram[3683]) );
  DFF ram_reg_1587__2_ ( .D(n7923), .CP(wclk), .Q(ram[3682]) );
  DFF ram_reg_1587__1_ ( .D(n7922), .CP(wclk), .Q(ram[3681]) );
  DFF ram_reg_1587__0_ ( .D(n7921), .CP(wclk), .Q(ram[3680]) );
  DFF ram_reg_1595__7_ ( .D(n7864), .CP(wclk), .Q(ram[3623]) );
  DFF ram_reg_1595__6_ ( .D(n7863), .CP(wclk), .Q(ram[3622]) );
  DFF ram_reg_1595__5_ ( .D(n7862), .CP(wclk), .Q(ram[3621]) );
  DFF ram_reg_1595__4_ ( .D(n7861), .CP(wclk), .Q(ram[3620]) );
  DFF ram_reg_1595__3_ ( .D(n7860), .CP(wclk), .Q(ram[3619]) );
  DFF ram_reg_1595__2_ ( .D(n7859), .CP(wclk), .Q(ram[3618]) );
  DFF ram_reg_1595__1_ ( .D(n7858), .CP(wclk), .Q(ram[3617]) );
  DFF ram_reg_1595__0_ ( .D(n7857), .CP(wclk), .Q(ram[3616]) );
  DFF ram_reg_1599__7_ ( .D(n7832), .CP(wclk), .Q(ram[3591]) );
  DFF ram_reg_1599__6_ ( .D(n7831), .CP(wclk), .Q(ram[3590]) );
  DFF ram_reg_1599__5_ ( .D(n7830), .CP(wclk), .Q(ram[3589]) );
  DFF ram_reg_1599__4_ ( .D(n7829), .CP(wclk), .Q(ram[3588]) );
  DFF ram_reg_1599__3_ ( .D(n7828), .CP(wclk), .Q(ram[3587]) );
  DFF ram_reg_1599__2_ ( .D(n7827), .CP(wclk), .Q(ram[3586]) );
  DFF ram_reg_1599__1_ ( .D(n7826), .CP(wclk), .Q(ram[3585]) );
  DFF ram_reg_1599__0_ ( .D(n7825), .CP(wclk), .Q(ram[3584]) );
  DFF ram_reg_1643__7_ ( .D(n7480), .CP(wclk), .Q(ram[3239]) );
  DFF ram_reg_1643__6_ ( .D(n7479), .CP(wclk), .Q(ram[3238]) );
  DFF ram_reg_1643__5_ ( .D(n7478), .CP(wclk), .Q(ram[3237]) );
  DFF ram_reg_1643__4_ ( .D(n7477), .CP(wclk), .Q(ram[3236]) );
  DFF ram_reg_1643__3_ ( .D(n7476), .CP(wclk), .Q(ram[3235]) );
  DFF ram_reg_1643__2_ ( .D(n7475), .CP(wclk), .Q(ram[3234]) );
  DFF ram_reg_1643__1_ ( .D(n7474), .CP(wclk), .Q(ram[3233]) );
  DFF ram_reg_1643__0_ ( .D(n7473), .CP(wclk), .Q(ram[3232]) );
  DFF ram_reg_1659__7_ ( .D(n7352), .CP(wclk), .Q(ram[3111]) );
  DFF ram_reg_1659__6_ ( .D(n7351), .CP(wclk), .Q(ram[3110]) );
  DFF ram_reg_1659__5_ ( .D(n7350), .CP(wclk), .Q(ram[3109]) );
  DFF ram_reg_1659__4_ ( .D(n7349), .CP(wclk), .Q(ram[3108]) );
  DFF ram_reg_1659__3_ ( .D(n7348), .CP(wclk), .Q(ram[3107]) );
  DFF ram_reg_1659__2_ ( .D(n7347), .CP(wclk), .Q(ram[3106]) );
  DFF ram_reg_1659__1_ ( .D(n7346), .CP(wclk), .Q(ram[3105]) );
  DFF ram_reg_1659__0_ ( .D(n7345), .CP(wclk), .Q(ram[3104]) );
  DFF ram_reg_1663__7_ ( .D(n7320), .CP(wclk), .Q(ram[3079]) );
  DFF ram_reg_1663__6_ ( .D(n7319), .CP(wclk), .Q(ram[3078]) );
  DFF ram_reg_1663__5_ ( .D(n7318), .CP(wclk), .Q(ram[3077]) );
  DFF ram_reg_1663__4_ ( .D(n7317), .CP(wclk), .Q(ram[3076]) );
  DFF ram_reg_1663__3_ ( .D(n7316), .CP(wclk), .Q(ram[3075]) );
  DFF ram_reg_1663__2_ ( .D(n7315), .CP(wclk), .Q(ram[3074]) );
  DFF ram_reg_1663__1_ ( .D(n7314), .CP(wclk), .Q(ram[3073]) );
  DFF ram_reg_1663__0_ ( .D(n7313), .CP(wclk), .Q(ram[3072]) );
  DFF ram_reg_1667__7_ ( .D(n7288), .CP(wclk), .Q(ram[3047]) );
  DFF ram_reg_1667__6_ ( .D(n7287), .CP(wclk), .Q(ram[3046]) );
  DFF ram_reg_1667__5_ ( .D(n7286), .CP(wclk), .Q(ram[3045]) );
  DFF ram_reg_1667__4_ ( .D(n7285), .CP(wclk), .Q(ram[3044]) );
  DFF ram_reg_1667__3_ ( .D(n7284), .CP(wclk), .Q(ram[3043]) );
  DFF ram_reg_1667__2_ ( .D(n7283), .CP(wclk), .Q(ram[3042]) );
  DFF ram_reg_1667__1_ ( .D(n7282), .CP(wclk), .Q(ram[3041]) );
  DFF ram_reg_1667__0_ ( .D(n7281), .CP(wclk), .Q(ram[3040]) );
  DFF ram_reg_1675__7_ ( .D(n7224), .CP(wclk), .Q(ram[2983]) );
  DFF ram_reg_1675__6_ ( .D(n7223), .CP(wclk), .Q(ram[2982]) );
  DFF ram_reg_1675__5_ ( .D(n7222), .CP(wclk), .Q(ram[2981]) );
  DFF ram_reg_1675__4_ ( .D(n7221), .CP(wclk), .Q(ram[2980]) );
  DFF ram_reg_1675__3_ ( .D(n7220), .CP(wclk), .Q(ram[2979]) );
  DFF ram_reg_1675__2_ ( .D(n7219), .CP(wclk), .Q(ram[2978]) );
  DFF ram_reg_1675__1_ ( .D(n7218), .CP(wclk), .Q(ram[2977]) );
  DFF ram_reg_1675__0_ ( .D(n7217), .CP(wclk), .Q(ram[2976]) );
  DFF ram_reg_1679__7_ ( .D(n7192), .CP(wclk), .Q(ram[2951]) );
  DFF ram_reg_1679__6_ ( .D(n7191), .CP(wclk), .Q(ram[2950]) );
  DFF ram_reg_1679__5_ ( .D(n7190), .CP(wclk), .Q(ram[2949]) );
  DFF ram_reg_1679__4_ ( .D(n7189), .CP(wclk), .Q(ram[2948]) );
  DFF ram_reg_1679__3_ ( .D(n7188), .CP(wclk), .Q(ram[2947]) );
  DFF ram_reg_1679__2_ ( .D(n7187), .CP(wclk), .Q(ram[2946]) );
  DFF ram_reg_1679__1_ ( .D(n7186), .CP(wclk), .Q(ram[2945]) );
  DFF ram_reg_1679__0_ ( .D(n7185), .CP(wclk), .Q(ram[2944]) );
  DFF ram_reg_1683__7_ ( .D(n7160), .CP(wclk), .Q(ram[2919]) );
  DFF ram_reg_1683__6_ ( .D(n7159), .CP(wclk), .Q(ram[2918]) );
  DFF ram_reg_1683__5_ ( .D(n7158), .CP(wclk), .Q(ram[2917]) );
  DFF ram_reg_1683__4_ ( .D(n7157), .CP(wclk), .Q(ram[2916]) );
  DFF ram_reg_1683__3_ ( .D(n7156), .CP(wclk), .Q(ram[2915]) );
  DFF ram_reg_1683__2_ ( .D(n7155), .CP(wclk), .Q(ram[2914]) );
  DFF ram_reg_1683__1_ ( .D(n7154), .CP(wclk), .Q(ram[2913]) );
  DFF ram_reg_1683__0_ ( .D(n7153), .CP(wclk), .Q(ram[2912]) );
  DFF ram_reg_1691__7_ ( .D(n7096), .CP(wclk), .Q(ram[2855]) );
  DFF ram_reg_1691__6_ ( .D(n7095), .CP(wclk), .Q(ram[2854]) );
  DFF ram_reg_1691__5_ ( .D(n7094), .CP(wclk), .Q(ram[2853]) );
  DFF ram_reg_1691__4_ ( .D(n7093), .CP(wclk), .Q(ram[2852]) );
  DFF ram_reg_1691__3_ ( .D(n7092), .CP(wclk), .Q(ram[2851]) );
  DFF ram_reg_1691__2_ ( .D(n7091), .CP(wclk), .Q(ram[2850]) );
  DFF ram_reg_1691__1_ ( .D(n7090), .CP(wclk), .Q(ram[2849]) );
  DFF ram_reg_1691__0_ ( .D(n7089), .CP(wclk), .Q(ram[2848]) );
  DFF ram_reg_1695__7_ ( .D(n7064), .CP(wclk), .Q(ram[2823]) );
  DFF ram_reg_1695__6_ ( .D(n7063), .CP(wclk), .Q(ram[2822]) );
  DFF ram_reg_1695__5_ ( .D(n7062), .CP(wclk), .Q(ram[2821]) );
  DFF ram_reg_1695__4_ ( .D(n7061), .CP(wclk), .Q(ram[2820]) );
  DFF ram_reg_1695__3_ ( .D(n7060), .CP(wclk), .Q(ram[2819]) );
  DFF ram_reg_1695__2_ ( .D(n7059), .CP(wclk), .Q(ram[2818]) );
  DFF ram_reg_1695__1_ ( .D(n7058), .CP(wclk), .Q(ram[2817]) );
  DFF ram_reg_1695__0_ ( .D(n7057), .CP(wclk), .Q(ram[2816]) );
  DFF ram_reg_1699__7_ ( .D(n7032), .CP(wclk), .Q(ram[2791]) );
  DFF ram_reg_1699__6_ ( .D(n7031), .CP(wclk), .Q(ram[2790]) );
  DFF ram_reg_1699__5_ ( .D(n7030), .CP(wclk), .Q(ram[2789]) );
  DFF ram_reg_1699__4_ ( .D(n7029), .CP(wclk), .Q(ram[2788]) );
  DFF ram_reg_1699__3_ ( .D(n7028), .CP(wclk), .Q(ram[2787]) );
  DFF ram_reg_1699__2_ ( .D(n7027), .CP(wclk), .Q(ram[2786]) );
  DFF ram_reg_1699__1_ ( .D(n7026), .CP(wclk), .Q(ram[2785]) );
  DFF ram_reg_1699__0_ ( .D(n7025), .CP(wclk), .Q(ram[2784]) );
  DFF ram_reg_1703__7_ ( .D(n7000), .CP(wclk), .Q(ram[2759]) );
  DFF ram_reg_1703__6_ ( .D(n6999), .CP(wclk), .Q(ram[2758]) );
  DFF ram_reg_1703__5_ ( .D(n6998), .CP(wclk), .Q(ram[2757]) );
  DFF ram_reg_1703__4_ ( .D(n6997), .CP(wclk), .Q(ram[2756]) );
  DFF ram_reg_1703__3_ ( .D(n6996), .CP(wclk), .Q(ram[2755]) );
  DFF ram_reg_1703__2_ ( .D(n6995), .CP(wclk), .Q(ram[2754]) );
  DFF ram_reg_1703__1_ ( .D(n6994), .CP(wclk), .Q(ram[2753]) );
  DFF ram_reg_1703__0_ ( .D(n6993), .CP(wclk), .Q(ram[2752]) );
  DFF ram_reg_1707__7_ ( .D(n6968), .CP(wclk), .Q(ram[2727]) );
  DFF ram_reg_1707__6_ ( .D(n6967), .CP(wclk), .Q(ram[2726]) );
  DFF ram_reg_1707__5_ ( .D(n6966), .CP(wclk), .Q(ram[2725]) );
  DFF ram_reg_1707__4_ ( .D(n6965), .CP(wclk), .Q(ram[2724]) );
  DFF ram_reg_1707__3_ ( .D(n6964), .CP(wclk), .Q(ram[2723]) );
  DFF ram_reg_1707__2_ ( .D(n6963), .CP(wclk), .Q(ram[2722]) );
  DFF ram_reg_1707__1_ ( .D(n6962), .CP(wclk), .Q(ram[2721]) );
  DFF ram_reg_1707__0_ ( .D(n6961), .CP(wclk), .Q(ram[2720]) );
  DFF ram_reg_1711__7_ ( .D(n6936), .CP(wclk), .Q(ram[2695]) );
  DFF ram_reg_1711__6_ ( .D(n6935), .CP(wclk), .Q(ram[2694]) );
  DFF ram_reg_1711__5_ ( .D(n6934), .CP(wclk), .Q(ram[2693]) );
  DFF ram_reg_1711__4_ ( .D(n6933), .CP(wclk), .Q(ram[2692]) );
  DFF ram_reg_1711__3_ ( .D(n6932), .CP(wclk), .Q(ram[2691]) );
  DFF ram_reg_1711__2_ ( .D(n6931), .CP(wclk), .Q(ram[2690]) );
  DFF ram_reg_1711__1_ ( .D(n6930), .CP(wclk), .Q(ram[2689]) );
  DFF ram_reg_1711__0_ ( .D(n6929), .CP(wclk), .Q(ram[2688]) );
  DFF ram_reg_1715__7_ ( .D(n6904), .CP(wclk), .Q(ram[2663]) );
  DFF ram_reg_1715__6_ ( .D(n6903), .CP(wclk), .Q(ram[2662]) );
  DFF ram_reg_1715__5_ ( .D(n6902), .CP(wclk), .Q(ram[2661]) );
  DFF ram_reg_1715__4_ ( .D(n6901), .CP(wclk), .Q(ram[2660]) );
  DFF ram_reg_1715__3_ ( .D(n6900), .CP(wclk), .Q(ram[2659]) );
  DFF ram_reg_1715__2_ ( .D(n6899), .CP(wclk), .Q(ram[2658]) );
  DFF ram_reg_1715__1_ ( .D(n6898), .CP(wclk), .Q(ram[2657]) );
  DFF ram_reg_1715__0_ ( .D(n6897), .CP(wclk), .Q(ram[2656]) );
  DFF ram_reg_1719__7_ ( .D(n6872), .CP(wclk), .Q(ram[2631]) );
  DFF ram_reg_1719__6_ ( .D(n6871), .CP(wclk), .Q(ram[2630]) );
  DFF ram_reg_1719__5_ ( .D(n6870), .CP(wclk), .Q(ram[2629]) );
  DFF ram_reg_1719__4_ ( .D(n6869), .CP(wclk), .Q(ram[2628]) );
  DFF ram_reg_1719__3_ ( .D(n6868), .CP(wclk), .Q(ram[2627]) );
  DFF ram_reg_1719__2_ ( .D(n6867), .CP(wclk), .Q(ram[2626]) );
  DFF ram_reg_1719__1_ ( .D(n6866), .CP(wclk), .Q(ram[2625]) );
  DFF ram_reg_1719__0_ ( .D(n6865), .CP(wclk), .Q(ram[2624]) );
  DFF ram_reg_1723__7_ ( .D(n6840), .CP(wclk), .Q(ram[2599]) );
  DFF ram_reg_1723__6_ ( .D(n6839), .CP(wclk), .Q(ram[2598]) );
  DFF ram_reg_1723__5_ ( .D(n6838), .CP(wclk), .Q(ram[2597]) );
  DFF ram_reg_1723__4_ ( .D(n6837), .CP(wclk), .Q(ram[2596]) );
  DFF ram_reg_1723__3_ ( .D(n6836), .CP(wclk), .Q(ram[2595]) );
  DFF ram_reg_1723__2_ ( .D(n6835), .CP(wclk), .Q(ram[2594]) );
  DFF ram_reg_1723__1_ ( .D(n6834), .CP(wclk), .Q(ram[2593]) );
  DFF ram_reg_1723__0_ ( .D(n6833), .CP(wclk), .Q(ram[2592]) );
  DFF ram_reg_1727__7_ ( .D(n6808), .CP(wclk), .Q(ram[2567]) );
  DFF ram_reg_1727__6_ ( .D(n6807), .CP(wclk), .Q(ram[2566]) );
  DFF ram_reg_1727__5_ ( .D(n6806), .CP(wclk), .Q(ram[2565]) );
  DFF ram_reg_1727__4_ ( .D(n6805), .CP(wclk), .Q(ram[2564]) );
  DFF ram_reg_1727__3_ ( .D(n6804), .CP(wclk), .Q(ram[2563]) );
  DFF ram_reg_1727__2_ ( .D(n6803), .CP(wclk), .Q(ram[2562]) );
  DFF ram_reg_1727__1_ ( .D(n6802), .CP(wclk), .Q(ram[2561]) );
  DFF ram_reg_1727__0_ ( .D(n6801), .CP(wclk), .Q(ram[2560]) );
  DFF ram_reg_1731__7_ ( .D(n6776), .CP(wclk), .Q(ram[2535]) );
  DFF ram_reg_1731__6_ ( .D(n6775), .CP(wclk), .Q(ram[2534]) );
  DFF ram_reg_1731__5_ ( .D(n6774), .CP(wclk), .Q(ram[2533]) );
  DFF ram_reg_1731__4_ ( .D(n6773), .CP(wclk), .Q(ram[2532]) );
  DFF ram_reg_1731__3_ ( .D(n6772), .CP(wclk), .Q(ram[2531]) );
  DFF ram_reg_1731__2_ ( .D(n6771), .CP(wclk), .Q(ram[2530]) );
  DFF ram_reg_1731__1_ ( .D(n6770), .CP(wclk), .Q(ram[2529]) );
  DFF ram_reg_1731__0_ ( .D(n6769), .CP(wclk), .Q(ram[2528]) );
  DFF ram_reg_1739__7_ ( .D(n6712), .CP(wclk), .Q(ram[2471]) );
  DFF ram_reg_1739__6_ ( .D(n6711), .CP(wclk), .Q(ram[2470]) );
  DFF ram_reg_1739__5_ ( .D(n6710), .CP(wclk), .Q(ram[2469]) );
  DFF ram_reg_1739__4_ ( .D(n6709), .CP(wclk), .Q(ram[2468]) );
  DFF ram_reg_1739__3_ ( .D(n6708), .CP(wclk), .Q(ram[2467]) );
  DFF ram_reg_1739__2_ ( .D(n6707), .CP(wclk), .Q(ram[2466]) );
  DFF ram_reg_1739__1_ ( .D(n6706), .CP(wclk), .Q(ram[2465]) );
  DFF ram_reg_1739__0_ ( .D(n6705), .CP(wclk), .Q(ram[2464]) );
  DFF ram_reg_1743__7_ ( .D(n6680), .CP(wclk), .Q(ram[2439]) );
  DFF ram_reg_1743__6_ ( .D(n6679), .CP(wclk), .Q(ram[2438]) );
  DFF ram_reg_1743__5_ ( .D(n6678), .CP(wclk), .Q(ram[2437]) );
  DFF ram_reg_1743__4_ ( .D(n6677), .CP(wclk), .Q(ram[2436]) );
  DFF ram_reg_1743__3_ ( .D(n6676), .CP(wclk), .Q(ram[2435]) );
  DFF ram_reg_1743__2_ ( .D(n6675), .CP(wclk), .Q(ram[2434]) );
  DFF ram_reg_1743__1_ ( .D(n6674), .CP(wclk), .Q(ram[2433]) );
  DFF ram_reg_1743__0_ ( .D(n6673), .CP(wclk), .Q(ram[2432]) );
  DFF ram_reg_1755__7_ ( .D(n6584), .CP(wclk), .Q(ram[2343]) );
  DFF ram_reg_1755__6_ ( .D(n6583), .CP(wclk), .Q(ram[2342]) );
  DFF ram_reg_1755__5_ ( .D(n6582), .CP(wclk), .Q(ram[2341]) );
  DFF ram_reg_1755__4_ ( .D(n6581), .CP(wclk), .Q(ram[2340]) );
  DFF ram_reg_1755__3_ ( .D(n6580), .CP(wclk), .Q(ram[2339]) );
  DFF ram_reg_1755__2_ ( .D(n6579), .CP(wclk), .Q(ram[2338]) );
  DFF ram_reg_1755__1_ ( .D(n6578), .CP(wclk), .Q(ram[2337]) );
  DFF ram_reg_1755__0_ ( .D(n6577), .CP(wclk), .Q(ram[2336]) );
  DFF ram_reg_1759__7_ ( .D(n6552), .CP(wclk), .Q(ram[2311]) );
  DFF ram_reg_1759__6_ ( .D(n6551), .CP(wclk), .Q(ram[2310]) );
  DFF ram_reg_1759__5_ ( .D(n6550), .CP(wclk), .Q(ram[2309]) );
  DFF ram_reg_1759__4_ ( .D(n6549), .CP(wclk), .Q(ram[2308]) );
  DFF ram_reg_1759__3_ ( .D(n6548), .CP(wclk), .Q(ram[2307]) );
  DFF ram_reg_1759__2_ ( .D(n6547), .CP(wclk), .Q(ram[2306]) );
  DFF ram_reg_1759__1_ ( .D(n6546), .CP(wclk), .Q(ram[2305]) );
  DFF ram_reg_1759__0_ ( .D(n6545), .CP(wclk), .Q(ram[2304]) );
  DFF ram_reg_1763__7_ ( .D(n6520), .CP(wclk), .Q(ram[2279]) );
  DFF ram_reg_1763__6_ ( .D(n6519), .CP(wclk), .Q(ram[2278]) );
  DFF ram_reg_1763__5_ ( .D(n6518), .CP(wclk), .Q(ram[2277]) );
  DFF ram_reg_1763__4_ ( .D(n6517), .CP(wclk), .Q(ram[2276]) );
  DFF ram_reg_1763__3_ ( .D(n6516), .CP(wclk), .Q(ram[2275]) );
  DFF ram_reg_1763__2_ ( .D(n6515), .CP(wclk), .Q(ram[2274]) );
  DFF ram_reg_1763__1_ ( .D(n6514), .CP(wclk), .Q(ram[2273]) );
  DFF ram_reg_1763__0_ ( .D(n6513), .CP(wclk), .Q(ram[2272]) );
  DFF ram_reg_1771__7_ ( .D(n6456), .CP(wclk), .Q(ram[2215]) );
  DFF ram_reg_1771__6_ ( .D(n6455), .CP(wclk), .Q(ram[2214]) );
  DFF ram_reg_1771__5_ ( .D(n6454), .CP(wclk), .Q(ram[2213]) );
  DFF ram_reg_1771__4_ ( .D(n6453), .CP(wclk), .Q(ram[2212]) );
  DFF ram_reg_1771__3_ ( .D(n6452), .CP(wclk), .Q(ram[2211]) );
  DFF ram_reg_1771__2_ ( .D(n6451), .CP(wclk), .Q(ram[2210]) );
  DFF ram_reg_1771__1_ ( .D(n6450), .CP(wclk), .Q(ram[2209]) );
  DFF ram_reg_1771__0_ ( .D(n6449), .CP(wclk), .Q(ram[2208]) );
  DFF ram_reg_1775__7_ ( .D(n6424), .CP(wclk), .Q(ram[2183]) );
  DFF ram_reg_1775__6_ ( .D(n6423), .CP(wclk), .Q(ram[2182]) );
  DFF ram_reg_1775__5_ ( .D(n6422), .CP(wclk), .Q(ram[2181]) );
  DFF ram_reg_1775__4_ ( .D(n6421), .CP(wclk), .Q(ram[2180]) );
  DFF ram_reg_1775__3_ ( .D(n6420), .CP(wclk), .Q(ram[2179]) );
  DFF ram_reg_1775__2_ ( .D(n6419), .CP(wclk), .Q(ram[2178]) );
  DFF ram_reg_1775__1_ ( .D(n6418), .CP(wclk), .Q(ram[2177]) );
  DFF ram_reg_1775__0_ ( .D(n6417), .CP(wclk), .Q(ram[2176]) );
  DFF ram_reg_1779__7_ ( .D(n6392), .CP(wclk), .Q(ram[2151]) );
  DFF ram_reg_1779__6_ ( .D(n6391), .CP(wclk), .Q(ram[2150]) );
  DFF ram_reg_1779__5_ ( .D(n6390), .CP(wclk), .Q(ram[2149]) );
  DFF ram_reg_1779__4_ ( .D(n6389), .CP(wclk), .Q(ram[2148]) );
  DFF ram_reg_1779__3_ ( .D(n6388), .CP(wclk), .Q(ram[2147]) );
  DFF ram_reg_1779__2_ ( .D(n6387), .CP(wclk), .Q(ram[2146]) );
  DFF ram_reg_1779__1_ ( .D(n6386), .CP(wclk), .Q(ram[2145]) );
  DFF ram_reg_1779__0_ ( .D(n6385), .CP(wclk), .Q(ram[2144]) );
  DFF ram_reg_1783__7_ ( .D(n6360), .CP(wclk), .Q(ram[2119]) );
  DFF ram_reg_1783__6_ ( .D(n6359), .CP(wclk), .Q(ram[2118]) );
  DFF ram_reg_1783__5_ ( .D(n6358), .CP(wclk), .Q(ram[2117]) );
  DFF ram_reg_1783__4_ ( .D(n6357), .CP(wclk), .Q(ram[2116]) );
  DFF ram_reg_1783__3_ ( .D(n6356), .CP(wclk), .Q(ram[2115]) );
  DFF ram_reg_1783__2_ ( .D(n6355), .CP(wclk), .Q(ram[2114]) );
  DFF ram_reg_1783__1_ ( .D(n6354), .CP(wclk), .Q(ram[2113]) );
  DFF ram_reg_1783__0_ ( .D(n6353), .CP(wclk), .Q(ram[2112]) );
  DFF ram_reg_1787__7_ ( .D(n6328), .CP(wclk), .Q(ram[2087]) );
  DFF ram_reg_1787__6_ ( .D(n6327), .CP(wclk), .Q(ram[2086]) );
  DFF ram_reg_1787__5_ ( .D(n6326), .CP(wclk), .Q(ram[2085]) );
  DFF ram_reg_1787__4_ ( .D(n6325), .CP(wclk), .Q(ram[2084]) );
  DFF ram_reg_1787__3_ ( .D(n6324), .CP(wclk), .Q(ram[2083]) );
  DFF ram_reg_1787__2_ ( .D(n6323), .CP(wclk), .Q(ram[2082]) );
  DFF ram_reg_1787__1_ ( .D(n6322), .CP(wclk), .Q(ram[2081]) );
  DFF ram_reg_1787__0_ ( .D(n6321), .CP(wclk), .Q(ram[2080]) );
  DFF ram_reg_1791__7_ ( .D(n6296), .CP(wclk), .Q(ram[2055]) );
  DFF ram_reg_1791__6_ ( .D(n6295), .CP(wclk), .Q(ram[2054]) );
  DFF ram_reg_1791__5_ ( .D(n6294), .CP(wclk), .Q(ram[2053]) );
  DFF ram_reg_1791__4_ ( .D(n6293), .CP(wclk), .Q(ram[2052]) );
  DFF ram_reg_1791__3_ ( .D(n6292), .CP(wclk), .Q(ram[2051]) );
  DFF ram_reg_1791__2_ ( .D(n6291), .CP(wclk), .Q(ram[2050]) );
  DFF ram_reg_1791__1_ ( .D(n6290), .CP(wclk), .Q(ram[2049]) );
  DFF ram_reg_1791__0_ ( .D(n6289), .CP(wclk), .Q(ram[2048]) );
  DFF ram_reg_1803__7_ ( .D(n6200), .CP(wclk), .Q(ram[1959]) );
  DFF ram_reg_1803__6_ ( .D(n6199), .CP(wclk), .Q(ram[1958]) );
  DFF ram_reg_1803__5_ ( .D(n6198), .CP(wclk), .Q(ram[1957]) );
  DFF ram_reg_1803__4_ ( .D(n6197), .CP(wclk), .Q(ram[1956]) );
  DFF ram_reg_1803__3_ ( .D(n6196), .CP(wclk), .Q(ram[1955]) );
  DFF ram_reg_1803__2_ ( .D(n6195), .CP(wclk), .Q(ram[1954]) );
  DFF ram_reg_1803__1_ ( .D(n6194), .CP(wclk), .Q(ram[1953]) );
  DFF ram_reg_1803__0_ ( .D(n6193), .CP(wclk), .Q(ram[1952]) );
  DFF ram_reg_1807__7_ ( .D(n6168), .CP(wclk), .Q(ram[1927]) );
  DFF ram_reg_1807__6_ ( .D(n6167), .CP(wclk), .Q(ram[1926]) );
  DFF ram_reg_1807__5_ ( .D(n6166), .CP(wclk), .Q(ram[1925]) );
  DFF ram_reg_1807__4_ ( .D(n6165), .CP(wclk), .Q(ram[1924]) );
  DFF ram_reg_1807__3_ ( .D(n6164), .CP(wclk), .Q(ram[1923]) );
  DFF ram_reg_1807__2_ ( .D(n6163), .CP(wclk), .Q(ram[1922]) );
  DFF ram_reg_1807__1_ ( .D(n6162), .CP(wclk), .Q(ram[1921]) );
  DFF ram_reg_1807__0_ ( .D(n6161), .CP(wclk), .Q(ram[1920]) );
  DFF ram_reg_1819__7_ ( .D(n6072), .CP(wclk), .Q(ram[1831]) );
  DFF ram_reg_1819__6_ ( .D(n6071), .CP(wclk), .Q(ram[1830]) );
  DFF ram_reg_1819__5_ ( .D(n6070), .CP(wclk), .Q(ram[1829]) );
  DFF ram_reg_1819__4_ ( .D(n6069), .CP(wclk), .Q(ram[1828]) );
  DFF ram_reg_1819__3_ ( .D(n6068), .CP(wclk), .Q(ram[1827]) );
  DFF ram_reg_1819__2_ ( .D(n6067), .CP(wclk), .Q(ram[1826]) );
  DFF ram_reg_1819__1_ ( .D(n6066), .CP(wclk), .Q(ram[1825]) );
  DFF ram_reg_1819__0_ ( .D(n6065), .CP(wclk), .Q(ram[1824]) );
  DFF ram_reg_1823__7_ ( .D(n6040), .CP(wclk), .Q(ram[1799]) );
  DFF ram_reg_1823__6_ ( .D(n6039), .CP(wclk), .Q(ram[1798]) );
  DFF ram_reg_1823__5_ ( .D(n6038), .CP(wclk), .Q(ram[1797]) );
  DFF ram_reg_1823__4_ ( .D(n6037), .CP(wclk), .Q(ram[1796]) );
  DFF ram_reg_1823__3_ ( .D(n6036), .CP(wclk), .Q(ram[1795]) );
  DFF ram_reg_1823__2_ ( .D(n6035), .CP(wclk), .Q(ram[1794]) );
  DFF ram_reg_1823__1_ ( .D(n6034), .CP(wclk), .Q(ram[1793]) );
  DFF ram_reg_1823__0_ ( .D(n6033), .CP(wclk), .Q(ram[1792]) );
  DFF ram_reg_1827__7_ ( .D(n6008), .CP(wclk), .Q(ram[1767]) );
  DFF ram_reg_1827__6_ ( .D(n6007), .CP(wclk), .Q(ram[1766]) );
  DFF ram_reg_1827__5_ ( .D(n6006), .CP(wclk), .Q(ram[1765]) );
  DFF ram_reg_1827__4_ ( .D(n6005), .CP(wclk), .Q(ram[1764]) );
  DFF ram_reg_1827__3_ ( .D(n6004), .CP(wclk), .Q(ram[1763]) );
  DFF ram_reg_1827__2_ ( .D(n6003), .CP(wclk), .Q(ram[1762]) );
  DFF ram_reg_1827__1_ ( .D(n6002), .CP(wclk), .Q(ram[1761]) );
  DFF ram_reg_1827__0_ ( .D(n6001), .CP(wclk), .Q(ram[1760]) );
  DFF ram_reg_1835__7_ ( .D(n5944), .CP(wclk), .Q(ram[1703]) );
  DFF ram_reg_1835__6_ ( .D(n5943), .CP(wclk), .Q(ram[1702]) );
  DFF ram_reg_1835__5_ ( .D(n5942), .CP(wclk), .Q(ram[1701]) );
  DFF ram_reg_1835__4_ ( .D(n5941), .CP(wclk), .Q(ram[1700]) );
  DFF ram_reg_1835__3_ ( .D(n5940), .CP(wclk), .Q(ram[1699]) );
  DFF ram_reg_1835__2_ ( .D(n5939), .CP(wclk), .Q(ram[1698]) );
  DFF ram_reg_1835__1_ ( .D(n5938), .CP(wclk), .Q(ram[1697]) );
  DFF ram_reg_1835__0_ ( .D(n5937), .CP(wclk), .Q(ram[1696]) );
  DFF ram_reg_1839__7_ ( .D(n5912), .CP(wclk), .Q(ram[1671]) );
  DFF ram_reg_1839__6_ ( .D(n5911), .CP(wclk), .Q(ram[1670]) );
  DFF ram_reg_1839__5_ ( .D(n5910), .CP(wclk), .Q(ram[1669]) );
  DFF ram_reg_1839__4_ ( .D(n5909), .CP(wclk), .Q(ram[1668]) );
  DFF ram_reg_1839__3_ ( .D(n5908), .CP(wclk), .Q(ram[1667]) );
  DFF ram_reg_1839__2_ ( .D(n5907), .CP(wclk), .Q(ram[1666]) );
  DFF ram_reg_1839__1_ ( .D(n5906), .CP(wclk), .Q(ram[1665]) );
  DFF ram_reg_1839__0_ ( .D(n5905), .CP(wclk), .Q(ram[1664]) );
  DFF ram_reg_1843__7_ ( .D(n5880), .CP(wclk), .Q(ram[1639]) );
  DFF ram_reg_1843__6_ ( .D(n5879), .CP(wclk), .Q(ram[1638]) );
  DFF ram_reg_1843__5_ ( .D(n5878), .CP(wclk), .Q(ram[1637]) );
  DFF ram_reg_1843__4_ ( .D(n5877), .CP(wclk), .Q(ram[1636]) );
  DFF ram_reg_1843__3_ ( .D(n5876), .CP(wclk), .Q(ram[1635]) );
  DFF ram_reg_1843__2_ ( .D(n5875), .CP(wclk), .Q(ram[1634]) );
  DFF ram_reg_1843__1_ ( .D(n5874), .CP(wclk), .Q(ram[1633]) );
  DFF ram_reg_1843__0_ ( .D(n5873), .CP(wclk), .Q(ram[1632]) );
  DFF ram_reg_1851__7_ ( .D(n5816), .CP(wclk), .Q(ram[1575]) );
  DFF ram_reg_1851__6_ ( .D(n5815), .CP(wclk), .Q(ram[1574]) );
  DFF ram_reg_1851__5_ ( .D(n5814), .CP(wclk), .Q(ram[1573]) );
  DFF ram_reg_1851__4_ ( .D(n5813), .CP(wclk), .Q(ram[1572]) );
  DFF ram_reg_1851__3_ ( .D(n5812), .CP(wclk), .Q(ram[1571]) );
  DFF ram_reg_1851__2_ ( .D(n5811), .CP(wclk), .Q(ram[1570]) );
  DFF ram_reg_1851__1_ ( .D(n5810), .CP(wclk), .Q(ram[1569]) );
  DFF ram_reg_1851__0_ ( .D(n5809), .CP(wclk), .Q(ram[1568]) );
  DFF ram_reg_1855__7_ ( .D(n5784), .CP(wclk), .Q(ram[1543]) );
  DFF ram_reg_1855__6_ ( .D(n5783), .CP(wclk), .Q(ram[1542]) );
  DFF ram_reg_1855__5_ ( .D(n5782), .CP(wclk), .Q(ram[1541]) );
  DFF ram_reg_1855__4_ ( .D(n5781), .CP(wclk), .Q(ram[1540]) );
  DFF ram_reg_1855__3_ ( .D(n5780), .CP(wclk), .Q(ram[1539]) );
  DFF ram_reg_1855__2_ ( .D(n5779), .CP(wclk), .Q(ram[1538]) );
  DFF ram_reg_1855__1_ ( .D(n5778), .CP(wclk), .Q(ram[1537]) );
  DFF ram_reg_1855__0_ ( .D(n5777), .CP(wclk), .Q(ram[1536]) );
  DFF ram_reg_1867__7_ ( .D(n5688), .CP(wclk), .Q(ram[1447]) );
  DFF ram_reg_1867__6_ ( .D(n5687), .CP(wclk), .Q(ram[1446]) );
  DFF ram_reg_1867__5_ ( .D(n5686), .CP(wclk), .Q(ram[1445]) );
  DFF ram_reg_1867__4_ ( .D(n5685), .CP(wclk), .Q(ram[1444]) );
  DFF ram_reg_1867__3_ ( .D(n5684), .CP(wclk), .Q(ram[1443]) );
  DFF ram_reg_1867__2_ ( .D(n5683), .CP(wclk), .Q(ram[1442]) );
  DFF ram_reg_1867__1_ ( .D(n5682), .CP(wclk), .Q(ram[1441]) );
  DFF ram_reg_1867__0_ ( .D(n5681), .CP(wclk), .Q(ram[1440]) );
  DFF ram_reg_1899__7_ ( .D(n5432), .CP(wclk), .Q(ram[1191]) );
  DFF ram_reg_1899__6_ ( .D(n5431), .CP(wclk), .Q(ram[1190]) );
  DFF ram_reg_1899__5_ ( .D(n5430), .CP(wclk), .Q(ram[1189]) );
  DFF ram_reg_1899__4_ ( .D(n5429), .CP(wclk), .Q(ram[1188]) );
  DFF ram_reg_1899__3_ ( .D(n5428), .CP(wclk), .Q(ram[1187]) );
  DFF ram_reg_1899__2_ ( .D(n5427), .CP(wclk), .Q(ram[1186]) );
  DFF ram_reg_1899__1_ ( .D(n5426), .CP(wclk), .Q(ram[1185]) );
  DFF ram_reg_1899__0_ ( .D(n5425), .CP(wclk), .Q(ram[1184]) );
  DFF ram_reg_1903__7_ ( .D(n5400), .CP(wclk), .Q(ram[1159]) );
  DFF ram_reg_1903__6_ ( .D(n5399), .CP(wclk), .Q(ram[1158]) );
  DFF ram_reg_1903__5_ ( .D(n5398), .CP(wclk), .Q(ram[1157]) );
  DFF ram_reg_1903__4_ ( .D(n5397), .CP(wclk), .Q(ram[1156]) );
  DFF ram_reg_1903__3_ ( .D(n5396), .CP(wclk), .Q(ram[1155]) );
  DFF ram_reg_1903__2_ ( .D(n5395), .CP(wclk), .Q(ram[1154]) );
  DFF ram_reg_1903__1_ ( .D(n5394), .CP(wclk), .Q(ram[1153]) );
  DFF ram_reg_1903__0_ ( .D(n5393), .CP(wclk), .Q(ram[1152]) );
  DFF ram_reg_1915__7_ ( .D(n5304), .CP(wclk), .Q(ram[1063]) );
  DFF ram_reg_1915__6_ ( .D(n5303), .CP(wclk), .Q(ram[1062]) );
  DFF ram_reg_1915__5_ ( .D(n5302), .CP(wclk), .Q(ram[1061]) );
  DFF ram_reg_1915__4_ ( .D(n5301), .CP(wclk), .Q(ram[1060]) );
  DFF ram_reg_1915__3_ ( .D(n5300), .CP(wclk), .Q(ram[1059]) );
  DFF ram_reg_1915__2_ ( .D(n5299), .CP(wclk), .Q(ram[1058]) );
  DFF ram_reg_1915__1_ ( .D(n5298), .CP(wclk), .Q(ram[1057]) );
  DFF ram_reg_1915__0_ ( .D(n5297), .CP(wclk), .Q(ram[1056]) );
  DFF ram_reg_1919__7_ ( .D(n5272), .CP(wclk), .Q(ram[1031]) );
  DFF ram_reg_1919__6_ ( .D(n5271), .CP(wclk), .Q(ram[1030]) );
  DFF ram_reg_1919__5_ ( .D(n5270), .CP(wclk), .Q(ram[1029]) );
  DFF ram_reg_1919__4_ ( .D(n5269), .CP(wclk), .Q(ram[1028]) );
  DFF ram_reg_1919__3_ ( .D(n5268), .CP(wclk), .Q(ram[1027]) );
  DFF ram_reg_1919__2_ ( .D(n5267), .CP(wclk), .Q(ram[1026]) );
  DFF ram_reg_1919__1_ ( .D(n5266), .CP(wclk), .Q(ram[1025]) );
  DFF ram_reg_1919__0_ ( .D(n5265), .CP(wclk), .Q(ram[1024]) );
  DFF ram_reg_1923__7_ ( .D(n5240), .CP(wclk), .Q(ram[999]) );
  DFF ram_reg_1923__6_ ( .D(n5239), .CP(wclk), .Q(ram[998]) );
  DFF ram_reg_1923__5_ ( .D(n5238), .CP(wclk), .Q(ram[997]) );
  DFF ram_reg_1923__4_ ( .D(n5237), .CP(wclk), .Q(ram[996]) );
  DFF ram_reg_1923__3_ ( .D(n5236), .CP(wclk), .Q(ram[995]) );
  DFF ram_reg_1923__2_ ( .D(n5235), .CP(wclk), .Q(ram[994]) );
  DFF ram_reg_1923__1_ ( .D(n5234), .CP(wclk), .Q(ram[993]) );
  DFF ram_reg_1923__0_ ( .D(n5233), .CP(wclk), .Q(ram[992]) );
  DFF ram_reg_1927__7_ ( .D(n5208), .CP(wclk), .Q(ram[967]) );
  DFF ram_reg_1927__6_ ( .D(n5207), .CP(wclk), .Q(ram[966]) );
  DFF ram_reg_1927__5_ ( .D(n5206), .CP(wclk), .Q(ram[965]) );
  DFF ram_reg_1927__4_ ( .D(n5205), .CP(wclk), .Q(ram[964]) );
  DFF ram_reg_1927__3_ ( .D(n5204), .CP(wclk), .Q(ram[963]) );
  DFF ram_reg_1927__2_ ( .D(n5203), .CP(wclk), .Q(ram[962]) );
  DFF ram_reg_1927__1_ ( .D(n5202), .CP(wclk), .Q(ram[961]) );
  DFF ram_reg_1927__0_ ( .D(n5201), .CP(wclk), .Q(ram[960]) );
  DFF ram_reg_1931__7_ ( .D(n5176), .CP(wclk), .Q(ram[935]) );
  DFF ram_reg_1931__6_ ( .D(n5175), .CP(wclk), .Q(ram[934]) );
  DFF ram_reg_1931__5_ ( .D(n5174), .CP(wclk), .Q(ram[933]) );
  DFF ram_reg_1931__4_ ( .D(n5173), .CP(wclk), .Q(ram[932]) );
  DFF ram_reg_1931__3_ ( .D(n5172), .CP(wclk), .Q(ram[931]) );
  DFF ram_reg_1931__2_ ( .D(n5171), .CP(wclk), .Q(ram[930]) );
  DFF ram_reg_1931__1_ ( .D(n5170), .CP(wclk), .Q(ram[929]) );
  DFF ram_reg_1931__0_ ( .D(n5169), .CP(wclk), .Q(ram[928]) );
  DFF ram_reg_1935__7_ ( .D(n5144), .CP(wclk), .Q(ram[903]) );
  DFF ram_reg_1935__6_ ( .D(n5143), .CP(wclk), .Q(ram[902]) );
  DFF ram_reg_1935__5_ ( .D(n5142), .CP(wclk), .Q(ram[901]) );
  DFF ram_reg_1935__4_ ( .D(n5141), .CP(wclk), .Q(ram[900]) );
  DFF ram_reg_1935__3_ ( .D(n5140), .CP(wclk), .Q(ram[899]) );
  DFF ram_reg_1935__2_ ( .D(n5139), .CP(wclk), .Q(ram[898]) );
  DFF ram_reg_1935__1_ ( .D(n5138), .CP(wclk), .Q(ram[897]) );
  DFF ram_reg_1935__0_ ( .D(n5137), .CP(wclk), .Q(ram[896]) );
  DFF ram_reg_1939__7_ ( .D(n5112), .CP(wclk), .Q(ram[871]) );
  DFF ram_reg_1939__6_ ( .D(n5111), .CP(wclk), .Q(ram[870]) );
  DFF ram_reg_1939__5_ ( .D(n5110), .CP(wclk), .Q(ram[869]) );
  DFF ram_reg_1939__4_ ( .D(n5109), .CP(wclk), .Q(ram[868]) );
  DFF ram_reg_1939__3_ ( .D(n5108), .CP(wclk), .Q(ram[867]) );
  DFF ram_reg_1939__2_ ( .D(n5107), .CP(wclk), .Q(ram[866]) );
  DFF ram_reg_1939__1_ ( .D(n5106), .CP(wclk), .Q(ram[865]) );
  DFF ram_reg_1939__0_ ( .D(n5105), .CP(wclk), .Q(ram[864]) );
  DFF ram_reg_1947__7_ ( .D(n5048), .CP(wclk), .Q(ram[807]) );
  DFF ram_reg_1947__6_ ( .D(n5047), .CP(wclk), .Q(ram[806]) );
  DFF ram_reg_1947__5_ ( .D(n5046), .CP(wclk), .Q(ram[805]) );
  DFF ram_reg_1947__4_ ( .D(n5045), .CP(wclk), .Q(ram[804]) );
  DFF ram_reg_1947__3_ ( .D(n5044), .CP(wclk), .Q(ram[803]) );
  DFF ram_reg_1947__2_ ( .D(n5043), .CP(wclk), .Q(ram[802]) );
  DFF ram_reg_1947__1_ ( .D(n5042), .CP(wclk), .Q(ram[801]) );
  DFF ram_reg_1947__0_ ( .D(n5041), .CP(wclk), .Q(ram[800]) );
  DFF ram_reg_1951__7_ ( .D(n5016), .CP(wclk), .Q(ram[775]) );
  DFF ram_reg_1951__6_ ( .D(n5015), .CP(wclk), .Q(ram[774]) );
  DFF ram_reg_1951__5_ ( .D(n5014), .CP(wclk), .Q(ram[773]) );
  DFF ram_reg_1951__4_ ( .D(n5013), .CP(wclk), .Q(ram[772]) );
  DFF ram_reg_1951__3_ ( .D(n5012), .CP(wclk), .Q(ram[771]) );
  DFF ram_reg_1951__2_ ( .D(n5011), .CP(wclk), .Q(ram[770]) );
  DFF ram_reg_1951__1_ ( .D(n5010), .CP(wclk), .Q(ram[769]) );
  DFF ram_reg_1951__0_ ( .D(n5009), .CP(wclk), .Q(ram[768]) );
  DFF ram_reg_1955__7_ ( .D(n4984), .CP(wclk), .Q(ram[743]) );
  DFF ram_reg_1955__6_ ( .D(n4983), .CP(wclk), .Q(ram[742]) );
  DFF ram_reg_1955__5_ ( .D(n4982), .CP(wclk), .Q(ram[741]) );
  DFF ram_reg_1955__4_ ( .D(n4981), .CP(wclk), .Q(ram[740]) );
  DFF ram_reg_1955__3_ ( .D(n4980), .CP(wclk), .Q(ram[739]) );
  DFF ram_reg_1955__2_ ( .D(n4979), .CP(wclk), .Q(ram[738]) );
  DFF ram_reg_1955__1_ ( .D(n4978), .CP(wclk), .Q(ram[737]) );
  DFF ram_reg_1955__0_ ( .D(n4977), .CP(wclk), .Q(ram[736]) );
  DFF ram_reg_1959__7_ ( .D(n4952), .CP(wclk), .Q(ram[711]) );
  DFF ram_reg_1959__6_ ( .D(n4951), .CP(wclk), .Q(ram[710]) );
  DFF ram_reg_1959__5_ ( .D(n4950), .CP(wclk), .Q(ram[709]) );
  DFF ram_reg_1959__4_ ( .D(n4949), .CP(wclk), .Q(ram[708]) );
  DFF ram_reg_1959__3_ ( .D(n4948), .CP(wclk), .Q(ram[707]) );
  DFF ram_reg_1959__2_ ( .D(n4947), .CP(wclk), .Q(ram[706]) );
  DFF ram_reg_1959__1_ ( .D(n4946), .CP(wclk), .Q(ram[705]) );
  DFF ram_reg_1959__0_ ( .D(n4945), .CP(wclk), .Q(ram[704]) );
  DFF ram_reg_1963__7_ ( .D(n4920), .CP(wclk), .Q(ram[679]) );
  DFF ram_reg_1963__6_ ( .D(n4919), .CP(wclk), .Q(ram[678]) );
  DFF ram_reg_1963__5_ ( .D(n4918), .CP(wclk), .Q(ram[677]) );
  DFF ram_reg_1963__4_ ( .D(n4917), .CP(wclk), .Q(ram[676]) );
  DFF ram_reg_1963__3_ ( .D(n4916), .CP(wclk), .Q(ram[675]) );
  DFF ram_reg_1963__2_ ( .D(n4915), .CP(wclk), .Q(ram[674]) );
  DFF ram_reg_1963__1_ ( .D(n4914), .CP(wclk), .Q(ram[673]) );
  DFF ram_reg_1963__0_ ( .D(n4913), .CP(wclk), .Q(ram[672]) );
  DFF ram_reg_1967__7_ ( .D(n4888), .CP(wclk), .Q(ram[647]) );
  DFF ram_reg_1967__6_ ( .D(n4887), .CP(wclk), .Q(ram[646]) );
  DFF ram_reg_1967__5_ ( .D(n4886), .CP(wclk), .Q(ram[645]) );
  DFF ram_reg_1967__4_ ( .D(n4885), .CP(wclk), .Q(ram[644]) );
  DFF ram_reg_1967__3_ ( .D(n4884), .CP(wclk), .Q(ram[643]) );
  DFF ram_reg_1967__2_ ( .D(n4883), .CP(wclk), .Q(ram[642]) );
  DFF ram_reg_1967__1_ ( .D(n4882), .CP(wclk), .Q(ram[641]) );
  DFF ram_reg_1967__0_ ( .D(n4881), .CP(wclk), .Q(ram[640]) );
  DFF ram_reg_1971__7_ ( .D(n4856), .CP(wclk), .Q(ram[615]) );
  DFF ram_reg_1971__6_ ( .D(n4855), .CP(wclk), .Q(ram[614]) );
  DFF ram_reg_1971__5_ ( .D(n4854), .CP(wclk), .Q(ram[613]) );
  DFF ram_reg_1971__4_ ( .D(n4853), .CP(wclk), .Q(ram[612]) );
  DFF ram_reg_1971__3_ ( .D(n4852), .CP(wclk), .Q(ram[611]) );
  DFF ram_reg_1971__2_ ( .D(n4851), .CP(wclk), .Q(ram[610]) );
  DFF ram_reg_1971__1_ ( .D(n4850), .CP(wclk), .Q(ram[609]) );
  DFF ram_reg_1971__0_ ( .D(n4849), .CP(wclk), .Q(ram[608]) );
  DFF ram_reg_1975__7_ ( .D(n4824), .CP(wclk), .Q(ram[583]) );
  DFF ram_reg_1975__6_ ( .D(n4823), .CP(wclk), .Q(ram[582]) );
  DFF ram_reg_1975__5_ ( .D(n4822), .CP(wclk), .Q(ram[581]) );
  DFF ram_reg_1975__4_ ( .D(n4821), .CP(wclk), .Q(ram[580]) );
  DFF ram_reg_1975__3_ ( .D(n4820), .CP(wclk), .Q(ram[579]) );
  DFF ram_reg_1975__2_ ( .D(n4819), .CP(wclk), .Q(ram[578]) );
  DFF ram_reg_1975__1_ ( .D(n4818), .CP(wclk), .Q(ram[577]) );
  DFF ram_reg_1975__0_ ( .D(n4817), .CP(wclk), .Q(ram[576]) );
  DFF ram_reg_1979__7_ ( .D(n4792), .CP(wclk), .Q(ram[551]) );
  DFF ram_reg_1979__6_ ( .D(n4791), .CP(wclk), .Q(ram[550]) );
  DFF ram_reg_1979__5_ ( .D(n4790), .CP(wclk), .Q(ram[549]) );
  DFF ram_reg_1979__4_ ( .D(n4789), .CP(wclk), .Q(ram[548]) );
  DFF ram_reg_1979__3_ ( .D(n4788), .CP(wclk), .Q(ram[547]) );
  DFF ram_reg_1979__2_ ( .D(n4787), .CP(wclk), .Q(ram[546]) );
  DFF ram_reg_1979__1_ ( .D(n4786), .CP(wclk), .Q(ram[545]) );
  DFF ram_reg_1979__0_ ( .D(n4785), .CP(wclk), .Q(ram[544]) );
  DFF ram_reg_1983__7_ ( .D(n4760), .CP(wclk), .Q(ram[519]) );
  DFF ram_reg_1983__6_ ( .D(n4759), .CP(wclk), .Q(ram[518]) );
  DFF ram_reg_1983__5_ ( .D(n4758), .CP(wclk), .Q(ram[517]) );
  DFF ram_reg_1983__4_ ( .D(n4757), .CP(wclk), .Q(ram[516]) );
  DFF ram_reg_1983__3_ ( .D(n4756), .CP(wclk), .Q(ram[515]) );
  DFF ram_reg_1983__2_ ( .D(n4755), .CP(wclk), .Q(ram[514]) );
  DFF ram_reg_1983__1_ ( .D(n4754), .CP(wclk), .Q(ram[513]) );
  DFF ram_reg_1983__0_ ( .D(n4753), .CP(wclk), .Q(ram[512]) );
  DFF ram_reg_1987__7_ ( .D(n4728), .CP(wclk), .Q(ram[487]) );
  DFF ram_reg_1987__6_ ( .D(n4727), .CP(wclk), .Q(ram[486]) );
  DFF ram_reg_1987__5_ ( .D(n4726), .CP(wclk), .Q(ram[485]) );
  DFF ram_reg_1987__4_ ( .D(n4725), .CP(wclk), .Q(ram[484]) );
  DFF ram_reg_1987__3_ ( .D(n4724), .CP(wclk), .Q(ram[483]) );
  DFF ram_reg_1987__2_ ( .D(n4723), .CP(wclk), .Q(ram[482]) );
  DFF ram_reg_1987__1_ ( .D(n4722), .CP(wclk), .Q(ram[481]) );
  DFF ram_reg_1987__0_ ( .D(n4721), .CP(wclk), .Q(ram[480]) );
  DFF ram_reg_1995__7_ ( .D(n4664), .CP(wclk), .Q(ram[423]) );
  DFF ram_reg_1995__6_ ( .D(n4663), .CP(wclk), .Q(ram[422]) );
  DFF ram_reg_1995__5_ ( .D(n4662), .CP(wclk), .Q(ram[421]) );
  DFF ram_reg_1995__4_ ( .D(n4661), .CP(wclk), .Q(ram[420]) );
  DFF ram_reg_1995__3_ ( .D(n4660), .CP(wclk), .Q(ram[419]) );
  DFF ram_reg_1995__2_ ( .D(n4659), .CP(wclk), .Q(ram[418]) );
  DFF ram_reg_1995__1_ ( .D(n4658), .CP(wclk), .Q(ram[417]) );
  DFF ram_reg_1995__0_ ( .D(n4657), .CP(wclk), .Q(ram[416]) );
  DFF ram_reg_1999__7_ ( .D(n4632), .CP(wclk), .Q(ram[391]) );
  DFF ram_reg_1999__6_ ( .D(n4631), .CP(wclk), .Q(ram[390]) );
  DFF ram_reg_1999__5_ ( .D(n4630), .CP(wclk), .Q(ram[389]) );
  DFF ram_reg_1999__4_ ( .D(n4629), .CP(wclk), .Q(ram[388]) );
  DFF ram_reg_1999__3_ ( .D(n4628), .CP(wclk), .Q(ram[387]) );
  DFF ram_reg_1999__2_ ( .D(n4627), .CP(wclk), .Q(ram[386]) );
  DFF ram_reg_1999__1_ ( .D(n4626), .CP(wclk), .Q(ram[385]) );
  DFF ram_reg_1999__0_ ( .D(n4625), .CP(wclk), .Q(ram[384]) );
  DFF ram_reg_2003__7_ ( .D(n4600), .CP(wclk), .Q(ram[359]) );
  DFF ram_reg_2003__6_ ( .D(n4599), .CP(wclk), .Q(ram[358]) );
  DFF ram_reg_2003__5_ ( .D(n4598), .CP(wclk), .Q(ram[357]) );
  DFF ram_reg_2003__4_ ( .D(n4597), .CP(wclk), .Q(ram[356]) );
  DFF ram_reg_2003__3_ ( .D(n4596), .CP(wclk), .Q(ram[355]) );
  DFF ram_reg_2003__2_ ( .D(n4595), .CP(wclk), .Q(ram[354]) );
  DFF ram_reg_2003__1_ ( .D(n4594), .CP(wclk), .Q(ram[353]) );
  DFF ram_reg_2003__0_ ( .D(n4593), .CP(wclk), .Q(ram[352]) );
  DFF ram_reg_2011__7_ ( .D(n4536), .CP(wclk), .Q(ram[295]) );
  DFF ram_reg_2011__6_ ( .D(n4535), .CP(wclk), .Q(ram[294]) );
  DFF ram_reg_2011__5_ ( .D(n4534), .CP(wclk), .Q(ram[293]) );
  DFF ram_reg_2011__4_ ( .D(n4533), .CP(wclk), .Q(ram[292]) );
  DFF ram_reg_2011__3_ ( .D(n4532), .CP(wclk), .Q(ram[291]) );
  DFF ram_reg_2011__2_ ( .D(n4531), .CP(wclk), .Q(ram[290]) );
  DFF ram_reg_2011__1_ ( .D(n4530), .CP(wclk), .Q(ram[289]) );
  DFF ram_reg_2011__0_ ( .D(n4529), .CP(wclk), .Q(ram[288]) );
  DFF ram_reg_2015__7_ ( .D(n4504), .CP(wclk), .Q(ram[263]) );
  DFF ram_reg_2015__6_ ( .D(n4503), .CP(wclk), .Q(ram[262]) );
  DFF ram_reg_2015__5_ ( .D(n4502), .CP(wclk), .Q(ram[261]) );
  DFF ram_reg_2015__4_ ( .D(n4501), .CP(wclk), .Q(ram[260]) );
  DFF ram_reg_2015__3_ ( .D(n4500), .CP(wclk), .Q(ram[259]) );
  DFF ram_reg_2015__2_ ( .D(n4499), .CP(wclk), .Q(ram[258]) );
  DFF ram_reg_2015__1_ ( .D(n4498), .CP(wclk), .Q(ram[257]) );
  DFF ram_reg_2015__0_ ( .D(n4497), .CP(wclk), .Q(ram[256]) );
  DFF ram_reg_2019__7_ ( .D(n4472), .CP(wclk), .Q(ram[231]) );
  DFF ram_reg_2019__6_ ( .D(n4471), .CP(wclk), .Q(ram[230]) );
  DFF ram_reg_2019__5_ ( .D(n4470), .CP(wclk), .Q(ram[229]) );
  DFF ram_reg_2019__4_ ( .D(n4469), .CP(wclk), .Q(ram[228]) );
  DFF ram_reg_2019__3_ ( .D(n4468), .CP(wclk), .Q(ram[227]) );
  DFF ram_reg_2019__2_ ( .D(n4467), .CP(wclk), .Q(ram[226]) );
  DFF ram_reg_2019__1_ ( .D(n4466), .CP(wclk), .Q(ram[225]) );
  DFF ram_reg_2019__0_ ( .D(n4465), .CP(wclk), .Q(ram[224]) );
  DFF ram_reg_2023__7_ ( .D(n4440), .CP(wclk), .Q(ram[199]) );
  DFF ram_reg_2023__6_ ( .D(n4439), .CP(wclk), .Q(ram[198]) );
  DFF ram_reg_2023__5_ ( .D(n4438), .CP(wclk), .Q(ram[197]) );
  DFF ram_reg_2023__4_ ( .D(n4437), .CP(wclk), .Q(ram[196]) );
  DFF ram_reg_2023__3_ ( .D(n4436), .CP(wclk), .Q(ram[195]) );
  DFF ram_reg_2023__2_ ( .D(n4435), .CP(wclk), .Q(ram[194]) );
  DFF ram_reg_2023__1_ ( .D(n4434), .CP(wclk), .Q(ram[193]) );
  DFF ram_reg_2023__0_ ( .D(n4433), .CP(wclk), .Q(ram[192]) );
  DFF ram_reg_2027__7_ ( .D(n4408), .CP(wclk), .Q(ram[167]) );
  DFF ram_reg_2027__6_ ( .D(n4407), .CP(wclk), .Q(ram[166]) );
  DFF ram_reg_2027__5_ ( .D(n4406), .CP(wclk), .Q(ram[165]) );
  DFF ram_reg_2027__4_ ( .D(n4405), .CP(wclk), .Q(ram[164]) );
  DFF ram_reg_2027__3_ ( .D(n4404), .CP(wclk), .Q(ram[163]) );
  DFF ram_reg_2027__2_ ( .D(n4403), .CP(wclk), .Q(ram[162]) );
  DFF ram_reg_2027__1_ ( .D(n4402), .CP(wclk), .Q(ram[161]) );
  DFF ram_reg_2027__0_ ( .D(n4401), .CP(wclk), .Q(ram[160]) );
  DFF ram_reg_2031__7_ ( .D(n4376), .CP(wclk), .Q(ram[135]) );
  DFF ram_reg_2031__6_ ( .D(n4375), .CP(wclk), .Q(ram[134]) );
  DFF ram_reg_2031__5_ ( .D(n4374), .CP(wclk), .Q(ram[133]) );
  DFF ram_reg_2031__4_ ( .D(n4373), .CP(wclk), .Q(ram[132]) );
  DFF ram_reg_2031__3_ ( .D(n4372), .CP(wclk), .Q(ram[131]) );
  DFF ram_reg_2031__2_ ( .D(n4371), .CP(wclk), .Q(ram[130]) );
  DFF ram_reg_2031__1_ ( .D(n4370), .CP(wclk), .Q(ram[129]) );
  DFF ram_reg_2031__0_ ( .D(n4369), .CP(wclk), .Q(ram[128]) );
  DFF ram_reg_2035__7_ ( .D(n4344), .CP(wclk), .Q(ram[103]) );
  DFF ram_reg_2035__6_ ( .D(n4343), .CP(wclk), .Q(ram[102]) );
  DFF ram_reg_2035__5_ ( .D(n4342), .CP(wclk), .Q(ram[101]) );
  DFF ram_reg_2035__4_ ( .D(n4341), .CP(wclk), .Q(ram[100]) );
  DFF ram_reg_2035__3_ ( .D(n4340), .CP(wclk), .Q(ram[99]) );
  DFF ram_reg_2035__2_ ( .D(n4339), .CP(wclk), .Q(ram[98]) );
  DFF ram_reg_2035__1_ ( .D(n4338), .CP(wclk), .Q(ram[97]) );
  DFF ram_reg_2035__0_ ( .D(n4337), .CP(wclk), .Q(ram[96]) );
  DFF ram_reg_2039__7_ ( .D(n4312), .CP(wclk), .Q(ram[71]) );
  DFF ram_reg_2039__6_ ( .D(n4311), .CP(wclk), .Q(ram[70]) );
  DFF ram_reg_2039__5_ ( .D(n4310), .CP(wclk), .Q(ram[69]) );
  DFF ram_reg_2039__4_ ( .D(n4309), .CP(wclk), .Q(ram[68]) );
  DFF ram_reg_2039__3_ ( .D(n4308), .CP(wclk), .Q(ram[67]) );
  DFF ram_reg_2039__2_ ( .D(n4307), .CP(wclk), .Q(ram[66]) );
  DFF ram_reg_2039__1_ ( .D(n4306), .CP(wclk), .Q(ram[65]) );
  DFF ram_reg_2039__0_ ( .D(n4305), .CP(wclk), .Q(ram[64]) );
  DFF ram_reg_2043__7_ ( .D(n4280), .CP(wclk), .Q(ram[39]) );
  DFF ram_reg_2043__6_ ( .D(n4279), .CP(wclk), .Q(ram[38]) );
  DFF ram_reg_2043__5_ ( .D(n4278), .CP(wclk), .Q(ram[37]) );
  DFF ram_reg_2043__4_ ( .D(n4277), .CP(wclk), .Q(ram[36]) );
  DFF ram_reg_2043__3_ ( .D(n4276), .CP(wclk), .Q(ram[35]) );
  DFF ram_reg_2043__2_ ( .D(n4275), .CP(wclk), .Q(ram[34]) );
  DFF ram_reg_2043__1_ ( .D(n4274), .CP(wclk), .Q(ram[33]) );
  DFF ram_reg_2043__0_ ( .D(n4273), .CP(wclk), .Q(ram[32]) );
  DFF ram_reg_2047__7_ ( .D(n4248), .CP(wclk), .Q(ram[7]) );
  DFF ram_reg_2047__6_ ( .D(n4247), .CP(wclk), .Q(ram[6]) );
  DFF ram_reg_2047__5_ ( .D(n4246), .CP(wclk), .Q(ram[5]) );
  DFF ram_reg_2047__4_ ( .D(n4245), .CP(wclk), .Q(ram[4]) );
  DFF ram_reg_2047__3_ ( .D(n4244), .CP(wclk), .Q(ram[3]) );
  DFF ram_reg_2047__2_ ( .D(n4243), .CP(wclk), .Q(ram[2]) );
  DFF ram_reg_2047__1_ ( .D(n4242), .CP(wclk), .Q(ram[1]) );
  DFF ram_reg_2047__0_ ( .D(n4241), .CP(wclk), .Q(ram[0]) );
  DFF ram_reg_0__7_ ( .D(n20624), .CP(wclk), .Q(ram[16383]) );
  DFF ram_reg_0__6_ ( .D(n20623), .CP(wclk), .Q(ram[16382]) );
  DFF ram_reg_0__5_ ( .D(n20622), .CP(wclk), .Q(ram[16381]) );
  DFF ram_reg_0__4_ ( .D(n20621), .CP(wclk), .Q(ram[16380]) );
  DFF ram_reg_0__3_ ( .D(n20620), .CP(wclk), .Q(ram[16379]) );
  DFF ram_reg_0__2_ ( .D(n20619), .CP(wclk), .Q(ram[16378]) );
  DFF ram_reg_0__1_ ( .D(n20618), .CP(wclk), .Q(ram[16377]) );
  DFF ram_reg_0__0_ ( .D(n20617), .CP(wclk), .Q(ram[16376]) );
  DFF ram_reg_4__7_ ( .D(n20592), .CP(wclk), .Q(ram[16351]) );
  DFF ram_reg_4__6_ ( .D(n20591), .CP(wclk), .Q(ram[16350]) );
  DFF ram_reg_4__5_ ( .D(n20590), .CP(wclk), .Q(ram[16349]) );
  DFF ram_reg_4__4_ ( .D(n20589), .CP(wclk), .Q(ram[16348]) );
  DFF ram_reg_4__3_ ( .D(n20588), .CP(wclk), .Q(ram[16347]) );
  DFF ram_reg_4__2_ ( .D(n20587), .CP(wclk), .Q(ram[16346]) );
  DFF ram_reg_4__1_ ( .D(n20586), .CP(wclk), .Q(ram[16345]) );
  DFF ram_reg_4__0_ ( .D(n20585), .CP(wclk), .Q(ram[16344]) );
  DFF ram_reg_8__7_ ( .D(n20560), .CP(wclk), .Q(ram[16319]) );
  DFF ram_reg_8__6_ ( .D(n20559), .CP(wclk), .Q(ram[16318]) );
  DFF ram_reg_8__5_ ( .D(n20558), .CP(wclk), .Q(ram[16317]) );
  DFF ram_reg_8__4_ ( .D(n20557), .CP(wclk), .Q(ram[16316]) );
  DFF ram_reg_8__3_ ( .D(n20556), .CP(wclk), .Q(ram[16315]) );
  DFF ram_reg_8__2_ ( .D(n20555), .CP(wclk), .Q(ram[16314]) );
  DFF ram_reg_8__1_ ( .D(n20554), .CP(wclk), .Q(ram[16313]) );
  DFF ram_reg_8__0_ ( .D(n20553), .CP(wclk), .Q(ram[16312]) );
  DFF ram_reg_12__7_ ( .D(n20528), .CP(wclk), .Q(ram[16287]) );
  DFF ram_reg_12__6_ ( .D(n20527), .CP(wclk), .Q(ram[16286]) );
  DFF ram_reg_12__5_ ( .D(n20526), .CP(wclk), .Q(ram[16285]) );
  DFF ram_reg_12__4_ ( .D(n20525), .CP(wclk), .Q(ram[16284]) );
  DFF ram_reg_12__3_ ( .D(n20524), .CP(wclk), .Q(ram[16283]) );
  DFF ram_reg_12__2_ ( .D(n20523), .CP(wclk), .Q(ram[16282]) );
  DFF ram_reg_12__1_ ( .D(n20522), .CP(wclk), .Q(ram[16281]) );
  DFF ram_reg_12__0_ ( .D(n20521), .CP(wclk), .Q(ram[16280]) );
  DFF ram_reg_16__7_ ( .D(n20496), .CP(wclk), .Q(ram[16255]) );
  DFF ram_reg_16__6_ ( .D(n20495), .CP(wclk), .Q(ram[16254]) );
  DFF ram_reg_16__5_ ( .D(n20494), .CP(wclk), .Q(ram[16253]) );
  DFF ram_reg_16__4_ ( .D(n20493), .CP(wclk), .Q(ram[16252]) );
  DFF ram_reg_16__3_ ( .D(n20492), .CP(wclk), .Q(ram[16251]) );
  DFF ram_reg_16__2_ ( .D(n20491), .CP(wclk), .Q(ram[16250]) );
  DFF ram_reg_16__1_ ( .D(n20490), .CP(wclk), .Q(ram[16249]) );
  DFF ram_reg_16__0_ ( .D(n20489), .CP(wclk), .Q(ram[16248]) );
  DFF ram_reg_20__7_ ( .D(n20464), .CP(wclk), .Q(ram[16223]) );
  DFF ram_reg_20__6_ ( .D(n20463), .CP(wclk), .Q(ram[16222]) );
  DFF ram_reg_20__5_ ( .D(n20462), .CP(wclk), .Q(ram[16221]) );
  DFF ram_reg_20__4_ ( .D(n20461), .CP(wclk), .Q(ram[16220]) );
  DFF ram_reg_20__3_ ( .D(n20460), .CP(wclk), .Q(ram[16219]) );
  DFF ram_reg_20__2_ ( .D(n20459), .CP(wclk), .Q(ram[16218]) );
  DFF ram_reg_20__1_ ( .D(n20458), .CP(wclk), .Q(ram[16217]) );
  DFF ram_reg_20__0_ ( .D(n20457), .CP(wclk), .Q(ram[16216]) );
  DFF ram_reg_24__7_ ( .D(n20432), .CP(wclk), .Q(ram[16191]) );
  DFF ram_reg_24__6_ ( .D(n20431), .CP(wclk), .Q(ram[16190]) );
  DFF ram_reg_24__5_ ( .D(n20430), .CP(wclk), .Q(ram[16189]) );
  DFF ram_reg_24__4_ ( .D(n20429), .CP(wclk), .Q(ram[16188]) );
  DFF ram_reg_24__3_ ( .D(n20428), .CP(wclk), .Q(ram[16187]) );
  DFF ram_reg_24__2_ ( .D(n20427), .CP(wclk), .Q(ram[16186]) );
  DFF ram_reg_24__1_ ( .D(n20426), .CP(wclk), .Q(ram[16185]) );
  DFF ram_reg_24__0_ ( .D(n20425), .CP(wclk), .Q(ram[16184]) );
  DFF ram_reg_28__7_ ( .D(n20400), .CP(wclk), .Q(ram[16159]) );
  DFF ram_reg_28__6_ ( .D(n20399), .CP(wclk), .Q(ram[16158]) );
  DFF ram_reg_28__5_ ( .D(n20398), .CP(wclk), .Q(ram[16157]) );
  DFF ram_reg_28__4_ ( .D(n20397), .CP(wclk), .Q(ram[16156]) );
  DFF ram_reg_28__3_ ( .D(n20396), .CP(wclk), .Q(ram[16155]) );
  DFF ram_reg_28__2_ ( .D(n20395), .CP(wclk), .Q(ram[16154]) );
  DFF ram_reg_28__1_ ( .D(n20394), .CP(wclk), .Q(ram[16153]) );
  DFF ram_reg_28__0_ ( .D(n20393), .CP(wclk), .Q(ram[16152]) );
  DFF ram_reg_32__7_ ( .D(n20368), .CP(wclk), .Q(ram[16127]) );
  DFF ram_reg_32__6_ ( .D(n20367), .CP(wclk), .Q(ram[16126]) );
  DFF ram_reg_32__5_ ( .D(n20366), .CP(wclk), .Q(ram[16125]) );
  DFF ram_reg_32__4_ ( .D(n20365), .CP(wclk), .Q(ram[16124]) );
  DFF ram_reg_32__3_ ( .D(n20364), .CP(wclk), .Q(ram[16123]) );
  DFF ram_reg_32__2_ ( .D(n20363), .CP(wclk), .Q(ram[16122]) );
  DFF ram_reg_32__1_ ( .D(n20362), .CP(wclk), .Q(ram[16121]) );
  DFF ram_reg_32__0_ ( .D(n20361), .CP(wclk), .Q(ram[16120]) );
  DFF ram_reg_36__7_ ( .D(n20336), .CP(wclk), .Q(ram[16095]) );
  DFF ram_reg_36__6_ ( .D(n20335), .CP(wclk), .Q(ram[16094]) );
  DFF ram_reg_36__5_ ( .D(n20334), .CP(wclk), .Q(ram[16093]) );
  DFF ram_reg_36__4_ ( .D(n20333), .CP(wclk), .Q(ram[16092]) );
  DFF ram_reg_36__3_ ( .D(n20332), .CP(wclk), .Q(ram[16091]) );
  DFF ram_reg_36__2_ ( .D(n20331), .CP(wclk), .Q(ram[16090]) );
  DFF ram_reg_36__1_ ( .D(n20330), .CP(wclk), .Q(ram[16089]) );
  DFF ram_reg_36__0_ ( .D(n20329), .CP(wclk), .Q(ram[16088]) );
  DFF ram_reg_44__7_ ( .D(n20272), .CP(wclk), .Q(ram[16031]) );
  DFF ram_reg_44__6_ ( .D(n20271), .CP(wclk), .Q(ram[16030]) );
  DFF ram_reg_44__5_ ( .D(n20270), .CP(wclk), .Q(ram[16029]) );
  DFF ram_reg_44__4_ ( .D(n20269), .CP(wclk), .Q(ram[16028]) );
  DFF ram_reg_44__3_ ( .D(n20268), .CP(wclk), .Q(ram[16027]) );
  DFF ram_reg_44__2_ ( .D(n20267), .CP(wclk), .Q(ram[16026]) );
  DFF ram_reg_44__1_ ( .D(n20266), .CP(wclk), .Q(ram[16025]) );
  DFF ram_reg_44__0_ ( .D(n20265), .CP(wclk), .Q(ram[16024]) );
  DFF ram_reg_48__7_ ( .D(n20240), .CP(wclk), .Q(ram[15999]) );
  DFF ram_reg_48__6_ ( .D(n20239), .CP(wclk), .Q(ram[15998]) );
  DFF ram_reg_48__5_ ( .D(n20238), .CP(wclk), .Q(ram[15997]) );
  DFF ram_reg_48__4_ ( .D(n20237), .CP(wclk), .Q(ram[15996]) );
  DFF ram_reg_48__3_ ( .D(n20236), .CP(wclk), .Q(ram[15995]) );
  DFF ram_reg_48__2_ ( .D(n20235), .CP(wclk), .Q(ram[15994]) );
  DFF ram_reg_48__1_ ( .D(n20234), .CP(wclk), .Q(ram[15993]) );
  DFF ram_reg_48__0_ ( .D(n20233), .CP(wclk), .Q(ram[15992]) );
  DFF ram_reg_52__7_ ( .D(n20208), .CP(wclk), .Q(ram[15967]) );
  DFF ram_reg_52__6_ ( .D(n20207), .CP(wclk), .Q(ram[15966]) );
  DFF ram_reg_52__5_ ( .D(n20206), .CP(wclk), .Q(ram[15965]) );
  DFF ram_reg_52__4_ ( .D(n20205), .CP(wclk), .Q(ram[15964]) );
  DFF ram_reg_52__3_ ( .D(n20204), .CP(wclk), .Q(ram[15963]) );
  DFF ram_reg_52__2_ ( .D(n20203), .CP(wclk), .Q(ram[15962]) );
  DFF ram_reg_52__1_ ( .D(n20202), .CP(wclk), .Q(ram[15961]) );
  DFF ram_reg_52__0_ ( .D(n20201), .CP(wclk), .Q(ram[15960]) );
  DFF ram_reg_60__7_ ( .D(n20144), .CP(wclk), .Q(ram[15903]) );
  DFF ram_reg_60__6_ ( .D(n20143), .CP(wclk), .Q(ram[15902]) );
  DFF ram_reg_60__5_ ( .D(n20142), .CP(wclk), .Q(ram[15901]) );
  DFF ram_reg_60__4_ ( .D(n20141), .CP(wclk), .Q(ram[15900]) );
  DFF ram_reg_60__3_ ( .D(n20140), .CP(wclk), .Q(ram[15899]) );
  DFF ram_reg_60__2_ ( .D(n20139), .CP(wclk), .Q(ram[15898]) );
  DFF ram_reg_60__1_ ( .D(n20138), .CP(wclk), .Q(ram[15897]) );
  DFF ram_reg_60__0_ ( .D(n20137), .CP(wclk), .Q(ram[15896]) );
  DFF ram_reg_64__7_ ( .D(n20112), .CP(wclk), .Q(ram[15871]) );
  DFF ram_reg_64__6_ ( .D(n20111), .CP(wclk), .Q(ram[15870]) );
  DFF ram_reg_64__5_ ( .D(n20110), .CP(wclk), .Q(ram[15869]) );
  DFF ram_reg_64__4_ ( .D(n20109), .CP(wclk), .Q(ram[15868]) );
  DFF ram_reg_64__3_ ( .D(n20108), .CP(wclk), .Q(ram[15867]) );
  DFF ram_reg_64__2_ ( .D(n20107), .CP(wclk), .Q(ram[15866]) );
  DFF ram_reg_64__1_ ( .D(n20106), .CP(wclk), .Q(ram[15865]) );
  DFF ram_reg_64__0_ ( .D(n20105), .CP(wclk), .Q(ram[15864]) );
  DFF ram_reg_68__7_ ( .D(n20080), .CP(wclk), .Q(ram[15839]) );
  DFF ram_reg_68__6_ ( .D(n20079), .CP(wclk), .Q(ram[15838]) );
  DFF ram_reg_68__5_ ( .D(n20078), .CP(wclk), .Q(ram[15837]) );
  DFF ram_reg_68__4_ ( .D(n20077), .CP(wclk), .Q(ram[15836]) );
  DFF ram_reg_68__3_ ( .D(n20076), .CP(wclk), .Q(ram[15835]) );
  DFF ram_reg_68__2_ ( .D(n20075), .CP(wclk), .Q(ram[15834]) );
  DFF ram_reg_68__1_ ( .D(n20074), .CP(wclk), .Q(ram[15833]) );
  DFF ram_reg_68__0_ ( .D(n20073), .CP(wclk), .Q(ram[15832]) );
  DFF ram_reg_72__7_ ( .D(n20048), .CP(wclk), .Q(ram[15807]) );
  DFF ram_reg_72__6_ ( .D(n20047), .CP(wclk), .Q(ram[15806]) );
  DFF ram_reg_72__5_ ( .D(n20046), .CP(wclk), .Q(ram[15805]) );
  DFF ram_reg_72__4_ ( .D(n20045), .CP(wclk), .Q(ram[15804]) );
  DFF ram_reg_72__3_ ( .D(n20044), .CP(wclk), .Q(ram[15803]) );
  DFF ram_reg_72__2_ ( .D(n20043), .CP(wclk), .Q(ram[15802]) );
  DFF ram_reg_72__1_ ( .D(n20042), .CP(wclk), .Q(ram[15801]) );
  DFF ram_reg_72__0_ ( .D(n20041), .CP(wclk), .Q(ram[15800]) );
  DFF ram_reg_76__7_ ( .D(n20016), .CP(wclk), .Q(ram[15775]) );
  DFF ram_reg_76__6_ ( .D(n20015), .CP(wclk), .Q(ram[15774]) );
  DFF ram_reg_76__5_ ( .D(n20014), .CP(wclk), .Q(ram[15773]) );
  DFF ram_reg_76__4_ ( .D(n20013), .CP(wclk), .Q(ram[15772]) );
  DFF ram_reg_76__3_ ( .D(n20012), .CP(wclk), .Q(ram[15771]) );
  DFF ram_reg_76__2_ ( .D(n20011), .CP(wclk), .Q(ram[15770]) );
  DFF ram_reg_76__1_ ( .D(n20010), .CP(wclk), .Q(ram[15769]) );
  DFF ram_reg_76__0_ ( .D(n20009), .CP(wclk), .Q(ram[15768]) );
  DFF ram_reg_80__7_ ( .D(n19984), .CP(wclk), .Q(ram[15743]) );
  DFF ram_reg_80__6_ ( .D(n19983), .CP(wclk), .Q(ram[15742]) );
  DFF ram_reg_80__5_ ( .D(n19982), .CP(wclk), .Q(ram[15741]) );
  DFF ram_reg_80__4_ ( .D(n19981), .CP(wclk), .Q(ram[15740]) );
  DFF ram_reg_80__3_ ( .D(n19980), .CP(wclk), .Q(ram[15739]) );
  DFF ram_reg_80__2_ ( .D(n19979), .CP(wclk), .Q(ram[15738]) );
  DFF ram_reg_80__1_ ( .D(n19978), .CP(wclk), .Q(ram[15737]) );
  DFF ram_reg_80__0_ ( .D(n19977), .CP(wclk), .Q(ram[15736]) );
  DFF ram_reg_84__7_ ( .D(n19952), .CP(wclk), .Q(ram[15711]) );
  DFF ram_reg_84__6_ ( .D(n19951), .CP(wclk), .Q(ram[15710]) );
  DFF ram_reg_84__5_ ( .D(n19950), .CP(wclk), .Q(ram[15709]) );
  DFF ram_reg_84__4_ ( .D(n19949), .CP(wclk), .Q(ram[15708]) );
  DFF ram_reg_84__3_ ( .D(n19948), .CP(wclk), .Q(ram[15707]) );
  DFF ram_reg_84__2_ ( .D(n19947), .CP(wclk), .Q(ram[15706]) );
  DFF ram_reg_84__1_ ( .D(n19946), .CP(wclk), .Q(ram[15705]) );
  DFF ram_reg_84__0_ ( .D(n19945), .CP(wclk), .Q(ram[15704]) );
  DFF ram_reg_88__7_ ( .D(n19920), .CP(wclk), .Q(ram[15679]) );
  DFF ram_reg_88__6_ ( .D(n19919), .CP(wclk), .Q(ram[15678]) );
  DFF ram_reg_88__5_ ( .D(n19918), .CP(wclk), .Q(ram[15677]) );
  DFF ram_reg_88__4_ ( .D(n19917), .CP(wclk), .Q(ram[15676]) );
  DFF ram_reg_88__3_ ( .D(n19916), .CP(wclk), .Q(ram[15675]) );
  DFF ram_reg_88__2_ ( .D(n19915), .CP(wclk), .Q(ram[15674]) );
  DFF ram_reg_88__1_ ( .D(n19914), .CP(wclk), .Q(ram[15673]) );
  DFF ram_reg_88__0_ ( .D(n19913), .CP(wclk), .Q(ram[15672]) );
  DFF ram_reg_92__7_ ( .D(n19888), .CP(wclk), .Q(ram[15647]) );
  DFF ram_reg_92__6_ ( .D(n19887), .CP(wclk), .Q(ram[15646]) );
  DFF ram_reg_92__5_ ( .D(n19886), .CP(wclk), .Q(ram[15645]) );
  DFF ram_reg_92__4_ ( .D(n19885), .CP(wclk), .Q(ram[15644]) );
  DFF ram_reg_92__3_ ( .D(n19884), .CP(wclk), .Q(ram[15643]) );
  DFF ram_reg_92__2_ ( .D(n19883), .CP(wclk), .Q(ram[15642]) );
  DFF ram_reg_92__1_ ( .D(n19882), .CP(wclk), .Q(ram[15641]) );
  DFF ram_reg_92__0_ ( .D(n19881), .CP(wclk), .Q(ram[15640]) );
  DFF ram_reg_96__7_ ( .D(n19856), .CP(wclk), .Q(ram[15615]) );
  DFF ram_reg_96__6_ ( .D(n19855), .CP(wclk), .Q(ram[15614]) );
  DFF ram_reg_96__5_ ( .D(n19854), .CP(wclk), .Q(ram[15613]) );
  DFF ram_reg_96__4_ ( .D(n19853), .CP(wclk), .Q(ram[15612]) );
  DFF ram_reg_96__3_ ( .D(n19852), .CP(wclk), .Q(ram[15611]) );
  DFF ram_reg_96__2_ ( .D(n19851), .CP(wclk), .Q(ram[15610]) );
  DFF ram_reg_96__1_ ( .D(n19850), .CP(wclk), .Q(ram[15609]) );
  DFF ram_reg_96__0_ ( .D(n19849), .CP(wclk), .Q(ram[15608]) );
  DFF ram_reg_100__7_ ( .D(n19824), .CP(wclk), .Q(ram[15583]) );
  DFF ram_reg_100__6_ ( .D(n19823), .CP(wclk), .Q(ram[15582]) );
  DFF ram_reg_100__5_ ( .D(n19822), .CP(wclk), .Q(ram[15581]) );
  DFF ram_reg_100__4_ ( .D(n19821), .CP(wclk), .Q(ram[15580]) );
  DFF ram_reg_100__3_ ( .D(n19820), .CP(wclk), .Q(ram[15579]) );
  DFF ram_reg_100__2_ ( .D(n19819), .CP(wclk), .Q(ram[15578]) );
  DFF ram_reg_100__1_ ( .D(n19818), .CP(wclk), .Q(ram[15577]) );
  DFF ram_reg_100__0_ ( .D(n19817), .CP(wclk), .Q(ram[15576]) );
  DFF ram_reg_104__7_ ( .D(n19792), .CP(wclk), .Q(ram[15551]) );
  DFF ram_reg_104__6_ ( .D(n19791), .CP(wclk), .Q(ram[15550]) );
  DFF ram_reg_104__5_ ( .D(n19790), .CP(wclk), .Q(ram[15549]) );
  DFF ram_reg_104__4_ ( .D(n19789), .CP(wclk), .Q(ram[15548]) );
  DFF ram_reg_104__3_ ( .D(n19788), .CP(wclk), .Q(ram[15547]) );
  DFF ram_reg_104__2_ ( .D(n19787), .CP(wclk), .Q(ram[15546]) );
  DFF ram_reg_104__1_ ( .D(n19786), .CP(wclk), .Q(ram[15545]) );
  DFF ram_reg_104__0_ ( .D(n19785), .CP(wclk), .Q(ram[15544]) );
  DFF ram_reg_108__7_ ( .D(n19760), .CP(wclk), .Q(ram[15519]) );
  DFF ram_reg_108__6_ ( .D(n19759), .CP(wclk), .Q(ram[15518]) );
  DFF ram_reg_108__5_ ( .D(n19758), .CP(wclk), .Q(ram[15517]) );
  DFF ram_reg_108__4_ ( .D(n19757), .CP(wclk), .Q(ram[15516]) );
  DFF ram_reg_108__3_ ( .D(n19756), .CP(wclk), .Q(ram[15515]) );
  DFF ram_reg_108__2_ ( .D(n19755), .CP(wclk), .Q(ram[15514]) );
  DFF ram_reg_108__1_ ( .D(n19754), .CP(wclk), .Q(ram[15513]) );
  DFF ram_reg_108__0_ ( .D(n19753), .CP(wclk), .Q(ram[15512]) );
  DFF ram_reg_112__7_ ( .D(n19728), .CP(wclk), .Q(ram[15487]) );
  DFF ram_reg_112__6_ ( .D(n19727), .CP(wclk), .Q(ram[15486]) );
  DFF ram_reg_112__5_ ( .D(n19726), .CP(wclk), .Q(ram[15485]) );
  DFF ram_reg_112__4_ ( .D(n19725), .CP(wclk), .Q(ram[15484]) );
  DFF ram_reg_112__3_ ( .D(n19724), .CP(wclk), .Q(ram[15483]) );
  DFF ram_reg_112__2_ ( .D(n19723), .CP(wclk), .Q(ram[15482]) );
  DFF ram_reg_112__1_ ( .D(n19722), .CP(wclk), .Q(ram[15481]) );
  DFF ram_reg_112__0_ ( .D(n19721), .CP(wclk), .Q(ram[15480]) );
  DFF ram_reg_116__7_ ( .D(n19696), .CP(wclk), .Q(ram[15455]) );
  DFF ram_reg_116__6_ ( .D(n19695), .CP(wclk), .Q(ram[15454]) );
  DFF ram_reg_116__5_ ( .D(n19694), .CP(wclk), .Q(ram[15453]) );
  DFF ram_reg_116__4_ ( .D(n19693), .CP(wclk), .Q(ram[15452]) );
  DFF ram_reg_116__3_ ( .D(n19692), .CP(wclk), .Q(ram[15451]) );
  DFF ram_reg_116__2_ ( .D(n19691), .CP(wclk), .Q(ram[15450]) );
  DFF ram_reg_116__1_ ( .D(n19690), .CP(wclk), .Q(ram[15449]) );
  DFF ram_reg_116__0_ ( .D(n19689), .CP(wclk), .Q(ram[15448]) );
  DFF ram_reg_120__7_ ( .D(n19664), .CP(wclk), .Q(ram[15423]) );
  DFF ram_reg_120__6_ ( .D(n19663), .CP(wclk), .Q(ram[15422]) );
  DFF ram_reg_120__5_ ( .D(n19662), .CP(wclk), .Q(ram[15421]) );
  DFF ram_reg_120__4_ ( .D(n19661), .CP(wclk), .Q(ram[15420]) );
  DFF ram_reg_120__3_ ( .D(n19660), .CP(wclk), .Q(ram[15419]) );
  DFF ram_reg_120__2_ ( .D(n19659), .CP(wclk), .Q(ram[15418]) );
  DFF ram_reg_120__1_ ( .D(n19658), .CP(wclk), .Q(ram[15417]) );
  DFF ram_reg_120__0_ ( .D(n19657), .CP(wclk), .Q(ram[15416]) );
  DFF ram_reg_124__7_ ( .D(n19632), .CP(wclk), .Q(ram[15391]) );
  DFF ram_reg_124__6_ ( .D(n19631), .CP(wclk), .Q(ram[15390]) );
  DFF ram_reg_124__5_ ( .D(n19630), .CP(wclk), .Q(ram[15389]) );
  DFF ram_reg_124__4_ ( .D(n19629), .CP(wclk), .Q(ram[15388]) );
  DFF ram_reg_124__3_ ( .D(n19628), .CP(wclk), .Q(ram[15387]) );
  DFF ram_reg_124__2_ ( .D(n19627), .CP(wclk), .Q(ram[15386]) );
  DFF ram_reg_124__1_ ( .D(n19626), .CP(wclk), .Q(ram[15385]) );
  DFF ram_reg_124__0_ ( .D(n19625), .CP(wclk), .Q(ram[15384]) );
  DFF ram_reg_128__7_ ( .D(n19600), .CP(wclk), .Q(ram[15359]) );
  DFF ram_reg_128__6_ ( .D(n19599), .CP(wclk), .Q(ram[15358]) );
  DFF ram_reg_128__5_ ( .D(n19598), .CP(wclk), .Q(ram[15357]) );
  DFF ram_reg_128__4_ ( .D(n19597), .CP(wclk), .Q(ram[15356]) );
  DFF ram_reg_128__3_ ( .D(n19596), .CP(wclk), .Q(ram[15355]) );
  DFF ram_reg_128__2_ ( .D(n19595), .CP(wclk), .Q(ram[15354]) );
  DFF ram_reg_128__1_ ( .D(n19594), .CP(wclk), .Q(ram[15353]) );
  DFF ram_reg_128__0_ ( .D(n19593), .CP(wclk), .Q(ram[15352]) );
  DFF ram_reg_132__7_ ( .D(n19568), .CP(wclk), .Q(ram[15327]) );
  DFF ram_reg_132__6_ ( .D(n19567), .CP(wclk), .Q(ram[15326]) );
  DFF ram_reg_132__5_ ( .D(n19566), .CP(wclk), .Q(ram[15325]) );
  DFF ram_reg_132__4_ ( .D(n19565), .CP(wclk), .Q(ram[15324]) );
  DFF ram_reg_132__3_ ( .D(n19564), .CP(wclk), .Q(ram[15323]) );
  DFF ram_reg_132__2_ ( .D(n19563), .CP(wclk), .Q(ram[15322]) );
  DFF ram_reg_132__1_ ( .D(n19562), .CP(wclk), .Q(ram[15321]) );
  DFF ram_reg_132__0_ ( .D(n19561), .CP(wclk), .Q(ram[15320]) );
  DFF ram_reg_144__7_ ( .D(n19472), .CP(wclk), .Q(ram[15231]) );
  DFF ram_reg_144__6_ ( .D(n19471), .CP(wclk), .Q(ram[15230]) );
  DFF ram_reg_144__5_ ( .D(n19470), .CP(wclk), .Q(ram[15229]) );
  DFF ram_reg_144__4_ ( .D(n19469), .CP(wclk), .Q(ram[15228]) );
  DFF ram_reg_144__3_ ( .D(n19468), .CP(wclk), .Q(ram[15227]) );
  DFF ram_reg_144__2_ ( .D(n19467), .CP(wclk), .Q(ram[15226]) );
  DFF ram_reg_144__1_ ( .D(n19466), .CP(wclk), .Q(ram[15225]) );
  DFF ram_reg_144__0_ ( .D(n19465), .CP(wclk), .Q(ram[15224]) );
  DFF ram_reg_148__7_ ( .D(n19440), .CP(wclk), .Q(ram[15199]) );
  DFF ram_reg_148__6_ ( .D(n19439), .CP(wclk), .Q(ram[15198]) );
  DFF ram_reg_148__5_ ( .D(n19438), .CP(wclk), .Q(ram[15197]) );
  DFF ram_reg_148__4_ ( .D(n19437), .CP(wclk), .Q(ram[15196]) );
  DFF ram_reg_148__3_ ( .D(n19436), .CP(wclk), .Q(ram[15195]) );
  DFF ram_reg_148__2_ ( .D(n19435), .CP(wclk), .Q(ram[15194]) );
  DFF ram_reg_148__1_ ( .D(n19434), .CP(wclk), .Q(ram[15193]) );
  DFF ram_reg_148__0_ ( .D(n19433), .CP(wclk), .Q(ram[15192]) );
  DFF ram_reg_156__7_ ( .D(n19376), .CP(wclk), .Q(ram[15135]) );
  DFF ram_reg_156__6_ ( .D(n19375), .CP(wclk), .Q(ram[15134]) );
  DFF ram_reg_156__5_ ( .D(n19374), .CP(wclk), .Q(ram[15133]) );
  DFF ram_reg_156__4_ ( .D(n19373), .CP(wclk), .Q(ram[15132]) );
  DFF ram_reg_156__3_ ( .D(n19372), .CP(wclk), .Q(ram[15131]) );
  DFF ram_reg_156__2_ ( .D(n19371), .CP(wclk), .Q(ram[15130]) );
  DFF ram_reg_156__1_ ( .D(n19370), .CP(wclk), .Q(ram[15129]) );
  DFF ram_reg_156__0_ ( .D(n19369), .CP(wclk), .Q(ram[15128]) );
  DFF ram_reg_164__7_ ( .D(n19312), .CP(wclk), .Q(ram[15071]) );
  DFF ram_reg_164__6_ ( .D(n19311), .CP(wclk), .Q(ram[15070]) );
  DFF ram_reg_164__5_ ( .D(n19310), .CP(wclk), .Q(ram[15069]) );
  DFF ram_reg_164__4_ ( .D(n19309), .CP(wclk), .Q(ram[15068]) );
  DFF ram_reg_164__3_ ( .D(n19308), .CP(wclk), .Q(ram[15067]) );
  DFF ram_reg_164__2_ ( .D(n19307), .CP(wclk), .Q(ram[15066]) );
  DFF ram_reg_164__1_ ( .D(n19306), .CP(wclk), .Q(ram[15065]) );
  DFF ram_reg_164__0_ ( .D(n19305), .CP(wclk), .Q(ram[15064]) );
  DFF ram_reg_180__7_ ( .D(n19184), .CP(wclk), .Q(ram[14943]) );
  DFF ram_reg_180__6_ ( .D(n19183), .CP(wclk), .Q(ram[14942]) );
  DFF ram_reg_180__5_ ( .D(n19182), .CP(wclk), .Q(ram[14941]) );
  DFF ram_reg_180__4_ ( .D(n19181), .CP(wclk), .Q(ram[14940]) );
  DFF ram_reg_180__3_ ( .D(n19180), .CP(wclk), .Q(ram[14939]) );
  DFF ram_reg_180__2_ ( .D(n19179), .CP(wclk), .Q(ram[14938]) );
  DFF ram_reg_180__1_ ( .D(n19178), .CP(wclk), .Q(ram[14937]) );
  DFF ram_reg_180__0_ ( .D(n19177), .CP(wclk), .Q(ram[14936]) );
  DFF ram_reg_192__7_ ( .D(n19088), .CP(wclk), .Q(ram[14847]) );
  DFF ram_reg_192__6_ ( .D(n19087), .CP(wclk), .Q(ram[14846]) );
  DFF ram_reg_192__5_ ( .D(n19086), .CP(wclk), .Q(ram[14845]) );
  DFF ram_reg_192__4_ ( .D(n19085), .CP(wclk), .Q(ram[14844]) );
  DFF ram_reg_192__3_ ( .D(n19084), .CP(wclk), .Q(ram[14843]) );
  DFF ram_reg_192__2_ ( .D(n19083), .CP(wclk), .Q(ram[14842]) );
  DFF ram_reg_192__1_ ( .D(n19082), .CP(wclk), .Q(ram[14841]) );
  DFF ram_reg_192__0_ ( .D(n19081), .CP(wclk), .Q(ram[14840]) );
  DFF ram_reg_196__7_ ( .D(n19056), .CP(wclk), .Q(ram[14815]) );
  DFF ram_reg_196__6_ ( .D(n19055), .CP(wclk), .Q(ram[14814]) );
  DFF ram_reg_196__5_ ( .D(n19054), .CP(wclk), .Q(ram[14813]) );
  DFF ram_reg_196__4_ ( .D(n19053), .CP(wclk), .Q(ram[14812]) );
  DFF ram_reg_196__3_ ( .D(n19052), .CP(wclk), .Q(ram[14811]) );
  DFF ram_reg_196__2_ ( .D(n19051), .CP(wclk), .Q(ram[14810]) );
  DFF ram_reg_196__1_ ( .D(n19050), .CP(wclk), .Q(ram[14809]) );
  DFF ram_reg_196__0_ ( .D(n19049), .CP(wclk), .Q(ram[14808]) );
  DFF ram_reg_204__7_ ( .D(n18992), .CP(wclk), .Q(ram[14751]) );
  DFF ram_reg_204__6_ ( .D(n18991), .CP(wclk), .Q(ram[14750]) );
  DFF ram_reg_204__5_ ( .D(n18990), .CP(wclk), .Q(ram[14749]) );
  DFF ram_reg_204__4_ ( .D(n18989), .CP(wclk), .Q(ram[14748]) );
  DFF ram_reg_204__3_ ( .D(n18988), .CP(wclk), .Q(ram[14747]) );
  DFF ram_reg_204__2_ ( .D(n18987), .CP(wclk), .Q(ram[14746]) );
  DFF ram_reg_204__1_ ( .D(n18986), .CP(wclk), .Q(ram[14745]) );
  DFF ram_reg_204__0_ ( .D(n18985), .CP(wclk), .Q(ram[14744]) );
  DFF ram_reg_208__7_ ( .D(n18960), .CP(wclk), .Q(ram[14719]) );
  DFF ram_reg_208__6_ ( .D(n18959), .CP(wclk), .Q(ram[14718]) );
  DFF ram_reg_208__5_ ( .D(n18958), .CP(wclk), .Q(ram[14717]) );
  DFF ram_reg_208__4_ ( .D(n18957), .CP(wclk), .Q(ram[14716]) );
  DFF ram_reg_208__3_ ( .D(n18956), .CP(wclk), .Q(ram[14715]) );
  DFF ram_reg_208__2_ ( .D(n18955), .CP(wclk), .Q(ram[14714]) );
  DFF ram_reg_208__1_ ( .D(n18954), .CP(wclk), .Q(ram[14713]) );
  DFF ram_reg_208__0_ ( .D(n18953), .CP(wclk), .Q(ram[14712]) );
  DFF ram_reg_212__7_ ( .D(n18928), .CP(wclk), .Q(ram[14687]) );
  DFF ram_reg_212__6_ ( .D(n18927), .CP(wclk), .Q(ram[14686]) );
  DFF ram_reg_212__5_ ( .D(n18926), .CP(wclk), .Q(ram[14685]) );
  DFF ram_reg_212__4_ ( .D(n18925), .CP(wclk), .Q(ram[14684]) );
  DFF ram_reg_212__3_ ( .D(n18924), .CP(wclk), .Q(ram[14683]) );
  DFF ram_reg_212__2_ ( .D(n18923), .CP(wclk), .Q(ram[14682]) );
  DFF ram_reg_212__1_ ( .D(n18922), .CP(wclk), .Q(ram[14681]) );
  DFF ram_reg_212__0_ ( .D(n18921), .CP(wclk), .Q(ram[14680]) );
  DFF ram_reg_216__7_ ( .D(n18896), .CP(wclk), .Q(ram[14655]) );
  DFF ram_reg_216__6_ ( .D(n18895), .CP(wclk), .Q(ram[14654]) );
  DFF ram_reg_216__5_ ( .D(n18894), .CP(wclk), .Q(ram[14653]) );
  DFF ram_reg_216__4_ ( .D(n18893), .CP(wclk), .Q(ram[14652]) );
  DFF ram_reg_216__3_ ( .D(n18892), .CP(wclk), .Q(ram[14651]) );
  DFF ram_reg_216__2_ ( .D(n18891), .CP(wclk), .Q(ram[14650]) );
  DFF ram_reg_216__1_ ( .D(n18890), .CP(wclk), .Q(ram[14649]) );
  DFF ram_reg_216__0_ ( .D(n18889), .CP(wclk), .Q(ram[14648]) );
  DFF ram_reg_220__7_ ( .D(n18864), .CP(wclk), .Q(ram[14623]) );
  DFF ram_reg_220__6_ ( .D(n18863), .CP(wclk), .Q(ram[14622]) );
  DFF ram_reg_220__5_ ( .D(n18862), .CP(wclk), .Q(ram[14621]) );
  DFF ram_reg_220__4_ ( .D(n18861), .CP(wclk), .Q(ram[14620]) );
  DFF ram_reg_220__3_ ( .D(n18860), .CP(wclk), .Q(ram[14619]) );
  DFF ram_reg_220__2_ ( .D(n18859), .CP(wclk), .Q(ram[14618]) );
  DFF ram_reg_220__1_ ( .D(n18858), .CP(wclk), .Q(ram[14617]) );
  DFF ram_reg_220__0_ ( .D(n18857), .CP(wclk), .Q(ram[14616]) );
  DFF ram_reg_224__7_ ( .D(n18832), .CP(wclk), .Q(ram[14591]) );
  DFF ram_reg_224__6_ ( .D(n18831), .CP(wclk), .Q(ram[14590]) );
  DFF ram_reg_224__5_ ( .D(n18830), .CP(wclk), .Q(ram[14589]) );
  DFF ram_reg_224__4_ ( .D(n18829), .CP(wclk), .Q(ram[14588]) );
  DFF ram_reg_224__3_ ( .D(n18828), .CP(wclk), .Q(ram[14587]) );
  DFF ram_reg_224__2_ ( .D(n18827), .CP(wclk), .Q(ram[14586]) );
  DFF ram_reg_224__1_ ( .D(n18826), .CP(wclk), .Q(ram[14585]) );
  DFF ram_reg_224__0_ ( .D(n18825), .CP(wclk), .Q(ram[14584]) );
  DFF ram_reg_228__7_ ( .D(n18800), .CP(wclk), .Q(ram[14559]) );
  DFF ram_reg_228__6_ ( .D(n18799), .CP(wclk), .Q(ram[14558]) );
  DFF ram_reg_228__5_ ( .D(n18798), .CP(wclk), .Q(ram[14557]) );
  DFF ram_reg_228__4_ ( .D(n18797), .CP(wclk), .Q(ram[14556]) );
  DFF ram_reg_228__3_ ( .D(n18796), .CP(wclk), .Q(ram[14555]) );
  DFF ram_reg_228__2_ ( .D(n18795), .CP(wclk), .Q(ram[14554]) );
  DFF ram_reg_228__1_ ( .D(n18794), .CP(wclk), .Q(ram[14553]) );
  DFF ram_reg_228__0_ ( .D(n18793), .CP(wclk), .Q(ram[14552]) );
  DFF ram_reg_240__7_ ( .D(n18704), .CP(wclk), .Q(ram[14463]) );
  DFF ram_reg_240__6_ ( .D(n18703), .CP(wclk), .Q(ram[14462]) );
  DFF ram_reg_240__5_ ( .D(n18702), .CP(wclk), .Q(ram[14461]) );
  DFF ram_reg_240__4_ ( .D(n18701), .CP(wclk), .Q(ram[14460]) );
  DFF ram_reg_240__3_ ( .D(n18700), .CP(wclk), .Q(ram[14459]) );
  DFF ram_reg_240__2_ ( .D(n18699), .CP(wclk), .Q(ram[14458]) );
  DFF ram_reg_240__1_ ( .D(n18698), .CP(wclk), .Q(ram[14457]) );
  DFF ram_reg_240__0_ ( .D(n18697), .CP(wclk), .Q(ram[14456]) );
  DFF ram_reg_244__7_ ( .D(n18672), .CP(wclk), .Q(ram[14431]) );
  DFF ram_reg_244__6_ ( .D(n18671), .CP(wclk), .Q(ram[14430]) );
  DFF ram_reg_244__5_ ( .D(n18670), .CP(wclk), .Q(ram[14429]) );
  DFF ram_reg_244__4_ ( .D(n18669), .CP(wclk), .Q(ram[14428]) );
  DFF ram_reg_244__3_ ( .D(n18668), .CP(wclk), .Q(ram[14427]) );
  DFF ram_reg_244__2_ ( .D(n18667), .CP(wclk), .Q(ram[14426]) );
  DFF ram_reg_244__1_ ( .D(n18666), .CP(wclk), .Q(ram[14425]) );
  DFF ram_reg_244__0_ ( .D(n18665), .CP(wclk), .Q(ram[14424]) );
  DFF ram_reg_256__7_ ( .D(n18576), .CP(wclk), .Q(ram[14335]) );
  DFF ram_reg_256__6_ ( .D(n18575), .CP(wclk), .Q(ram[14334]) );
  DFF ram_reg_256__5_ ( .D(n18574), .CP(wclk), .Q(ram[14333]) );
  DFF ram_reg_256__4_ ( .D(n18573), .CP(wclk), .Q(ram[14332]) );
  DFF ram_reg_256__3_ ( .D(n18572), .CP(wclk), .Q(ram[14331]) );
  DFF ram_reg_256__2_ ( .D(n18571), .CP(wclk), .Q(ram[14330]) );
  DFF ram_reg_256__1_ ( .D(n18570), .CP(wclk), .Q(ram[14329]) );
  DFF ram_reg_256__0_ ( .D(n18569), .CP(wclk), .Q(ram[14328]) );
  DFF ram_reg_260__7_ ( .D(n18544), .CP(wclk), .Q(ram[14303]) );
  DFF ram_reg_260__6_ ( .D(n18543), .CP(wclk), .Q(ram[14302]) );
  DFF ram_reg_260__5_ ( .D(n18542), .CP(wclk), .Q(ram[14301]) );
  DFF ram_reg_260__4_ ( .D(n18541), .CP(wclk), .Q(ram[14300]) );
  DFF ram_reg_260__3_ ( .D(n18540), .CP(wclk), .Q(ram[14299]) );
  DFF ram_reg_260__2_ ( .D(n18539), .CP(wclk), .Q(ram[14298]) );
  DFF ram_reg_260__1_ ( .D(n18538), .CP(wclk), .Q(ram[14297]) );
  DFF ram_reg_260__0_ ( .D(n18537), .CP(wclk), .Q(ram[14296]) );
  DFF ram_reg_264__7_ ( .D(n18512), .CP(wclk), .Q(ram[14271]) );
  DFF ram_reg_264__6_ ( .D(n18511), .CP(wclk), .Q(ram[14270]) );
  DFF ram_reg_264__5_ ( .D(n18510), .CP(wclk), .Q(ram[14269]) );
  DFF ram_reg_264__4_ ( .D(n18509), .CP(wclk), .Q(ram[14268]) );
  DFF ram_reg_264__3_ ( .D(n18508), .CP(wclk), .Q(ram[14267]) );
  DFF ram_reg_264__2_ ( .D(n18507), .CP(wclk), .Q(ram[14266]) );
  DFF ram_reg_264__1_ ( .D(n18506), .CP(wclk), .Q(ram[14265]) );
  DFF ram_reg_264__0_ ( .D(n18505), .CP(wclk), .Q(ram[14264]) );
  DFF ram_reg_268__7_ ( .D(n18480), .CP(wclk), .Q(ram[14239]) );
  DFF ram_reg_268__6_ ( .D(n18479), .CP(wclk), .Q(ram[14238]) );
  DFF ram_reg_268__5_ ( .D(n18478), .CP(wclk), .Q(ram[14237]) );
  DFF ram_reg_268__4_ ( .D(n18477), .CP(wclk), .Q(ram[14236]) );
  DFF ram_reg_268__3_ ( .D(n18476), .CP(wclk), .Q(ram[14235]) );
  DFF ram_reg_268__2_ ( .D(n18475), .CP(wclk), .Q(ram[14234]) );
  DFF ram_reg_268__1_ ( .D(n18474), .CP(wclk), .Q(ram[14233]) );
  DFF ram_reg_268__0_ ( .D(n18473), .CP(wclk), .Q(ram[14232]) );
  DFF ram_reg_272__7_ ( .D(n18448), .CP(wclk), .Q(ram[14207]) );
  DFF ram_reg_272__6_ ( .D(n18447), .CP(wclk), .Q(ram[14206]) );
  DFF ram_reg_272__5_ ( .D(n18446), .CP(wclk), .Q(ram[14205]) );
  DFF ram_reg_272__4_ ( .D(n18445), .CP(wclk), .Q(ram[14204]) );
  DFF ram_reg_272__3_ ( .D(n18444), .CP(wclk), .Q(ram[14203]) );
  DFF ram_reg_272__2_ ( .D(n18443), .CP(wclk), .Q(ram[14202]) );
  DFF ram_reg_272__1_ ( .D(n18442), .CP(wclk), .Q(ram[14201]) );
  DFF ram_reg_272__0_ ( .D(n18441), .CP(wclk), .Q(ram[14200]) );
  DFF ram_reg_276__7_ ( .D(n18416), .CP(wclk), .Q(ram[14175]) );
  DFF ram_reg_276__6_ ( .D(n18415), .CP(wclk), .Q(ram[14174]) );
  DFF ram_reg_276__5_ ( .D(n18414), .CP(wclk), .Q(ram[14173]) );
  DFF ram_reg_276__4_ ( .D(n18413), .CP(wclk), .Q(ram[14172]) );
  DFF ram_reg_276__3_ ( .D(n18412), .CP(wclk), .Q(ram[14171]) );
  DFF ram_reg_276__2_ ( .D(n18411), .CP(wclk), .Q(ram[14170]) );
  DFF ram_reg_276__1_ ( .D(n18410), .CP(wclk), .Q(ram[14169]) );
  DFF ram_reg_276__0_ ( .D(n18409), .CP(wclk), .Q(ram[14168]) );
  DFF ram_reg_280__7_ ( .D(n18384), .CP(wclk), .Q(ram[14143]) );
  DFF ram_reg_280__6_ ( .D(n18383), .CP(wclk), .Q(ram[14142]) );
  DFF ram_reg_280__5_ ( .D(n18382), .CP(wclk), .Q(ram[14141]) );
  DFF ram_reg_280__4_ ( .D(n18381), .CP(wclk), .Q(ram[14140]) );
  DFF ram_reg_280__3_ ( .D(n18380), .CP(wclk), .Q(ram[14139]) );
  DFF ram_reg_280__2_ ( .D(n18379), .CP(wclk), .Q(ram[14138]) );
  DFF ram_reg_280__1_ ( .D(n18378), .CP(wclk), .Q(ram[14137]) );
  DFF ram_reg_280__0_ ( .D(n18377), .CP(wclk), .Q(ram[14136]) );
  DFF ram_reg_284__7_ ( .D(n18352), .CP(wclk), .Q(ram[14111]) );
  DFF ram_reg_284__6_ ( .D(n18351), .CP(wclk), .Q(ram[14110]) );
  DFF ram_reg_284__5_ ( .D(n18350), .CP(wclk), .Q(ram[14109]) );
  DFF ram_reg_284__4_ ( .D(n18349), .CP(wclk), .Q(ram[14108]) );
  DFF ram_reg_284__3_ ( .D(n18348), .CP(wclk), .Q(ram[14107]) );
  DFF ram_reg_284__2_ ( .D(n18347), .CP(wclk), .Q(ram[14106]) );
  DFF ram_reg_284__1_ ( .D(n18346), .CP(wclk), .Q(ram[14105]) );
  DFF ram_reg_284__0_ ( .D(n18345), .CP(wclk), .Q(ram[14104]) );
  DFF ram_reg_288__7_ ( .D(n18320), .CP(wclk), .Q(ram[14079]) );
  DFF ram_reg_288__6_ ( .D(n18319), .CP(wclk), .Q(ram[14078]) );
  DFF ram_reg_288__5_ ( .D(n18318), .CP(wclk), .Q(ram[14077]) );
  DFF ram_reg_288__4_ ( .D(n18317), .CP(wclk), .Q(ram[14076]) );
  DFF ram_reg_288__3_ ( .D(n18316), .CP(wclk), .Q(ram[14075]) );
  DFF ram_reg_288__2_ ( .D(n18315), .CP(wclk), .Q(ram[14074]) );
  DFF ram_reg_288__1_ ( .D(n18314), .CP(wclk), .Q(ram[14073]) );
  DFF ram_reg_288__0_ ( .D(n18313), .CP(wclk), .Q(ram[14072]) );
  DFF ram_reg_292__7_ ( .D(n18288), .CP(wclk), .Q(ram[14047]) );
  DFF ram_reg_292__6_ ( .D(n18287), .CP(wclk), .Q(ram[14046]) );
  DFF ram_reg_292__5_ ( .D(n18286), .CP(wclk), .Q(ram[14045]) );
  DFF ram_reg_292__4_ ( .D(n18285), .CP(wclk), .Q(ram[14044]) );
  DFF ram_reg_292__3_ ( .D(n18284), .CP(wclk), .Q(ram[14043]) );
  DFF ram_reg_292__2_ ( .D(n18283), .CP(wclk), .Q(ram[14042]) );
  DFF ram_reg_292__1_ ( .D(n18282), .CP(wclk), .Q(ram[14041]) );
  DFF ram_reg_292__0_ ( .D(n18281), .CP(wclk), .Q(ram[14040]) );
  DFF ram_reg_300__7_ ( .D(n18224), .CP(wclk), .Q(ram[13983]) );
  DFF ram_reg_300__6_ ( .D(n18223), .CP(wclk), .Q(ram[13982]) );
  DFF ram_reg_300__5_ ( .D(n18222), .CP(wclk), .Q(ram[13981]) );
  DFF ram_reg_300__4_ ( .D(n18221), .CP(wclk), .Q(ram[13980]) );
  DFF ram_reg_300__3_ ( .D(n18220), .CP(wclk), .Q(ram[13979]) );
  DFF ram_reg_300__2_ ( .D(n18219), .CP(wclk), .Q(ram[13978]) );
  DFF ram_reg_300__1_ ( .D(n18218), .CP(wclk), .Q(ram[13977]) );
  DFF ram_reg_300__0_ ( .D(n18217), .CP(wclk), .Q(ram[13976]) );
  DFF ram_reg_304__7_ ( .D(n18192), .CP(wclk), .Q(ram[13951]) );
  DFF ram_reg_304__6_ ( .D(n18191), .CP(wclk), .Q(ram[13950]) );
  DFF ram_reg_304__5_ ( .D(n18190), .CP(wclk), .Q(ram[13949]) );
  DFF ram_reg_304__4_ ( .D(n18189), .CP(wclk), .Q(ram[13948]) );
  DFF ram_reg_304__3_ ( .D(n18188), .CP(wclk), .Q(ram[13947]) );
  DFF ram_reg_304__2_ ( .D(n18187), .CP(wclk), .Q(ram[13946]) );
  DFF ram_reg_304__1_ ( .D(n18186), .CP(wclk), .Q(ram[13945]) );
  DFF ram_reg_304__0_ ( .D(n18185), .CP(wclk), .Q(ram[13944]) );
  DFF ram_reg_308__7_ ( .D(n18160), .CP(wclk), .Q(ram[13919]) );
  DFF ram_reg_308__6_ ( .D(n18159), .CP(wclk), .Q(ram[13918]) );
  DFF ram_reg_308__5_ ( .D(n18158), .CP(wclk), .Q(ram[13917]) );
  DFF ram_reg_308__4_ ( .D(n18157), .CP(wclk), .Q(ram[13916]) );
  DFF ram_reg_308__3_ ( .D(n18156), .CP(wclk), .Q(ram[13915]) );
  DFF ram_reg_308__2_ ( .D(n18155), .CP(wclk), .Q(ram[13914]) );
  DFF ram_reg_308__1_ ( .D(n18154), .CP(wclk), .Q(ram[13913]) );
  DFF ram_reg_308__0_ ( .D(n18153), .CP(wclk), .Q(ram[13912]) );
  DFF ram_reg_320__7_ ( .D(n18064), .CP(wclk), .Q(ram[13823]) );
  DFF ram_reg_320__6_ ( .D(n18063), .CP(wclk), .Q(ram[13822]) );
  DFF ram_reg_320__5_ ( .D(n18062), .CP(wclk), .Q(ram[13821]) );
  DFF ram_reg_320__4_ ( .D(n18061), .CP(wclk), .Q(ram[13820]) );
  DFF ram_reg_320__3_ ( .D(n18060), .CP(wclk), .Q(ram[13819]) );
  DFF ram_reg_320__2_ ( .D(n18059), .CP(wclk), .Q(ram[13818]) );
  DFF ram_reg_320__1_ ( .D(n18058), .CP(wclk), .Q(ram[13817]) );
  DFF ram_reg_320__0_ ( .D(n18057), .CP(wclk), .Q(ram[13816]) );
  DFF ram_reg_324__7_ ( .D(n18032), .CP(wclk), .Q(ram[13791]) );
  DFF ram_reg_324__6_ ( .D(n18031), .CP(wclk), .Q(ram[13790]) );
  DFF ram_reg_324__5_ ( .D(n18030), .CP(wclk), .Q(ram[13789]) );
  DFF ram_reg_324__4_ ( .D(n18029), .CP(wclk), .Q(ram[13788]) );
  DFF ram_reg_324__3_ ( .D(n18028), .CP(wclk), .Q(ram[13787]) );
  DFF ram_reg_324__2_ ( .D(n18027), .CP(wclk), .Q(ram[13786]) );
  DFF ram_reg_324__1_ ( .D(n18026), .CP(wclk), .Q(ram[13785]) );
  DFF ram_reg_324__0_ ( .D(n18025), .CP(wclk), .Q(ram[13784]) );
  DFF ram_reg_328__7_ ( .D(n18000), .CP(wclk), .Q(ram[13759]) );
  DFF ram_reg_328__6_ ( .D(n17999), .CP(wclk), .Q(ram[13758]) );
  DFF ram_reg_328__5_ ( .D(n17998), .CP(wclk), .Q(ram[13757]) );
  DFF ram_reg_328__4_ ( .D(n17997), .CP(wclk), .Q(ram[13756]) );
  DFF ram_reg_328__3_ ( .D(n17996), .CP(wclk), .Q(ram[13755]) );
  DFF ram_reg_328__2_ ( .D(n17995), .CP(wclk), .Q(ram[13754]) );
  DFF ram_reg_328__1_ ( .D(n17994), .CP(wclk), .Q(ram[13753]) );
  DFF ram_reg_328__0_ ( .D(n17993), .CP(wclk), .Q(ram[13752]) );
  DFF ram_reg_332__7_ ( .D(n17968), .CP(wclk), .Q(ram[13727]) );
  DFF ram_reg_332__6_ ( .D(n17967), .CP(wclk), .Q(ram[13726]) );
  DFF ram_reg_332__5_ ( .D(n17966), .CP(wclk), .Q(ram[13725]) );
  DFF ram_reg_332__4_ ( .D(n17965), .CP(wclk), .Q(ram[13724]) );
  DFF ram_reg_332__3_ ( .D(n17964), .CP(wclk), .Q(ram[13723]) );
  DFF ram_reg_332__2_ ( .D(n17963), .CP(wclk), .Q(ram[13722]) );
  DFF ram_reg_332__1_ ( .D(n17962), .CP(wclk), .Q(ram[13721]) );
  DFF ram_reg_332__0_ ( .D(n17961), .CP(wclk), .Q(ram[13720]) );
  DFF ram_reg_336__7_ ( .D(n17936), .CP(wclk), .Q(ram[13695]) );
  DFF ram_reg_336__6_ ( .D(n17935), .CP(wclk), .Q(ram[13694]) );
  DFF ram_reg_336__5_ ( .D(n17934), .CP(wclk), .Q(ram[13693]) );
  DFF ram_reg_336__4_ ( .D(n17933), .CP(wclk), .Q(ram[13692]) );
  DFF ram_reg_336__3_ ( .D(n17932), .CP(wclk), .Q(ram[13691]) );
  DFF ram_reg_336__2_ ( .D(n17931), .CP(wclk), .Q(ram[13690]) );
  DFF ram_reg_336__1_ ( .D(n17930), .CP(wclk), .Q(ram[13689]) );
  DFF ram_reg_336__0_ ( .D(n17929), .CP(wclk), .Q(ram[13688]) );
  DFF ram_reg_340__7_ ( .D(n17904), .CP(wclk), .Q(ram[13663]) );
  DFF ram_reg_340__6_ ( .D(n17903), .CP(wclk), .Q(ram[13662]) );
  DFF ram_reg_340__5_ ( .D(n17902), .CP(wclk), .Q(ram[13661]) );
  DFF ram_reg_340__4_ ( .D(n17901), .CP(wclk), .Q(ram[13660]) );
  DFF ram_reg_340__3_ ( .D(n17900), .CP(wclk), .Q(ram[13659]) );
  DFF ram_reg_340__2_ ( .D(n17899), .CP(wclk), .Q(ram[13658]) );
  DFF ram_reg_340__1_ ( .D(n17898), .CP(wclk), .Q(ram[13657]) );
  DFF ram_reg_340__0_ ( .D(n17897), .CP(wclk), .Q(ram[13656]) );
  DFF ram_reg_344__7_ ( .D(n17872), .CP(wclk), .Q(ram[13631]) );
  DFF ram_reg_344__6_ ( .D(n17871), .CP(wclk), .Q(ram[13630]) );
  DFF ram_reg_344__5_ ( .D(n17870), .CP(wclk), .Q(ram[13629]) );
  DFF ram_reg_344__4_ ( .D(n17869), .CP(wclk), .Q(ram[13628]) );
  DFF ram_reg_344__3_ ( .D(n17868), .CP(wclk), .Q(ram[13627]) );
  DFF ram_reg_344__2_ ( .D(n17867), .CP(wclk), .Q(ram[13626]) );
  DFF ram_reg_344__1_ ( .D(n17866), .CP(wclk), .Q(ram[13625]) );
  DFF ram_reg_344__0_ ( .D(n17865), .CP(wclk), .Q(ram[13624]) );
  DFF ram_reg_348__7_ ( .D(n17840), .CP(wclk), .Q(ram[13599]) );
  DFF ram_reg_348__6_ ( .D(n17839), .CP(wclk), .Q(ram[13598]) );
  DFF ram_reg_348__5_ ( .D(n17838), .CP(wclk), .Q(ram[13597]) );
  DFF ram_reg_348__4_ ( .D(n17837), .CP(wclk), .Q(ram[13596]) );
  DFF ram_reg_348__3_ ( .D(n17836), .CP(wclk), .Q(ram[13595]) );
  DFF ram_reg_348__2_ ( .D(n17835), .CP(wclk), .Q(ram[13594]) );
  DFF ram_reg_348__1_ ( .D(n17834), .CP(wclk), .Q(ram[13593]) );
  DFF ram_reg_348__0_ ( .D(n17833), .CP(wclk), .Q(ram[13592]) );
  DFF ram_reg_352__7_ ( .D(n17808), .CP(wclk), .Q(ram[13567]) );
  DFF ram_reg_352__6_ ( .D(n17807), .CP(wclk), .Q(ram[13566]) );
  DFF ram_reg_352__5_ ( .D(n17806), .CP(wclk), .Q(ram[13565]) );
  DFF ram_reg_352__4_ ( .D(n17805), .CP(wclk), .Q(ram[13564]) );
  DFF ram_reg_352__3_ ( .D(n17804), .CP(wclk), .Q(ram[13563]) );
  DFF ram_reg_352__2_ ( .D(n17803), .CP(wclk), .Q(ram[13562]) );
  DFF ram_reg_352__1_ ( .D(n17802), .CP(wclk), .Q(ram[13561]) );
  DFF ram_reg_352__0_ ( .D(n17801), .CP(wclk), .Q(ram[13560]) );
  DFF ram_reg_356__7_ ( .D(n17776), .CP(wclk), .Q(ram[13535]) );
  DFF ram_reg_356__6_ ( .D(n17775), .CP(wclk), .Q(ram[13534]) );
  DFF ram_reg_356__5_ ( .D(n17774), .CP(wclk), .Q(ram[13533]) );
  DFF ram_reg_356__4_ ( .D(n17773), .CP(wclk), .Q(ram[13532]) );
  DFF ram_reg_356__3_ ( .D(n17772), .CP(wclk), .Q(ram[13531]) );
  DFF ram_reg_356__2_ ( .D(n17771), .CP(wclk), .Q(ram[13530]) );
  DFF ram_reg_356__1_ ( .D(n17770), .CP(wclk), .Q(ram[13529]) );
  DFF ram_reg_356__0_ ( .D(n17769), .CP(wclk), .Q(ram[13528]) );
  DFF ram_reg_360__7_ ( .D(n17744), .CP(wclk), .Q(ram[13503]) );
  DFF ram_reg_360__6_ ( .D(n17743), .CP(wclk), .Q(ram[13502]) );
  DFF ram_reg_360__5_ ( .D(n17742), .CP(wclk), .Q(ram[13501]) );
  DFF ram_reg_360__4_ ( .D(n17741), .CP(wclk), .Q(ram[13500]) );
  DFF ram_reg_360__3_ ( .D(n17740), .CP(wclk), .Q(ram[13499]) );
  DFF ram_reg_360__2_ ( .D(n17739), .CP(wclk), .Q(ram[13498]) );
  DFF ram_reg_360__1_ ( .D(n17738), .CP(wclk), .Q(ram[13497]) );
  DFF ram_reg_360__0_ ( .D(n17737), .CP(wclk), .Q(ram[13496]) );
  DFF ram_reg_364__7_ ( .D(n17712), .CP(wclk), .Q(ram[13471]) );
  DFF ram_reg_364__6_ ( .D(n17711), .CP(wclk), .Q(ram[13470]) );
  DFF ram_reg_364__5_ ( .D(n17710), .CP(wclk), .Q(ram[13469]) );
  DFF ram_reg_364__4_ ( .D(n17709), .CP(wclk), .Q(ram[13468]) );
  DFF ram_reg_364__3_ ( .D(n17708), .CP(wclk), .Q(ram[13467]) );
  DFF ram_reg_364__2_ ( .D(n17707), .CP(wclk), .Q(ram[13466]) );
  DFF ram_reg_364__1_ ( .D(n17706), .CP(wclk), .Q(ram[13465]) );
  DFF ram_reg_364__0_ ( .D(n17705), .CP(wclk), .Q(ram[13464]) );
  DFF ram_reg_368__7_ ( .D(n17680), .CP(wclk), .Q(ram[13439]) );
  DFF ram_reg_368__6_ ( .D(n17679), .CP(wclk), .Q(ram[13438]) );
  DFF ram_reg_368__5_ ( .D(n17678), .CP(wclk), .Q(ram[13437]) );
  DFF ram_reg_368__4_ ( .D(n17677), .CP(wclk), .Q(ram[13436]) );
  DFF ram_reg_368__3_ ( .D(n17676), .CP(wclk), .Q(ram[13435]) );
  DFF ram_reg_368__2_ ( .D(n17675), .CP(wclk), .Q(ram[13434]) );
  DFF ram_reg_368__1_ ( .D(n17674), .CP(wclk), .Q(ram[13433]) );
  DFF ram_reg_368__0_ ( .D(n17673), .CP(wclk), .Q(ram[13432]) );
  DFF ram_reg_372__7_ ( .D(n17648), .CP(wclk), .Q(ram[13407]) );
  DFF ram_reg_372__6_ ( .D(n17647), .CP(wclk), .Q(ram[13406]) );
  DFF ram_reg_372__5_ ( .D(n17646), .CP(wclk), .Q(ram[13405]) );
  DFF ram_reg_372__4_ ( .D(n17645), .CP(wclk), .Q(ram[13404]) );
  DFF ram_reg_372__3_ ( .D(n17644), .CP(wclk), .Q(ram[13403]) );
  DFF ram_reg_372__2_ ( .D(n17643), .CP(wclk), .Q(ram[13402]) );
  DFF ram_reg_372__1_ ( .D(n17642), .CP(wclk), .Q(ram[13401]) );
  DFF ram_reg_372__0_ ( .D(n17641), .CP(wclk), .Q(ram[13400]) );
  DFF ram_reg_376__7_ ( .D(n17616), .CP(wclk), .Q(ram[13375]) );
  DFF ram_reg_376__6_ ( .D(n17615), .CP(wclk), .Q(ram[13374]) );
  DFF ram_reg_376__5_ ( .D(n17614), .CP(wclk), .Q(ram[13373]) );
  DFF ram_reg_376__4_ ( .D(n17613), .CP(wclk), .Q(ram[13372]) );
  DFF ram_reg_376__3_ ( .D(n17612), .CP(wclk), .Q(ram[13371]) );
  DFF ram_reg_376__2_ ( .D(n17611), .CP(wclk), .Q(ram[13370]) );
  DFF ram_reg_376__1_ ( .D(n17610), .CP(wclk), .Q(ram[13369]) );
  DFF ram_reg_376__0_ ( .D(n17609), .CP(wclk), .Q(ram[13368]) );
  DFF ram_reg_380__7_ ( .D(n17584), .CP(wclk), .Q(ram[13343]) );
  DFF ram_reg_380__6_ ( .D(n17583), .CP(wclk), .Q(ram[13342]) );
  DFF ram_reg_380__5_ ( .D(n17582), .CP(wclk), .Q(ram[13341]) );
  DFF ram_reg_380__4_ ( .D(n17581), .CP(wclk), .Q(ram[13340]) );
  DFF ram_reg_380__3_ ( .D(n17580), .CP(wclk), .Q(ram[13339]) );
  DFF ram_reg_380__2_ ( .D(n17579), .CP(wclk), .Q(ram[13338]) );
  DFF ram_reg_380__1_ ( .D(n17578), .CP(wclk), .Q(ram[13337]) );
  DFF ram_reg_380__0_ ( .D(n17577), .CP(wclk), .Q(ram[13336]) );
  DFF ram_reg_384__7_ ( .D(n17552), .CP(wclk), .Q(ram[13311]) );
  DFF ram_reg_384__6_ ( .D(n17551), .CP(wclk), .Q(ram[13310]) );
  DFF ram_reg_384__5_ ( .D(n17550), .CP(wclk), .Q(ram[13309]) );
  DFF ram_reg_384__4_ ( .D(n17549), .CP(wclk), .Q(ram[13308]) );
  DFF ram_reg_384__3_ ( .D(n17548), .CP(wclk), .Q(ram[13307]) );
  DFF ram_reg_384__2_ ( .D(n17547), .CP(wclk), .Q(ram[13306]) );
  DFF ram_reg_384__1_ ( .D(n17546), .CP(wclk), .Q(ram[13305]) );
  DFF ram_reg_384__0_ ( .D(n17545), .CP(wclk), .Q(ram[13304]) );
  DFF ram_reg_388__7_ ( .D(n17520), .CP(wclk), .Q(ram[13279]) );
  DFF ram_reg_388__6_ ( .D(n17519), .CP(wclk), .Q(ram[13278]) );
  DFF ram_reg_388__5_ ( .D(n17518), .CP(wclk), .Q(ram[13277]) );
  DFF ram_reg_388__4_ ( .D(n17517), .CP(wclk), .Q(ram[13276]) );
  DFF ram_reg_388__3_ ( .D(n17516), .CP(wclk), .Q(ram[13275]) );
  DFF ram_reg_388__2_ ( .D(n17515), .CP(wclk), .Q(ram[13274]) );
  DFF ram_reg_388__1_ ( .D(n17514), .CP(wclk), .Q(ram[13273]) );
  DFF ram_reg_388__0_ ( .D(n17513), .CP(wclk), .Q(ram[13272]) );
  DFF ram_reg_400__7_ ( .D(n17424), .CP(wclk), .Q(ram[13183]) );
  DFF ram_reg_400__6_ ( .D(n17423), .CP(wclk), .Q(ram[13182]) );
  DFF ram_reg_400__5_ ( .D(n17422), .CP(wclk), .Q(ram[13181]) );
  DFF ram_reg_400__4_ ( .D(n17421), .CP(wclk), .Q(ram[13180]) );
  DFF ram_reg_400__3_ ( .D(n17420), .CP(wclk), .Q(ram[13179]) );
  DFF ram_reg_400__2_ ( .D(n17419), .CP(wclk), .Q(ram[13178]) );
  DFF ram_reg_400__1_ ( .D(n17418), .CP(wclk), .Q(ram[13177]) );
  DFF ram_reg_400__0_ ( .D(n17417), .CP(wclk), .Q(ram[13176]) );
  DFF ram_reg_404__7_ ( .D(n17392), .CP(wclk), .Q(ram[13151]) );
  DFF ram_reg_404__6_ ( .D(n17391), .CP(wclk), .Q(ram[13150]) );
  DFF ram_reg_404__5_ ( .D(n17390), .CP(wclk), .Q(ram[13149]) );
  DFF ram_reg_404__4_ ( .D(n17389), .CP(wclk), .Q(ram[13148]) );
  DFF ram_reg_404__3_ ( .D(n17388), .CP(wclk), .Q(ram[13147]) );
  DFF ram_reg_404__2_ ( .D(n17387), .CP(wclk), .Q(ram[13146]) );
  DFF ram_reg_404__1_ ( .D(n17386), .CP(wclk), .Q(ram[13145]) );
  DFF ram_reg_404__0_ ( .D(n17385), .CP(wclk), .Q(ram[13144]) );
  DFF ram_reg_420__7_ ( .D(n17264), .CP(wclk), .Q(ram[13023]) );
  DFF ram_reg_420__6_ ( .D(n17263), .CP(wclk), .Q(ram[13022]) );
  DFF ram_reg_420__5_ ( .D(n17262), .CP(wclk), .Q(ram[13021]) );
  DFF ram_reg_420__4_ ( .D(n17261), .CP(wclk), .Q(ram[13020]) );
  DFF ram_reg_420__3_ ( .D(n17260), .CP(wclk), .Q(ram[13019]) );
  DFF ram_reg_420__2_ ( .D(n17259), .CP(wclk), .Q(ram[13018]) );
  DFF ram_reg_420__1_ ( .D(n17258), .CP(wclk), .Q(ram[13017]) );
  DFF ram_reg_420__0_ ( .D(n17257), .CP(wclk), .Q(ram[13016]) );
  DFF ram_reg_436__7_ ( .D(n17136), .CP(wclk), .Q(ram[12895]) );
  DFF ram_reg_436__6_ ( .D(n17135), .CP(wclk), .Q(ram[12894]) );
  DFF ram_reg_436__5_ ( .D(n17134), .CP(wclk), .Q(ram[12893]) );
  DFF ram_reg_436__4_ ( .D(n17133), .CP(wclk), .Q(ram[12892]) );
  DFF ram_reg_436__3_ ( .D(n17132), .CP(wclk), .Q(ram[12891]) );
  DFF ram_reg_436__2_ ( .D(n17131), .CP(wclk), .Q(ram[12890]) );
  DFF ram_reg_436__1_ ( .D(n17130), .CP(wclk), .Q(ram[12889]) );
  DFF ram_reg_436__0_ ( .D(n17129), .CP(wclk), .Q(ram[12888]) );
  DFF ram_reg_448__7_ ( .D(n17040), .CP(wclk), .Q(ram[12799]) );
  DFF ram_reg_448__6_ ( .D(n17039), .CP(wclk), .Q(ram[12798]) );
  DFF ram_reg_448__5_ ( .D(n17038), .CP(wclk), .Q(ram[12797]) );
  DFF ram_reg_448__4_ ( .D(n17037), .CP(wclk), .Q(ram[12796]) );
  DFF ram_reg_448__3_ ( .D(n17036), .CP(wclk), .Q(ram[12795]) );
  DFF ram_reg_448__2_ ( .D(n17035), .CP(wclk), .Q(ram[12794]) );
  DFF ram_reg_448__1_ ( .D(n17034), .CP(wclk), .Q(ram[12793]) );
  DFF ram_reg_448__0_ ( .D(n17033), .CP(wclk), .Q(ram[12792]) );
  DFF ram_reg_452__7_ ( .D(n17008), .CP(wclk), .Q(ram[12767]) );
  DFF ram_reg_452__6_ ( .D(n17007), .CP(wclk), .Q(ram[12766]) );
  DFF ram_reg_452__5_ ( .D(n17006), .CP(wclk), .Q(ram[12765]) );
  DFF ram_reg_452__4_ ( .D(n17005), .CP(wclk), .Q(ram[12764]) );
  DFF ram_reg_452__3_ ( .D(n17004), .CP(wclk), .Q(ram[12763]) );
  DFF ram_reg_452__2_ ( .D(n17003), .CP(wclk), .Q(ram[12762]) );
  DFF ram_reg_452__1_ ( .D(n17002), .CP(wclk), .Q(ram[12761]) );
  DFF ram_reg_452__0_ ( .D(n17001), .CP(wclk), .Q(ram[12760]) );
  DFF ram_reg_464__7_ ( .D(n16912), .CP(wclk), .Q(ram[12671]) );
  DFF ram_reg_464__6_ ( .D(n16911), .CP(wclk), .Q(ram[12670]) );
  DFF ram_reg_464__5_ ( .D(n16910), .CP(wclk), .Q(ram[12669]) );
  DFF ram_reg_464__4_ ( .D(n16909), .CP(wclk), .Q(ram[12668]) );
  DFF ram_reg_464__3_ ( .D(n16908), .CP(wclk), .Q(ram[12667]) );
  DFF ram_reg_464__2_ ( .D(n16907), .CP(wclk), .Q(ram[12666]) );
  DFF ram_reg_464__1_ ( .D(n16906), .CP(wclk), .Q(ram[12665]) );
  DFF ram_reg_464__0_ ( .D(n16905), .CP(wclk), .Q(ram[12664]) );
  DFF ram_reg_468__7_ ( .D(n16880), .CP(wclk), .Q(ram[12639]) );
  DFF ram_reg_468__6_ ( .D(n16879), .CP(wclk), .Q(ram[12638]) );
  DFF ram_reg_468__5_ ( .D(n16878), .CP(wclk), .Q(ram[12637]) );
  DFF ram_reg_468__4_ ( .D(n16877), .CP(wclk), .Q(ram[12636]) );
  DFF ram_reg_468__3_ ( .D(n16876), .CP(wclk), .Q(ram[12635]) );
  DFF ram_reg_468__2_ ( .D(n16875), .CP(wclk), .Q(ram[12634]) );
  DFF ram_reg_468__1_ ( .D(n16874), .CP(wclk), .Q(ram[12633]) );
  DFF ram_reg_468__0_ ( .D(n16873), .CP(wclk), .Q(ram[12632]) );
  DFF ram_reg_476__7_ ( .D(n16816), .CP(wclk), .Q(ram[12575]) );
  DFF ram_reg_476__6_ ( .D(n16815), .CP(wclk), .Q(ram[12574]) );
  DFF ram_reg_476__5_ ( .D(n16814), .CP(wclk), .Q(ram[12573]) );
  DFF ram_reg_476__4_ ( .D(n16813), .CP(wclk), .Q(ram[12572]) );
  DFF ram_reg_476__3_ ( .D(n16812), .CP(wclk), .Q(ram[12571]) );
  DFF ram_reg_476__2_ ( .D(n16811), .CP(wclk), .Q(ram[12570]) );
  DFF ram_reg_476__1_ ( .D(n16810), .CP(wclk), .Q(ram[12569]) );
  DFF ram_reg_476__0_ ( .D(n16809), .CP(wclk), .Q(ram[12568]) );
  DFF ram_reg_480__7_ ( .D(n16784), .CP(wclk), .Q(ram[12543]) );
  DFF ram_reg_480__6_ ( .D(n16783), .CP(wclk), .Q(ram[12542]) );
  DFF ram_reg_480__5_ ( .D(n16782), .CP(wclk), .Q(ram[12541]) );
  DFF ram_reg_480__4_ ( .D(n16781), .CP(wclk), .Q(ram[12540]) );
  DFF ram_reg_480__3_ ( .D(n16780), .CP(wclk), .Q(ram[12539]) );
  DFF ram_reg_480__2_ ( .D(n16779), .CP(wclk), .Q(ram[12538]) );
  DFF ram_reg_480__1_ ( .D(n16778), .CP(wclk), .Q(ram[12537]) );
  DFF ram_reg_480__0_ ( .D(n16777), .CP(wclk), .Q(ram[12536]) );
  DFF ram_reg_484__7_ ( .D(n16752), .CP(wclk), .Q(ram[12511]) );
  DFF ram_reg_484__6_ ( .D(n16751), .CP(wclk), .Q(ram[12510]) );
  DFF ram_reg_484__5_ ( .D(n16750), .CP(wclk), .Q(ram[12509]) );
  DFF ram_reg_484__4_ ( .D(n16749), .CP(wclk), .Q(ram[12508]) );
  DFF ram_reg_484__3_ ( .D(n16748), .CP(wclk), .Q(ram[12507]) );
  DFF ram_reg_484__2_ ( .D(n16747), .CP(wclk), .Q(ram[12506]) );
  DFF ram_reg_484__1_ ( .D(n16746), .CP(wclk), .Q(ram[12505]) );
  DFF ram_reg_484__0_ ( .D(n16745), .CP(wclk), .Q(ram[12504]) );
  DFF ram_reg_500__7_ ( .D(n16624), .CP(wclk), .Q(ram[12383]) );
  DFF ram_reg_500__6_ ( .D(n16623), .CP(wclk), .Q(ram[12382]) );
  DFF ram_reg_500__5_ ( .D(n16622), .CP(wclk), .Q(ram[12381]) );
  DFF ram_reg_500__4_ ( .D(n16621), .CP(wclk), .Q(ram[12380]) );
  DFF ram_reg_500__3_ ( .D(n16620), .CP(wclk), .Q(ram[12379]) );
  DFF ram_reg_500__2_ ( .D(n16619), .CP(wclk), .Q(ram[12378]) );
  DFF ram_reg_500__1_ ( .D(n16618), .CP(wclk), .Q(ram[12377]) );
  DFF ram_reg_500__0_ ( .D(n16617), .CP(wclk), .Q(ram[12376]) );
  DFF ram_reg_512__7_ ( .D(n16528), .CP(wclk), .Q(ram[12287]) );
  DFF ram_reg_512__6_ ( .D(n16527), .CP(wclk), .Q(ram[12286]) );
  DFF ram_reg_512__5_ ( .D(n16526), .CP(wclk), .Q(ram[12285]) );
  DFF ram_reg_512__4_ ( .D(n16525), .CP(wclk), .Q(ram[12284]) );
  DFF ram_reg_512__3_ ( .D(n16524), .CP(wclk), .Q(ram[12283]) );
  DFF ram_reg_512__2_ ( .D(n16523), .CP(wclk), .Q(ram[12282]) );
  DFF ram_reg_512__1_ ( .D(n16522), .CP(wclk), .Q(ram[12281]) );
  DFF ram_reg_512__0_ ( .D(n16521), .CP(wclk), .Q(ram[12280]) );
  DFF ram_reg_516__7_ ( .D(n16496), .CP(wclk), .Q(ram[12255]) );
  DFF ram_reg_516__6_ ( .D(n16495), .CP(wclk), .Q(ram[12254]) );
  DFF ram_reg_516__5_ ( .D(n16494), .CP(wclk), .Q(ram[12253]) );
  DFF ram_reg_516__4_ ( .D(n16493), .CP(wclk), .Q(ram[12252]) );
  DFF ram_reg_516__3_ ( .D(n16492), .CP(wclk), .Q(ram[12251]) );
  DFF ram_reg_516__2_ ( .D(n16491), .CP(wclk), .Q(ram[12250]) );
  DFF ram_reg_516__1_ ( .D(n16490), .CP(wclk), .Q(ram[12249]) );
  DFF ram_reg_516__0_ ( .D(n16489), .CP(wclk), .Q(ram[12248]) );
  DFF ram_reg_524__7_ ( .D(n16432), .CP(wclk), .Q(ram[12191]) );
  DFF ram_reg_524__6_ ( .D(n16431), .CP(wclk), .Q(ram[12190]) );
  DFF ram_reg_524__5_ ( .D(n16430), .CP(wclk), .Q(ram[12189]) );
  DFF ram_reg_524__4_ ( .D(n16429), .CP(wclk), .Q(ram[12188]) );
  DFF ram_reg_524__3_ ( .D(n16428), .CP(wclk), .Q(ram[12187]) );
  DFF ram_reg_524__2_ ( .D(n16427), .CP(wclk), .Q(ram[12186]) );
  DFF ram_reg_524__1_ ( .D(n16426), .CP(wclk), .Q(ram[12185]) );
  DFF ram_reg_524__0_ ( .D(n16425), .CP(wclk), .Q(ram[12184]) );
  DFF ram_reg_528__7_ ( .D(n16400), .CP(wclk), .Q(ram[12159]) );
  DFF ram_reg_528__6_ ( .D(n16399), .CP(wclk), .Q(ram[12158]) );
  DFF ram_reg_528__5_ ( .D(n16398), .CP(wclk), .Q(ram[12157]) );
  DFF ram_reg_528__4_ ( .D(n16397), .CP(wclk), .Q(ram[12156]) );
  DFF ram_reg_528__3_ ( .D(n16396), .CP(wclk), .Q(ram[12155]) );
  DFF ram_reg_528__2_ ( .D(n16395), .CP(wclk), .Q(ram[12154]) );
  DFF ram_reg_528__1_ ( .D(n16394), .CP(wclk), .Q(ram[12153]) );
  DFF ram_reg_528__0_ ( .D(n16393), .CP(wclk), .Q(ram[12152]) );
  DFF ram_reg_532__7_ ( .D(n16368), .CP(wclk), .Q(ram[12127]) );
  DFF ram_reg_532__6_ ( .D(n16367), .CP(wclk), .Q(ram[12126]) );
  DFF ram_reg_532__5_ ( .D(n16366), .CP(wclk), .Q(ram[12125]) );
  DFF ram_reg_532__4_ ( .D(n16365), .CP(wclk), .Q(ram[12124]) );
  DFF ram_reg_532__3_ ( .D(n16364), .CP(wclk), .Q(ram[12123]) );
  DFF ram_reg_532__2_ ( .D(n16363), .CP(wclk), .Q(ram[12122]) );
  DFF ram_reg_532__1_ ( .D(n16362), .CP(wclk), .Q(ram[12121]) );
  DFF ram_reg_532__0_ ( .D(n16361), .CP(wclk), .Q(ram[12120]) );
  DFF ram_reg_540__7_ ( .D(n16304), .CP(wclk), .Q(ram[12063]) );
  DFF ram_reg_540__6_ ( .D(n16303), .CP(wclk), .Q(ram[12062]) );
  DFF ram_reg_540__5_ ( .D(n16302), .CP(wclk), .Q(ram[12061]) );
  DFF ram_reg_540__4_ ( .D(n16301), .CP(wclk), .Q(ram[12060]) );
  DFF ram_reg_540__3_ ( .D(n16300), .CP(wclk), .Q(ram[12059]) );
  DFF ram_reg_540__2_ ( .D(n16299), .CP(wclk), .Q(ram[12058]) );
  DFF ram_reg_540__1_ ( .D(n16298), .CP(wclk), .Q(ram[12057]) );
  DFF ram_reg_540__0_ ( .D(n16297), .CP(wclk), .Q(ram[12056]) );
  DFF ram_reg_544__7_ ( .D(n16272), .CP(wclk), .Q(ram[12031]) );
  DFF ram_reg_544__6_ ( .D(n16271), .CP(wclk), .Q(ram[12030]) );
  DFF ram_reg_544__5_ ( .D(n16270), .CP(wclk), .Q(ram[12029]) );
  DFF ram_reg_544__4_ ( .D(n16269), .CP(wclk), .Q(ram[12028]) );
  DFF ram_reg_544__3_ ( .D(n16268), .CP(wclk), .Q(ram[12027]) );
  DFF ram_reg_544__2_ ( .D(n16267), .CP(wclk), .Q(ram[12026]) );
  DFF ram_reg_544__1_ ( .D(n16266), .CP(wclk), .Q(ram[12025]) );
  DFF ram_reg_544__0_ ( .D(n16265), .CP(wclk), .Q(ram[12024]) );
  DFF ram_reg_548__7_ ( .D(n16240), .CP(wclk), .Q(ram[11999]) );
  DFF ram_reg_548__6_ ( .D(n16239), .CP(wclk), .Q(ram[11998]) );
  DFF ram_reg_548__5_ ( .D(n16238), .CP(wclk), .Q(ram[11997]) );
  DFF ram_reg_548__4_ ( .D(n16237), .CP(wclk), .Q(ram[11996]) );
  DFF ram_reg_548__3_ ( .D(n16236), .CP(wclk), .Q(ram[11995]) );
  DFF ram_reg_548__2_ ( .D(n16235), .CP(wclk), .Q(ram[11994]) );
  DFF ram_reg_548__1_ ( .D(n16234), .CP(wclk), .Q(ram[11993]) );
  DFF ram_reg_548__0_ ( .D(n16233), .CP(wclk), .Q(ram[11992]) );
  DFF ram_reg_560__7_ ( .D(n16144), .CP(wclk), .Q(ram[11903]) );
  DFF ram_reg_560__6_ ( .D(n16143), .CP(wclk), .Q(ram[11902]) );
  DFF ram_reg_560__5_ ( .D(n16142), .CP(wclk), .Q(ram[11901]) );
  DFF ram_reg_560__4_ ( .D(n16141), .CP(wclk), .Q(ram[11900]) );
  DFF ram_reg_560__3_ ( .D(n16140), .CP(wclk), .Q(ram[11899]) );
  DFF ram_reg_560__2_ ( .D(n16139), .CP(wclk), .Q(ram[11898]) );
  DFF ram_reg_560__1_ ( .D(n16138), .CP(wclk), .Q(ram[11897]) );
  DFF ram_reg_560__0_ ( .D(n16137), .CP(wclk), .Q(ram[11896]) );
  DFF ram_reg_564__7_ ( .D(n16112), .CP(wclk), .Q(ram[11871]) );
  DFF ram_reg_564__6_ ( .D(n16111), .CP(wclk), .Q(ram[11870]) );
  DFF ram_reg_564__5_ ( .D(n16110), .CP(wclk), .Q(ram[11869]) );
  DFF ram_reg_564__4_ ( .D(n16109), .CP(wclk), .Q(ram[11868]) );
  DFF ram_reg_564__3_ ( .D(n16108), .CP(wclk), .Q(ram[11867]) );
  DFF ram_reg_564__2_ ( .D(n16107), .CP(wclk), .Q(ram[11866]) );
  DFF ram_reg_564__1_ ( .D(n16106), .CP(wclk), .Q(ram[11865]) );
  DFF ram_reg_564__0_ ( .D(n16105), .CP(wclk), .Q(ram[11864]) );
  DFF ram_reg_576__7_ ( .D(n16016), .CP(wclk), .Q(ram[11775]) );
  DFF ram_reg_576__6_ ( .D(n16015), .CP(wclk), .Q(ram[11774]) );
  DFF ram_reg_576__5_ ( .D(n16014), .CP(wclk), .Q(ram[11773]) );
  DFF ram_reg_576__4_ ( .D(n16013), .CP(wclk), .Q(ram[11772]) );
  DFF ram_reg_576__3_ ( .D(n16012), .CP(wclk), .Q(ram[11771]) );
  DFF ram_reg_576__2_ ( .D(n16011), .CP(wclk), .Q(ram[11770]) );
  DFF ram_reg_576__1_ ( .D(n16010), .CP(wclk), .Q(ram[11769]) );
  DFF ram_reg_576__0_ ( .D(n16009), .CP(wclk), .Q(ram[11768]) );
  DFF ram_reg_580__7_ ( .D(n15984), .CP(wclk), .Q(ram[11743]) );
  DFF ram_reg_580__6_ ( .D(n15983), .CP(wclk), .Q(ram[11742]) );
  DFF ram_reg_580__5_ ( .D(n15982), .CP(wclk), .Q(ram[11741]) );
  DFF ram_reg_580__4_ ( .D(n15981), .CP(wclk), .Q(ram[11740]) );
  DFF ram_reg_580__3_ ( .D(n15980), .CP(wclk), .Q(ram[11739]) );
  DFF ram_reg_580__2_ ( .D(n15979), .CP(wclk), .Q(ram[11738]) );
  DFF ram_reg_580__1_ ( .D(n15978), .CP(wclk), .Q(ram[11737]) );
  DFF ram_reg_580__0_ ( .D(n15977), .CP(wclk), .Q(ram[11736]) );
  DFF ram_reg_584__7_ ( .D(n15952), .CP(wclk), .Q(ram[11711]) );
  DFF ram_reg_584__6_ ( .D(n15951), .CP(wclk), .Q(ram[11710]) );
  DFF ram_reg_584__5_ ( .D(n15950), .CP(wclk), .Q(ram[11709]) );
  DFF ram_reg_584__4_ ( .D(n15949), .CP(wclk), .Q(ram[11708]) );
  DFF ram_reg_584__3_ ( .D(n15948), .CP(wclk), .Q(ram[11707]) );
  DFF ram_reg_584__2_ ( .D(n15947), .CP(wclk), .Q(ram[11706]) );
  DFF ram_reg_584__1_ ( .D(n15946), .CP(wclk), .Q(ram[11705]) );
  DFF ram_reg_584__0_ ( .D(n15945), .CP(wclk), .Q(ram[11704]) );
  DFF ram_reg_588__7_ ( .D(n15920), .CP(wclk), .Q(ram[11679]) );
  DFF ram_reg_588__6_ ( .D(n15919), .CP(wclk), .Q(ram[11678]) );
  DFF ram_reg_588__5_ ( .D(n15918), .CP(wclk), .Q(ram[11677]) );
  DFF ram_reg_588__4_ ( .D(n15917), .CP(wclk), .Q(ram[11676]) );
  DFF ram_reg_588__3_ ( .D(n15916), .CP(wclk), .Q(ram[11675]) );
  DFF ram_reg_588__2_ ( .D(n15915), .CP(wclk), .Q(ram[11674]) );
  DFF ram_reg_588__1_ ( .D(n15914), .CP(wclk), .Q(ram[11673]) );
  DFF ram_reg_588__0_ ( .D(n15913), .CP(wclk), .Q(ram[11672]) );
  DFF ram_reg_592__7_ ( .D(n15888), .CP(wclk), .Q(ram[11647]) );
  DFF ram_reg_592__6_ ( .D(n15887), .CP(wclk), .Q(ram[11646]) );
  DFF ram_reg_592__5_ ( .D(n15886), .CP(wclk), .Q(ram[11645]) );
  DFF ram_reg_592__4_ ( .D(n15885), .CP(wclk), .Q(ram[11644]) );
  DFF ram_reg_592__3_ ( .D(n15884), .CP(wclk), .Q(ram[11643]) );
  DFF ram_reg_592__2_ ( .D(n15883), .CP(wclk), .Q(ram[11642]) );
  DFF ram_reg_592__1_ ( .D(n15882), .CP(wclk), .Q(ram[11641]) );
  DFF ram_reg_592__0_ ( .D(n15881), .CP(wclk), .Q(ram[11640]) );
  DFF ram_reg_596__7_ ( .D(n15856), .CP(wclk), .Q(ram[11615]) );
  DFF ram_reg_596__6_ ( .D(n15855), .CP(wclk), .Q(ram[11614]) );
  DFF ram_reg_596__5_ ( .D(n15854), .CP(wclk), .Q(ram[11613]) );
  DFF ram_reg_596__4_ ( .D(n15853), .CP(wclk), .Q(ram[11612]) );
  DFF ram_reg_596__3_ ( .D(n15852), .CP(wclk), .Q(ram[11611]) );
  DFF ram_reg_596__2_ ( .D(n15851), .CP(wclk), .Q(ram[11610]) );
  DFF ram_reg_596__1_ ( .D(n15850), .CP(wclk), .Q(ram[11609]) );
  DFF ram_reg_596__0_ ( .D(n15849), .CP(wclk), .Q(ram[11608]) );
  DFF ram_reg_600__7_ ( .D(n15824), .CP(wclk), .Q(ram[11583]) );
  DFF ram_reg_600__6_ ( .D(n15823), .CP(wclk), .Q(ram[11582]) );
  DFF ram_reg_600__5_ ( .D(n15822), .CP(wclk), .Q(ram[11581]) );
  DFF ram_reg_600__4_ ( .D(n15821), .CP(wclk), .Q(ram[11580]) );
  DFF ram_reg_600__3_ ( .D(n15820), .CP(wclk), .Q(ram[11579]) );
  DFF ram_reg_600__2_ ( .D(n15819), .CP(wclk), .Q(ram[11578]) );
  DFF ram_reg_600__1_ ( .D(n15818), .CP(wclk), .Q(ram[11577]) );
  DFF ram_reg_600__0_ ( .D(n15817), .CP(wclk), .Q(ram[11576]) );
  DFF ram_reg_604__7_ ( .D(n15792), .CP(wclk), .Q(ram[11551]) );
  DFF ram_reg_604__6_ ( .D(n15791), .CP(wclk), .Q(ram[11550]) );
  DFF ram_reg_604__5_ ( .D(n15790), .CP(wclk), .Q(ram[11549]) );
  DFF ram_reg_604__4_ ( .D(n15789), .CP(wclk), .Q(ram[11548]) );
  DFF ram_reg_604__3_ ( .D(n15788), .CP(wclk), .Q(ram[11547]) );
  DFF ram_reg_604__2_ ( .D(n15787), .CP(wclk), .Q(ram[11546]) );
  DFF ram_reg_604__1_ ( .D(n15786), .CP(wclk), .Q(ram[11545]) );
  DFF ram_reg_604__0_ ( .D(n15785), .CP(wclk), .Q(ram[11544]) );
  DFF ram_reg_608__7_ ( .D(n15760), .CP(wclk), .Q(ram[11519]) );
  DFF ram_reg_608__6_ ( .D(n15759), .CP(wclk), .Q(ram[11518]) );
  DFF ram_reg_608__5_ ( .D(n15758), .CP(wclk), .Q(ram[11517]) );
  DFF ram_reg_608__4_ ( .D(n15757), .CP(wclk), .Q(ram[11516]) );
  DFF ram_reg_608__3_ ( .D(n15756), .CP(wclk), .Q(ram[11515]) );
  DFF ram_reg_608__2_ ( .D(n15755), .CP(wclk), .Q(ram[11514]) );
  DFF ram_reg_608__1_ ( .D(n15754), .CP(wclk), .Q(ram[11513]) );
  DFF ram_reg_608__0_ ( .D(n15753), .CP(wclk), .Q(ram[11512]) );
  DFF ram_reg_612__7_ ( .D(n15728), .CP(wclk), .Q(ram[11487]) );
  DFF ram_reg_612__6_ ( .D(n15727), .CP(wclk), .Q(ram[11486]) );
  DFF ram_reg_612__5_ ( .D(n15726), .CP(wclk), .Q(ram[11485]) );
  DFF ram_reg_612__4_ ( .D(n15725), .CP(wclk), .Q(ram[11484]) );
  DFF ram_reg_612__3_ ( .D(n15724), .CP(wclk), .Q(ram[11483]) );
  DFF ram_reg_612__2_ ( .D(n15723), .CP(wclk), .Q(ram[11482]) );
  DFF ram_reg_612__1_ ( .D(n15722), .CP(wclk), .Q(ram[11481]) );
  DFF ram_reg_612__0_ ( .D(n15721), .CP(wclk), .Q(ram[11480]) );
  DFF ram_reg_616__7_ ( .D(n15696), .CP(wclk), .Q(ram[11455]) );
  DFF ram_reg_616__6_ ( .D(n15695), .CP(wclk), .Q(ram[11454]) );
  DFF ram_reg_616__5_ ( .D(n15694), .CP(wclk), .Q(ram[11453]) );
  DFF ram_reg_616__4_ ( .D(n15693), .CP(wclk), .Q(ram[11452]) );
  DFF ram_reg_616__3_ ( .D(n15692), .CP(wclk), .Q(ram[11451]) );
  DFF ram_reg_616__2_ ( .D(n15691), .CP(wclk), .Q(ram[11450]) );
  DFF ram_reg_616__1_ ( .D(n15690), .CP(wclk), .Q(ram[11449]) );
  DFF ram_reg_616__0_ ( .D(n15689), .CP(wclk), .Q(ram[11448]) );
  DFF ram_reg_620__7_ ( .D(n15664), .CP(wclk), .Q(ram[11423]) );
  DFF ram_reg_620__6_ ( .D(n15663), .CP(wclk), .Q(ram[11422]) );
  DFF ram_reg_620__5_ ( .D(n15662), .CP(wclk), .Q(ram[11421]) );
  DFF ram_reg_620__4_ ( .D(n15661), .CP(wclk), .Q(ram[11420]) );
  DFF ram_reg_620__3_ ( .D(n15660), .CP(wclk), .Q(ram[11419]) );
  DFF ram_reg_620__2_ ( .D(n15659), .CP(wclk), .Q(ram[11418]) );
  DFF ram_reg_620__1_ ( .D(n15658), .CP(wclk), .Q(ram[11417]) );
  DFF ram_reg_620__0_ ( .D(n15657), .CP(wclk), .Q(ram[11416]) );
  DFF ram_reg_624__7_ ( .D(n15632), .CP(wclk), .Q(ram[11391]) );
  DFF ram_reg_624__6_ ( .D(n15631), .CP(wclk), .Q(ram[11390]) );
  DFF ram_reg_624__5_ ( .D(n15630), .CP(wclk), .Q(ram[11389]) );
  DFF ram_reg_624__4_ ( .D(n15629), .CP(wclk), .Q(ram[11388]) );
  DFF ram_reg_624__3_ ( .D(n15628), .CP(wclk), .Q(ram[11387]) );
  DFF ram_reg_624__2_ ( .D(n15627), .CP(wclk), .Q(ram[11386]) );
  DFF ram_reg_624__1_ ( .D(n15626), .CP(wclk), .Q(ram[11385]) );
  DFF ram_reg_624__0_ ( .D(n15625), .CP(wclk), .Q(ram[11384]) );
  DFF ram_reg_628__7_ ( .D(n15600), .CP(wclk), .Q(ram[11359]) );
  DFF ram_reg_628__6_ ( .D(n15599), .CP(wclk), .Q(ram[11358]) );
  DFF ram_reg_628__5_ ( .D(n15598), .CP(wclk), .Q(ram[11357]) );
  DFF ram_reg_628__4_ ( .D(n15597), .CP(wclk), .Q(ram[11356]) );
  DFF ram_reg_628__3_ ( .D(n15596), .CP(wclk), .Q(ram[11355]) );
  DFF ram_reg_628__2_ ( .D(n15595), .CP(wclk), .Q(ram[11354]) );
  DFF ram_reg_628__1_ ( .D(n15594), .CP(wclk), .Q(ram[11353]) );
  DFF ram_reg_628__0_ ( .D(n15593), .CP(wclk), .Q(ram[11352]) );
  DFF ram_reg_636__7_ ( .D(n15536), .CP(wclk), .Q(ram[11295]) );
  DFF ram_reg_636__6_ ( .D(n15535), .CP(wclk), .Q(ram[11294]) );
  DFF ram_reg_636__5_ ( .D(n15534), .CP(wclk), .Q(ram[11293]) );
  DFF ram_reg_636__4_ ( .D(n15533), .CP(wclk), .Q(ram[11292]) );
  DFF ram_reg_636__3_ ( .D(n15532), .CP(wclk), .Q(ram[11291]) );
  DFF ram_reg_636__2_ ( .D(n15531), .CP(wclk), .Q(ram[11290]) );
  DFF ram_reg_636__1_ ( .D(n15530), .CP(wclk), .Q(ram[11289]) );
  DFF ram_reg_636__0_ ( .D(n15529), .CP(wclk), .Q(ram[11288]) );
  DFF ram_reg_644__7_ ( .D(n15472), .CP(wclk), .Q(ram[11231]) );
  DFF ram_reg_644__6_ ( .D(n15471), .CP(wclk), .Q(ram[11230]) );
  DFF ram_reg_644__5_ ( .D(n15470), .CP(wclk), .Q(ram[11229]) );
  DFF ram_reg_644__4_ ( .D(n15469), .CP(wclk), .Q(ram[11228]) );
  DFF ram_reg_644__3_ ( .D(n15468), .CP(wclk), .Q(ram[11227]) );
  DFF ram_reg_644__2_ ( .D(n15467), .CP(wclk), .Q(ram[11226]) );
  DFF ram_reg_644__1_ ( .D(n15466), .CP(wclk), .Q(ram[11225]) );
  DFF ram_reg_644__0_ ( .D(n15465), .CP(wclk), .Q(ram[11224]) );
  DFF ram_reg_660__7_ ( .D(n15344), .CP(wclk), .Q(ram[11103]) );
  DFF ram_reg_660__6_ ( .D(n15343), .CP(wclk), .Q(ram[11102]) );
  DFF ram_reg_660__5_ ( .D(n15342), .CP(wclk), .Q(ram[11101]) );
  DFF ram_reg_660__4_ ( .D(n15341), .CP(wclk), .Q(ram[11100]) );
  DFF ram_reg_660__3_ ( .D(n15340), .CP(wclk), .Q(ram[11099]) );
  DFF ram_reg_660__2_ ( .D(n15339), .CP(wclk), .Q(ram[11098]) );
  DFF ram_reg_660__1_ ( .D(n15338), .CP(wclk), .Q(ram[11097]) );
  DFF ram_reg_660__0_ ( .D(n15337), .CP(wclk), .Q(ram[11096]) );
  DFF ram_reg_676__7_ ( .D(n15216), .CP(wclk), .Q(ram[10975]) );
  DFF ram_reg_676__6_ ( .D(n15215), .CP(wclk), .Q(ram[10974]) );
  DFF ram_reg_676__5_ ( .D(n15214), .CP(wclk), .Q(ram[10973]) );
  DFF ram_reg_676__4_ ( .D(n15213), .CP(wclk), .Q(ram[10972]) );
  DFF ram_reg_676__3_ ( .D(n15212), .CP(wclk), .Q(ram[10971]) );
  DFF ram_reg_676__2_ ( .D(n15211), .CP(wclk), .Q(ram[10970]) );
  DFF ram_reg_676__1_ ( .D(n15210), .CP(wclk), .Q(ram[10969]) );
  DFF ram_reg_676__0_ ( .D(n15209), .CP(wclk), .Q(ram[10968]) );
  DFF ram_reg_704__7_ ( .D(n14992), .CP(wclk), .Q(ram[10751]) );
  DFF ram_reg_704__6_ ( .D(n14991), .CP(wclk), .Q(ram[10750]) );
  DFF ram_reg_704__5_ ( .D(n14990), .CP(wclk), .Q(ram[10749]) );
  DFF ram_reg_704__4_ ( .D(n14989), .CP(wclk), .Q(ram[10748]) );
  DFF ram_reg_704__3_ ( .D(n14988), .CP(wclk), .Q(ram[10747]) );
  DFF ram_reg_704__2_ ( .D(n14987), .CP(wclk), .Q(ram[10746]) );
  DFF ram_reg_704__1_ ( .D(n14986), .CP(wclk), .Q(ram[10745]) );
  DFF ram_reg_704__0_ ( .D(n14985), .CP(wclk), .Q(ram[10744]) );
  DFF ram_reg_708__7_ ( .D(n14960), .CP(wclk), .Q(ram[10719]) );
  DFF ram_reg_708__6_ ( .D(n14959), .CP(wclk), .Q(ram[10718]) );
  DFF ram_reg_708__5_ ( .D(n14958), .CP(wclk), .Q(ram[10717]) );
  DFF ram_reg_708__4_ ( .D(n14957), .CP(wclk), .Q(ram[10716]) );
  DFF ram_reg_708__3_ ( .D(n14956), .CP(wclk), .Q(ram[10715]) );
  DFF ram_reg_708__2_ ( .D(n14955), .CP(wclk), .Q(ram[10714]) );
  DFF ram_reg_708__1_ ( .D(n14954), .CP(wclk), .Q(ram[10713]) );
  DFF ram_reg_708__0_ ( .D(n14953), .CP(wclk), .Q(ram[10712]) );
  DFF ram_reg_720__7_ ( .D(n14864), .CP(wclk), .Q(ram[10623]) );
  DFF ram_reg_720__6_ ( .D(n14863), .CP(wclk), .Q(ram[10622]) );
  DFF ram_reg_720__5_ ( .D(n14862), .CP(wclk), .Q(ram[10621]) );
  DFF ram_reg_720__4_ ( .D(n14861), .CP(wclk), .Q(ram[10620]) );
  DFF ram_reg_720__3_ ( .D(n14860), .CP(wclk), .Q(ram[10619]) );
  DFF ram_reg_720__2_ ( .D(n14859), .CP(wclk), .Q(ram[10618]) );
  DFF ram_reg_720__1_ ( .D(n14858), .CP(wclk), .Q(ram[10617]) );
  DFF ram_reg_720__0_ ( .D(n14857), .CP(wclk), .Q(ram[10616]) );
  DFF ram_reg_724__7_ ( .D(n14832), .CP(wclk), .Q(ram[10591]) );
  DFF ram_reg_724__6_ ( .D(n14831), .CP(wclk), .Q(ram[10590]) );
  DFF ram_reg_724__5_ ( .D(n14830), .CP(wclk), .Q(ram[10589]) );
  DFF ram_reg_724__4_ ( .D(n14829), .CP(wclk), .Q(ram[10588]) );
  DFF ram_reg_724__3_ ( .D(n14828), .CP(wclk), .Q(ram[10587]) );
  DFF ram_reg_724__2_ ( .D(n14827), .CP(wclk), .Q(ram[10586]) );
  DFF ram_reg_724__1_ ( .D(n14826), .CP(wclk), .Q(ram[10585]) );
  DFF ram_reg_724__0_ ( .D(n14825), .CP(wclk), .Q(ram[10584]) );
  DFF ram_reg_740__7_ ( .D(n14704), .CP(wclk), .Q(ram[10463]) );
  DFF ram_reg_740__6_ ( .D(n14703), .CP(wclk), .Q(ram[10462]) );
  DFF ram_reg_740__5_ ( .D(n14702), .CP(wclk), .Q(ram[10461]) );
  DFF ram_reg_740__4_ ( .D(n14701), .CP(wclk), .Q(ram[10460]) );
  DFF ram_reg_740__3_ ( .D(n14700), .CP(wclk), .Q(ram[10459]) );
  DFF ram_reg_740__2_ ( .D(n14699), .CP(wclk), .Q(ram[10458]) );
  DFF ram_reg_740__1_ ( .D(n14698), .CP(wclk), .Q(ram[10457]) );
  DFF ram_reg_740__0_ ( .D(n14697), .CP(wclk), .Q(ram[10456]) );
  DFF ram_reg_756__7_ ( .D(n14576), .CP(wclk), .Q(ram[10335]) );
  DFF ram_reg_756__6_ ( .D(n14575), .CP(wclk), .Q(ram[10334]) );
  DFF ram_reg_756__5_ ( .D(n14574), .CP(wclk), .Q(ram[10333]) );
  DFF ram_reg_756__4_ ( .D(n14573), .CP(wclk), .Q(ram[10332]) );
  DFF ram_reg_756__3_ ( .D(n14572), .CP(wclk), .Q(ram[10331]) );
  DFF ram_reg_756__2_ ( .D(n14571), .CP(wclk), .Q(ram[10330]) );
  DFF ram_reg_756__1_ ( .D(n14570), .CP(wclk), .Q(ram[10329]) );
  DFF ram_reg_756__0_ ( .D(n14569), .CP(wclk), .Q(ram[10328]) );
  DFF ram_reg_768__7_ ( .D(n14480), .CP(wclk), .Q(ram[10239]) );
  DFF ram_reg_768__6_ ( .D(n14479), .CP(wclk), .Q(ram[10238]) );
  DFF ram_reg_768__5_ ( .D(n14478), .CP(wclk), .Q(ram[10237]) );
  DFF ram_reg_768__4_ ( .D(n14477), .CP(wclk), .Q(ram[10236]) );
  DFF ram_reg_768__3_ ( .D(n14476), .CP(wclk), .Q(ram[10235]) );
  DFF ram_reg_768__2_ ( .D(n14475), .CP(wclk), .Q(ram[10234]) );
  DFF ram_reg_768__1_ ( .D(n14474), .CP(wclk), .Q(ram[10233]) );
  DFF ram_reg_768__0_ ( .D(n14473), .CP(wclk), .Q(ram[10232]) );
  DFF ram_reg_772__7_ ( .D(n14448), .CP(wclk), .Q(ram[10207]) );
  DFF ram_reg_772__6_ ( .D(n14447), .CP(wclk), .Q(ram[10206]) );
  DFF ram_reg_772__5_ ( .D(n14446), .CP(wclk), .Q(ram[10205]) );
  DFF ram_reg_772__4_ ( .D(n14445), .CP(wclk), .Q(ram[10204]) );
  DFF ram_reg_772__3_ ( .D(n14444), .CP(wclk), .Q(ram[10203]) );
  DFF ram_reg_772__2_ ( .D(n14443), .CP(wclk), .Q(ram[10202]) );
  DFF ram_reg_772__1_ ( .D(n14442), .CP(wclk), .Q(ram[10201]) );
  DFF ram_reg_772__0_ ( .D(n14441), .CP(wclk), .Q(ram[10200]) );
  DFF ram_reg_784__7_ ( .D(n14352), .CP(wclk), .Q(ram[10111]) );
  DFF ram_reg_784__6_ ( .D(n14351), .CP(wclk), .Q(ram[10110]) );
  DFF ram_reg_784__5_ ( .D(n14350), .CP(wclk), .Q(ram[10109]) );
  DFF ram_reg_784__4_ ( .D(n14349), .CP(wclk), .Q(ram[10108]) );
  DFF ram_reg_784__3_ ( .D(n14348), .CP(wclk), .Q(ram[10107]) );
  DFF ram_reg_784__2_ ( .D(n14347), .CP(wclk), .Q(ram[10106]) );
  DFF ram_reg_784__1_ ( .D(n14346), .CP(wclk), .Q(ram[10105]) );
  DFF ram_reg_784__0_ ( .D(n14345), .CP(wclk), .Q(ram[10104]) );
  DFF ram_reg_788__7_ ( .D(n14320), .CP(wclk), .Q(ram[10079]) );
  DFF ram_reg_788__6_ ( .D(n14319), .CP(wclk), .Q(ram[10078]) );
  DFF ram_reg_788__5_ ( .D(n14318), .CP(wclk), .Q(ram[10077]) );
  DFF ram_reg_788__4_ ( .D(n14317), .CP(wclk), .Q(ram[10076]) );
  DFF ram_reg_788__3_ ( .D(n14316), .CP(wclk), .Q(ram[10075]) );
  DFF ram_reg_788__2_ ( .D(n14315), .CP(wclk), .Q(ram[10074]) );
  DFF ram_reg_788__1_ ( .D(n14314), .CP(wclk), .Q(ram[10073]) );
  DFF ram_reg_788__0_ ( .D(n14313), .CP(wclk), .Q(ram[10072]) );
  DFF ram_reg_796__7_ ( .D(n14256), .CP(wclk), .Q(ram[10015]) );
  DFF ram_reg_796__6_ ( .D(n14255), .CP(wclk), .Q(ram[10014]) );
  DFF ram_reg_796__5_ ( .D(n14254), .CP(wclk), .Q(ram[10013]) );
  DFF ram_reg_796__4_ ( .D(n14253), .CP(wclk), .Q(ram[10012]) );
  DFF ram_reg_796__3_ ( .D(n14252), .CP(wclk), .Q(ram[10011]) );
  DFF ram_reg_796__2_ ( .D(n14251), .CP(wclk), .Q(ram[10010]) );
  DFF ram_reg_796__1_ ( .D(n14250), .CP(wclk), .Q(ram[10009]) );
  DFF ram_reg_796__0_ ( .D(n14249), .CP(wclk), .Q(ram[10008]) );
  DFF ram_reg_800__7_ ( .D(n14224), .CP(wclk), .Q(ram[9983]) );
  DFF ram_reg_800__6_ ( .D(n14223), .CP(wclk), .Q(ram[9982]) );
  DFF ram_reg_800__5_ ( .D(n14222), .CP(wclk), .Q(ram[9981]) );
  DFF ram_reg_800__4_ ( .D(n14221), .CP(wclk), .Q(ram[9980]) );
  DFF ram_reg_800__3_ ( .D(n14220), .CP(wclk), .Q(ram[9979]) );
  DFF ram_reg_800__2_ ( .D(n14219), .CP(wclk), .Q(ram[9978]) );
  DFF ram_reg_800__1_ ( .D(n14218), .CP(wclk), .Q(ram[9977]) );
  DFF ram_reg_800__0_ ( .D(n14217), .CP(wclk), .Q(ram[9976]) );
  DFF ram_reg_804__7_ ( .D(n14192), .CP(wclk), .Q(ram[9951]) );
  DFF ram_reg_804__6_ ( .D(n14191), .CP(wclk), .Q(ram[9950]) );
  DFF ram_reg_804__5_ ( .D(n14190), .CP(wclk), .Q(ram[9949]) );
  DFF ram_reg_804__4_ ( .D(n14189), .CP(wclk), .Q(ram[9948]) );
  DFF ram_reg_804__3_ ( .D(n14188), .CP(wclk), .Q(ram[9947]) );
  DFF ram_reg_804__2_ ( .D(n14187), .CP(wclk), .Q(ram[9946]) );
  DFF ram_reg_804__1_ ( .D(n14186), .CP(wclk), .Q(ram[9945]) );
  DFF ram_reg_804__0_ ( .D(n14185), .CP(wclk), .Q(ram[9944]) );
  DFF ram_reg_820__7_ ( .D(n14064), .CP(wclk), .Q(ram[9823]) );
  DFF ram_reg_820__6_ ( .D(n14063), .CP(wclk), .Q(ram[9822]) );
  DFF ram_reg_820__5_ ( .D(n14062), .CP(wclk), .Q(ram[9821]) );
  DFF ram_reg_820__4_ ( .D(n14061), .CP(wclk), .Q(ram[9820]) );
  DFF ram_reg_820__3_ ( .D(n14060), .CP(wclk), .Q(ram[9819]) );
  DFF ram_reg_820__2_ ( .D(n14059), .CP(wclk), .Q(ram[9818]) );
  DFF ram_reg_820__1_ ( .D(n14058), .CP(wclk), .Q(ram[9817]) );
  DFF ram_reg_820__0_ ( .D(n14057), .CP(wclk), .Q(ram[9816]) );
  DFF ram_reg_832__7_ ( .D(n13968), .CP(wclk), .Q(ram[9727]) );
  DFF ram_reg_832__6_ ( .D(n13967), .CP(wclk), .Q(ram[9726]) );
  DFF ram_reg_832__5_ ( .D(n13966), .CP(wclk), .Q(ram[9725]) );
  DFF ram_reg_832__4_ ( .D(n13965), .CP(wclk), .Q(ram[9724]) );
  DFF ram_reg_832__3_ ( .D(n13964), .CP(wclk), .Q(ram[9723]) );
  DFF ram_reg_832__2_ ( .D(n13963), .CP(wclk), .Q(ram[9722]) );
  DFF ram_reg_832__1_ ( .D(n13962), .CP(wclk), .Q(ram[9721]) );
  DFF ram_reg_832__0_ ( .D(n13961), .CP(wclk), .Q(ram[9720]) );
  DFF ram_reg_836__7_ ( .D(n13936), .CP(wclk), .Q(ram[9695]) );
  DFF ram_reg_836__6_ ( .D(n13935), .CP(wclk), .Q(ram[9694]) );
  DFF ram_reg_836__5_ ( .D(n13934), .CP(wclk), .Q(ram[9693]) );
  DFF ram_reg_836__4_ ( .D(n13933), .CP(wclk), .Q(ram[9692]) );
  DFF ram_reg_836__3_ ( .D(n13932), .CP(wclk), .Q(ram[9691]) );
  DFF ram_reg_836__2_ ( .D(n13931), .CP(wclk), .Q(ram[9690]) );
  DFF ram_reg_836__1_ ( .D(n13930), .CP(wclk), .Q(ram[9689]) );
  DFF ram_reg_836__0_ ( .D(n13929), .CP(wclk), .Q(ram[9688]) );
  DFF ram_reg_840__7_ ( .D(n13904), .CP(wclk), .Q(ram[9663]) );
  DFF ram_reg_840__6_ ( .D(n13903), .CP(wclk), .Q(ram[9662]) );
  DFF ram_reg_840__5_ ( .D(n13902), .CP(wclk), .Q(ram[9661]) );
  DFF ram_reg_840__4_ ( .D(n13901), .CP(wclk), .Q(ram[9660]) );
  DFF ram_reg_840__3_ ( .D(n13900), .CP(wclk), .Q(ram[9659]) );
  DFF ram_reg_840__2_ ( .D(n13899), .CP(wclk), .Q(ram[9658]) );
  DFF ram_reg_840__1_ ( .D(n13898), .CP(wclk), .Q(ram[9657]) );
  DFF ram_reg_840__0_ ( .D(n13897), .CP(wclk), .Q(ram[9656]) );
  DFF ram_reg_844__7_ ( .D(n13872), .CP(wclk), .Q(ram[9631]) );
  DFF ram_reg_844__6_ ( .D(n13871), .CP(wclk), .Q(ram[9630]) );
  DFF ram_reg_844__5_ ( .D(n13870), .CP(wclk), .Q(ram[9629]) );
  DFF ram_reg_844__4_ ( .D(n13869), .CP(wclk), .Q(ram[9628]) );
  DFF ram_reg_844__3_ ( .D(n13868), .CP(wclk), .Q(ram[9627]) );
  DFF ram_reg_844__2_ ( .D(n13867), .CP(wclk), .Q(ram[9626]) );
  DFF ram_reg_844__1_ ( .D(n13866), .CP(wclk), .Q(ram[9625]) );
  DFF ram_reg_844__0_ ( .D(n13865), .CP(wclk), .Q(ram[9624]) );
  DFF ram_reg_848__7_ ( .D(n13840), .CP(wclk), .Q(ram[9599]) );
  DFF ram_reg_848__6_ ( .D(n13839), .CP(wclk), .Q(ram[9598]) );
  DFF ram_reg_848__5_ ( .D(n13838), .CP(wclk), .Q(ram[9597]) );
  DFF ram_reg_848__4_ ( .D(n13837), .CP(wclk), .Q(ram[9596]) );
  DFF ram_reg_848__3_ ( .D(n13836), .CP(wclk), .Q(ram[9595]) );
  DFF ram_reg_848__2_ ( .D(n13835), .CP(wclk), .Q(ram[9594]) );
  DFF ram_reg_848__1_ ( .D(n13834), .CP(wclk), .Q(ram[9593]) );
  DFF ram_reg_848__0_ ( .D(n13833), .CP(wclk), .Q(ram[9592]) );
  DFF ram_reg_852__7_ ( .D(n13808), .CP(wclk), .Q(ram[9567]) );
  DFF ram_reg_852__6_ ( .D(n13807), .CP(wclk), .Q(ram[9566]) );
  DFF ram_reg_852__5_ ( .D(n13806), .CP(wclk), .Q(ram[9565]) );
  DFF ram_reg_852__4_ ( .D(n13805), .CP(wclk), .Q(ram[9564]) );
  DFF ram_reg_852__3_ ( .D(n13804), .CP(wclk), .Q(ram[9563]) );
  DFF ram_reg_852__2_ ( .D(n13803), .CP(wclk), .Q(ram[9562]) );
  DFF ram_reg_852__1_ ( .D(n13802), .CP(wclk), .Q(ram[9561]) );
  DFF ram_reg_852__0_ ( .D(n13801), .CP(wclk), .Q(ram[9560]) );
  DFF ram_reg_856__7_ ( .D(n13776), .CP(wclk), .Q(ram[9535]) );
  DFF ram_reg_856__6_ ( .D(n13775), .CP(wclk), .Q(ram[9534]) );
  DFF ram_reg_856__5_ ( .D(n13774), .CP(wclk), .Q(ram[9533]) );
  DFF ram_reg_856__4_ ( .D(n13773), .CP(wclk), .Q(ram[9532]) );
  DFF ram_reg_856__3_ ( .D(n13772), .CP(wclk), .Q(ram[9531]) );
  DFF ram_reg_856__2_ ( .D(n13771), .CP(wclk), .Q(ram[9530]) );
  DFF ram_reg_856__1_ ( .D(n13770), .CP(wclk), .Q(ram[9529]) );
  DFF ram_reg_856__0_ ( .D(n13769), .CP(wclk), .Q(ram[9528]) );
  DFF ram_reg_860__7_ ( .D(n13744), .CP(wclk), .Q(ram[9503]) );
  DFF ram_reg_860__6_ ( .D(n13743), .CP(wclk), .Q(ram[9502]) );
  DFF ram_reg_860__5_ ( .D(n13742), .CP(wclk), .Q(ram[9501]) );
  DFF ram_reg_860__4_ ( .D(n13741), .CP(wclk), .Q(ram[9500]) );
  DFF ram_reg_860__3_ ( .D(n13740), .CP(wclk), .Q(ram[9499]) );
  DFF ram_reg_860__2_ ( .D(n13739), .CP(wclk), .Q(ram[9498]) );
  DFF ram_reg_860__1_ ( .D(n13738), .CP(wclk), .Q(ram[9497]) );
  DFF ram_reg_860__0_ ( .D(n13737), .CP(wclk), .Q(ram[9496]) );
  DFF ram_reg_864__7_ ( .D(n13712), .CP(wclk), .Q(ram[9471]) );
  DFF ram_reg_864__6_ ( .D(n13711), .CP(wclk), .Q(ram[9470]) );
  DFF ram_reg_864__5_ ( .D(n13710), .CP(wclk), .Q(ram[9469]) );
  DFF ram_reg_864__4_ ( .D(n13709), .CP(wclk), .Q(ram[9468]) );
  DFF ram_reg_864__3_ ( .D(n13708), .CP(wclk), .Q(ram[9467]) );
  DFF ram_reg_864__2_ ( .D(n13707), .CP(wclk), .Q(ram[9466]) );
  DFF ram_reg_864__1_ ( .D(n13706), .CP(wclk), .Q(ram[9465]) );
  DFF ram_reg_864__0_ ( .D(n13705), .CP(wclk), .Q(ram[9464]) );
  DFF ram_reg_868__7_ ( .D(n13680), .CP(wclk), .Q(ram[9439]) );
  DFF ram_reg_868__6_ ( .D(n13679), .CP(wclk), .Q(ram[9438]) );
  DFF ram_reg_868__5_ ( .D(n13678), .CP(wclk), .Q(ram[9437]) );
  DFF ram_reg_868__4_ ( .D(n13677), .CP(wclk), .Q(ram[9436]) );
  DFF ram_reg_868__3_ ( .D(n13676), .CP(wclk), .Q(ram[9435]) );
  DFF ram_reg_868__2_ ( .D(n13675), .CP(wclk), .Q(ram[9434]) );
  DFF ram_reg_868__1_ ( .D(n13674), .CP(wclk), .Q(ram[9433]) );
  DFF ram_reg_868__0_ ( .D(n13673), .CP(wclk), .Q(ram[9432]) );
  DFF ram_reg_876__7_ ( .D(n13616), .CP(wclk), .Q(ram[9375]) );
  DFF ram_reg_876__6_ ( .D(n13615), .CP(wclk), .Q(ram[9374]) );
  DFF ram_reg_876__5_ ( .D(n13614), .CP(wclk), .Q(ram[9373]) );
  DFF ram_reg_876__4_ ( .D(n13613), .CP(wclk), .Q(ram[9372]) );
  DFF ram_reg_876__3_ ( .D(n13612), .CP(wclk), .Q(ram[9371]) );
  DFF ram_reg_876__2_ ( .D(n13611), .CP(wclk), .Q(ram[9370]) );
  DFF ram_reg_876__1_ ( .D(n13610), .CP(wclk), .Q(ram[9369]) );
  DFF ram_reg_876__0_ ( .D(n13609), .CP(wclk), .Q(ram[9368]) );
  DFF ram_reg_880__7_ ( .D(n13584), .CP(wclk), .Q(ram[9343]) );
  DFF ram_reg_880__6_ ( .D(n13583), .CP(wclk), .Q(ram[9342]) );
  DFF ram_reg_880__5_ ( .D(n13582), .CP(wclk), .Q(ram[9341]) );
  DFF ram_reg_880__4_ ( .D(n13581), .CP(wclk), .Q(ram[9340]) );
  DFF ram_reg_880__3_ ( .D(n13580), .CP(wclk), .Q(ram[9339]) );
  DFF ram_reg_880__2_ ( .D(n13579), .CP(wclk), .Q(ram[9338]) );
  DFF ram_reg_880__1_ ( .D(n13578), .CP(wclk), .Q(ram[9337]) );
  DFF ram_reg_880__0_ ( .D(n13577), .CP(wclk), .Q(ram[9336]) );
  DFF ram_reg_884__7_ ( .D(n13552), .CP(wclk), .Q(ram[9311]) );
  DFF ram_reg_884__6_ ( .D(n13551), .CP(wclk), .Q(ram[9310]) );
  DFF ram_reg_884__5_ ( .D(n13550), .CP(wclk), .Q(ram[9309]) );
  DFF ram_reg_884__4_ ( .D(n13549), .CP(wclk), .Q(ram[9308]) );
  DFF ram_reg_884__3_ ( .D(n13548), .CP(wclk), .Q(ram[9307]) );
  DFF ram_reg_884__2_ ( .D(n13547), .CP(wclk), .Q(ram[9306]) );
  DFF ram_reg_884__1_ ( .D(n13546), .CP(wclk), .Q(ram[9305]) );
  DFF ram_reg_884__0_ ( .D(n13545), .CP(wclk), .Q(ram[9304]) );
  DFF ram_reg_892__7_ ( .D(n13488), .CP(wclk), .Q(ram[9247]) );
  DFF ram_reg_892__6_ ( .D(n13487), .CP(wclk), .Q(ram[9246]) );
  DFF ram_reg_892__5_ ( .D(n13486), .CP(wclk), .Q(ram[9245]) );
  DFF ram_reg_892__4_ ( .D(n13485), .CP(wclk), .Q(ram[9244]) );
  DFF ram_reg_892__3_ ( .D(n13484), .CP(wclk), .Q(ram[9243]) );
  DFF ram_reg_892__2_ ( .D(n13483), .CP(wclk), .Q(ram[9242]) );
  DFF ram_reg_892__1_ ( .D(n13482), .CP(wclk), .Q(ram[9241]) );
  DFF ram_reg_892__0_ ( .D(n13481), .CP(wclk), .Q(ram[9240]) );
  DFF ram_reg_900__7_ ( .D(n13424), .CP(wclk), .Q(ram[9183]) );
  DFF ram_reg_900__6_ ( .D(n13423), .CP(wclk), .Q(ram[9182]) );
  DFF ram_reg_900__5_ ( .D(n13422), .CP(wclk), .Q(ram[9181]) );
  DFF ram_reg_900__4_ ( .D(n13421), .CP(wclk), .Q(ram[9180]) );
  DFF ram_reg_900__3_ ( .D(n13420), .CP(wclk), .Q(ram[9179]) );
  DFF ram_reg_900__2_ ( .D(n13419), .CP(wclk), .Q(ram[9178]) );
  DFF ram_reg_900__1_ ( .D(n13418), .CP(wclk), .Q(ram[9177]) );
  DFF ram_reg_900__0_ ( .D(n13417), .CP(wclk), .Q(ram[9176]) );
  DFF ram_reg_916__7_ ( .D(n13296), .CP(wclk), .Q(ram[9055]) );
  DFF ram_reg_916__6_ ( .D(n13295), .CP(wclk), .Q(ram[9054]) );
  DFF ram_reg_916__5_ ( .D(n13294), .CP(wclk), .Q(ram[9053]) );
  DFF ram_reg_916__4_ ( .D(n13293), .CP(wclk), .Q(ram[9052]) );
  DFF ram_reg_916__3_ ( .D(n13292), .CP(wclk), .Q(ram[9051]) );
  DFF ram_reg_916__2_ ( .D(n13291), .CP(wclk), .Q(ram[9050]) );
  DFF ram_reg_916__1_ ( .D(n13290), .CP(wclk), .Q(ram[9049]) );
  DFF ram_reg_916__0_ ( .D(n13289), .CP(wclk), .Q(ram[9048]) );
  DFF ram_reg_964__7_ ( .D(n12912), .CP(wclk), .Q(ram[8671]) );
  DFF ram_reg_964__6_ ( .D(n12911), .CP(wclk), .Q(ram[8670]) );
  DFF ram_reg_964__5_ ( .D(n12910), .CP(wclk), .Q(ram[8669]) );
  DFF ram_reg_964__4_ ( .D(n12909), .CP(wclk), .Q(ram[8668]) );
  DFF ram_reg_964__3_ ( .D(n12908), .CP(wclk), .Q(ram[8667]) );
  DFF ram_reg_964__2_ ( .D(n12907), .CP(wclk), .Q(ram[8666]) );
  DFF ram_reg_964__1_ ( .D(n12906), .CP(wclk), .Q(ram[8665]) );
  DFF ram_reg_964__0_ ( .D(n12905), .CP(wclk), .Q(ram[8664]) );
  DFF ram_reg_976__7_ ( .D(n12816), .CP(wclk), .Q(ram[8575]) );
  DFF ram_reg_976__6_ ( .D(n12815), .CP(wclk), .Q(ram[8574]) );
  DFF ram_reg_976__5_ ( .D(n12814), .CP(wclk), .Q(ram[8573]) );
  DFF ram_reg_976__4_ ( .D(n12813), .CP(wclk), .Q(ram[8572]) );
  DFF ram_reg_976__3_ ( .D(n12812), .CP(wclk), .Q(ram[8571]) );
  DFF ram_reg_976__2_ ( .D(n12811), .CP(wclk), .Q(ram[8570]) );
  DFF ram_reg_976__1_ ( .D(n12810), .CP(wclk), .Q(ram[8569]) );
  DFF ram_reg_976__0_ ( .D(n12809), .CP(wclk), .Q(ram[8568]) );
  DFF ram_reg_980__7_ ( .D(n12784), .CP(wclk), .Q(ram[8543]) );
  DFF ram_reg_980__6_ ( .D(n12783), .CP(wclk), .Q(ram[8542]) );
  DFF ram_reg_980__5_ ( .D(n12782), .CP(wclk), .Q(ram[8541]) );
  DFF ram_reg_980__4_ ( .D(n12781), .CP(wclk), .Q(ram[8540]) );
  DFF ram_reg_980__3_ ( .D(n12780), .CP(wclk), .Q(ram[8539]) );
  DFF ram_reg_980__2_ ( .D(n12779), .CP(wclk), .Q(ram[8538]) );
  DFF ram_reg_980__1_ ( .D(n12778), .CP(wclk), .Q(ram[8537]) );
  DFF ram_reg_980__0_ ( .D(n12777), .CP(wclk), .Q(ram[8536]) );
  DFF ram_reg_996__7_ ( .D(n12656), .CP(wclk), .Q(ram[8415]) );
  DFF ram_reg_996__6_ ( .D(n12655), .CP(wclk), .Q(ram[8414]) );
  DFF ram_reg_996__5_ ( .D(n12654), .CP(wclk), .Q(ram[8413]) );
  DFF ram_reg_996__4_ ( .D(n12653), .CP(wclk), .Q(ram[8412]) );
  DFF ram_reg_996__3_ ( .D(n12652), .CP(wclk), .Q(ram[8411]) );
  DFF ram_reg_996__2_ ( .D(n12651), .CP(wclk), .Q(ram[8410]) );
  DFF ram_reg_996__1_ ( .D(n12650), .CP(wclk), .Q(ram[8409]) );
  DFF ram_reg_996__0_ ( .D(n12649), .CP(wclk), .Q(ram[8408]) );
  DFF ram_reg_1012__7_ ( .D(n12528), .CP(wclk), .Q(ram[8287]) );
  DFF ram_reg_1012__6_ ( .D(n12527), .CP(wclk), .Q(ram[8286]) );
  DFF ram_reg_1012__5_ ( .D(n12526), .CP(wclk), .Q(ram[8285]) );
  DFF ram_reg_1012__4_ ( .D(n12525), .CP(wclk), .Q(ram[8284]) );
  DFF ram_reg_1012__3_ ( .D(n12524), .CP(wclk), .Q(ram[8283]) );
  DFF ram_reg_1012__2_ ( .D(n12523), .CP(wclk), .Q(ram[8282]) );
  DFF ram_reg_1012__1_ ( .D(n12522), .CP(wclk), .Q(ram[8281]) );
  DFF ram_reg_1012__0_ ( .D(n12521), .CP(wclk), .Q(ram[8280]) );
  DFF ram_reg_1024__7_ ( .D(n12432), .CP(wclk), .Q(ram[8191]) );
  DFF ram_reg_1024__6_ ( .D(n12431), .CP(wclk), .Q(ram[8190]) );
  DFF ram_reg_1024__5_ ( .D(n12430), .CP(wclk), .Q(ram[8189]) );
  DFF ram_reg_1024__4_ ( .D(n12429), .CP(wclk), .Q(ram[8188]) );
  DFF ram_reg_1024__3_ ( .D(n12428), .CP(wclk), .Q(ram[8187]) );
  DFF ram_reg_1024__2_ ( .D(n12427), .CP(wclk), .Q(ram[8186]) );
  DFF ram_reg_1024__1_ ( .D(n12426), .CP(wclk), .Q(ram[8185]) );
  DFF ram_reg_1024__0_ ( .D(n12425), .CP(wclk), .Q(ram[8184]) );
  DFF ram_reg_1028__7_ ( .D(n12400), .CP(wclk), .Q(ram[8159]) );
  DFF ram_reg_1028__6_ ( .D(n12399), .CP(wclk), .Q(ram[8158]) );
  DFF ram_reg_1028__5_ ( .D(n12398), .CP(wclk), .Q(ram[8157]) );
  DFF ram_reg_1028__4_ ( .D(n12397), .CP(wclk), .Q(ram[8156]) );
  DFF ram_reg_1028__3_ ( .D(n12396), .CP(wclk), .Q(ram[8155]) );
  DFF ram_reg_1028__2_ ( .D(n12395), .CP(wclk), .Q(ram[8154]) );
  DFF ram_reg_1028__1_ ( .D(n12394), .CP(wclk), .Q(ram[8153]) );
  DFF ram_reg_1028__0_ ( .D(n12393), .CP(wclk), .Q(ram[8152]) );
  DFF ram_reg_1036__7_ ( .D(n12336), .CP(wclk), .Q(ram[8095]) );
  DFF ram_reg_1036__6_ ( .D(n12335), .CP(wclk), .Q(ram[8094]) );
  DFF ram_reg_1036__5_ ( .D(n12334), .CP(wclk), .Q(ram[8093]) );
  DFF ram_reg_1036__4_ ( .D(n12333), .CP(wclk), .Q(ram[8092]) );
  DFF ram_reg_1036__3_ ( .D(n12332), .CP(wclk), .Q(ram[8091]) );
  DFF ram_reg_1036__2_ ( .D(n12331), .CP(wclk), .Q(ram[8090]) );
  DFF ram_reg_1036__1_ ( .D(n12330), .CP(wclk), .Q(ram[8089]) );
  DFF ram_reg_1036__0_ ( .D(n12329), .CP(wclk), .Q(ram[8088]) );
  DFF ram_reg_1040__7_ ( .D(n12304), .CP(wclk), .Q(ram[8063]) );
  DFF ram_reg_1040__6_ ( .D(n12303), .CP(wclk), .Q(ram[8062]) );
  DFF ram_reg_1040__5_ ( .D(n12302), .CP(wclk), .Q(ram[8061]) );
  DFF ram_reg_1040__4_ ( .D(n12301), .CP(wclk), .Q(ram[8060]) );
  DFF ram_reg_1040__3_ ( .D(n12300), .CP(wclk), .Q(ram[8059]) );
  DFF ram_reg_1040__2_ ( .D(n12299), .CP(wclk), .Q(ram[8058]) );
  DFF ram_reg_1040__1_ ( .D(n12298), .CP(wclk), .Q(ram[8057]) );
  DFF ram_reg_1040__0_ ( .D(n12297), .CP(wclk), .Q(ram[8056]) );
  DFF ram_reg_1044__7_ ( .D(n12272), .CP(wclk), .Q(ram[8031]) );
  DFF ram_reg_1044__6_ ( .D(n12271), .CP(wclk), .Q(ram[8030]) );
  DFF ram_reg_1044__5_ ( .D(n12270), .CP(wclk), .Q(ram[8029]) );
  DFF ram_reg_1044__4_ ( .D(n12269), .CP(wclk), .Q(ram[8028]) );
  DFF ram_reg_1044__3_ ( .D(n12268), .CP(wclk), .Q(ram[8027]) );
  DFF ram_reg_1044__2_ ( .D(n12267), .CP(wclk), .Q(ram[8026]) );
  DFF ram_reg_1044__1_ ( .D(n12266), .CP(wclk), .Q(ram[8025]) );
  DFF ram_reg_1044__0_ ( .D(n12265), .CP(wclk), .Q(ram[8024]) );
  DFF ram_reg_1048__7_ ( .D(n12240), .CP(wclk), .Q(ram[7999]) );
  DFF ram_reg_1048__6_ ( .D(n12239), .CP(wclk), .Q(ram[7998]) );
  DFF ram_reg_1048__5_ ( .D(n12238), .CP(wclk), .Q(ram[7997]) );
  DFF ram_reg_1048__4_ ( .D(n12237), .CP(wclk), .Q(ram[7996]) );
  DFF ram_reg_1048__3_ ( .D(n12236), .CP(wclk), .Q(ram[7995]) );
  DFF ram_reg_1048__2_ ( .D(n12235), .CP(wclk), .Q(ram[7994]) );
  DFF ram_reg_1048__1_ ( .D(n12234), .CP(wclk), .Q(ram[7993]) );
  DFF ram_reg_1048__0_ ( .D(n12233), .CP(wclk), .Q(ram[7992]) );
  DFF ram_reg_1052__7_ ( .D(n12208), .CP(wclk), .Q(ram[7967]) );
  DFF ram_reg_1052__6_ ( .D(n12207), .CP(wclk), .Q(ram[7966]) );
  DFF ram_reg_1052__5_ ( .D(n12206), .CP(wclk), .Q(ram[7965]) );
  DFF ram_reg_1052__4_ ( .D(n12205), .CP(wclk), .Q(ram[7964]) );
  DFF ram_reg_1052__3_ ( .D(n12204), .CP(wclk), .Q(ram[7963]) );
  DFF ram_reg_1052__2_ ( .D(n12203), .CP(wclk), .Q(ram[7962]) );
  DFF ram_reg_1052__1_ ( .D(n12202), .CP(wclk), .Q(ram[7961]) );
  DFF ram_reg_1052__0_ ( .D(n12201), .CP(wclk), .Q(ram[7960]) );
  DFF ram_reg_1056__7_ ( .D(n12176), .CP(wclk), .Q(ram[7935]) );
  DFF ram_reg_1056__6_ ( .D(n12175), .CP(wclk), .Q(ram[7934]) );
  DFF ram_reg_1056__5_ ( .D(n12174), .CP(wclk), .Q(ram[7933]) );
  DFF ram_reg_1056__4_ ( .D(n12173), .CP(wclk), .Q(ram[7932]) );
  DFF ram_reg_1056__3_ ( .D(n12172), .CP(wclk), .Q(ram[7931]) );
  DFF ram_reg_1056__2_ ( .D(n12171), .CP(wclk), .Q(ram[7930]) );
  DFF ram_reg_1056__1_ ( .D(n12170), .CP(wclk), .Q(ram[7929]) );
  DFF ram_reg_1056__0_ ( .D(n12169), .CP(wclk), .Q(ram[7928]) );
  DFF ram_reg_1060__7_ ( .D(n12144), .CP(wclk), .Q(ram[7903]) );
  DFF ram_reg_1060__6_ ( .D(n12143), .CP(wclk), .Q(ram[7902]) );
  DFF ram_reg_1060__5_ ( .D(n12142), .CP(wclk), .Q(ram[7901]) );
  DFF ram_reg_1060__4_ ( .D(n12141), .CP(wclk), .Q(ram[7900]) );
  DFF ram_reg_1060__3_ ( .D(n12140), .CP(wclk), .Q(ram[7899]) );
  DFF ram_reg_1060__2_ ( .D(n12139), .CP(wclk), .Q(ram[7898]) );
  DFF ram_reg_1060__1_ ( .D(n12138), .CP(wclk), .Q(ram[7897]) );
  DFF ram_reg_1060__0_ ( .D(n12137), .CP(wclk), .Q(ram[7896]) );
  DFF ram_reg_1072__7_ ( .D(n12048), .CP(wclk), .Q(ram[7807]) );
  DFF ram_reg_1072__6_ ( .D(n12047), .CP(wclk), .Q(ram[7806]) );
  DFF ram_reg_1072__5_ ( .D(n12046), .CP(wclk), .Q(ram[7805]) );
  DFF ram_reg_1072__4_ ( .D(n12045), .CP(wclk), .Q(ram[7804]) );
  DFF ram_reg_1072__3_ ( .D(n12044), .CP(wclk), .Q(ram[7803]) );
  DFF ram_reg_1072__2_ ( .D(n12043), .CP(wclk), .Q(ram[7802]) );
  DFF ram_reg_1072__1_ ( .D(n12042), .CP(wclk), .Q(ram[7801]) );
  DFF ram_reg_1072__0_ ( .D(n12041), .CP(wclk), .Q(ram[7800]) );
  DFF ram_reg_1076__7_ ( .D(n12016), .CP(wclk), .Q(ram[7775]) );
  DFF ram_reg_1076__6_ ( .D(n12015), .CP(wclk), .Q(ram[7774]) );
  DFF ram_reg_1076__5_ ( .D(n12014), .CP(wclk), .Q(ram[7773]) );
  DFF ram_reg_1076__4_ ( .D(n12013), .CP(wclk), .Q(ram[7772]) );
  DFF ram_reg_1076__3_ ( .D(n12012), .CP(wclk), .Q(ram[7771]) );
  DFF ram_reg_1076__2_ ( .D(n12011), .CP(wclk), .Q(ram[7770]) );
  DFF ram_reg_1076__1_ ( .D(n12010), .CP(wclk), .Q(ram[7769]) );
  DFF ram_reg_1076__0_ ( .D(n12009), .CP(wclk), .Q(ram[7768]) );
  DFF ram_reg_1088__7_ ( .D(n11920), .CP(wclk), .Q(ram[7679]) );
  DFF ram_reg_1088__6_ ( .D(n11919), .CP(wclk), .Q(ram[7678]) );
  DFF ram_reg_1088__5_ ( .D(n11918), .CP(wclk), .Q(ram[7677]) );
  DFF ram_reg_1088__4_ ( .D(n11917), .CP(wclk), .Q(ram[7676]) );
  DFF ram_reg_1088__3_ ( .D(n11916), .CP(wclk), .Q(ram[7675]) );
  DFF ram_reg_1088__2_ ( .D(n11915), .CP(wclk), .Q(ram[7674]) );
  DFF ram_reg_1088__1_ ( .D(n11914), .CP(wclk), .Q(ram[7673]) );
  DFF ram_reg_1088__0_ ( .D(n11913), .CP(wclk), .Q(ram[7672]) );
  DFF ram_reg_1092__7_ ( .D(n11888), .CP(wclk), .Q(ram[7647]) );
  DFF ram_reg_1092__6_ ( .D(n11887), .CP(wclk), .Q(ram[7646]) );
  DFF ram_reg_1092__5_ ( .D(n11886), .CP(wclk), .Q(ram[7645]) );
  DFF ram_reg_1092__4_ ( .D(n11885), .CP(wclk), .Q(ram[7644]) );
  DFF ram_reg_1092__3_ ( .D(n11884), .CP(wclk), .Q(ram[7643]) );
  DFF ram_reg_1092__2_ ( .D(n11883), .CP(wclk), .Q(ram[7642]) );
  DFF ram_reg_1092__1_ ( .D(n11882), .CP(wclk), .Q(ram[7641]) );
  DFF ram_reg_1092__0_ ( .D(n11881), .CP(wclk), .Q(ram[7640]) );
  DFF ram_reg_1096__7_ ( .D(n11856), .CP(wclk), .Q(ram[7615]) );
  DFF ram_reg_1096__6_ ( .D(n11855), .CP(wclk), .Q(ram[7614]) );
  DFF ram_reg_1096__5_ ( .D(n11854), .CP(wclk), .Q(ram[7613]) );
  DFF ram_reg_1096__4_ ( .D(n11853), .CP(wclk), .Q(ram[7612]) );
  DFF ram_reg_1096__3_ ( .D(n11852), .CP(wclk), .Q(ram[7611]) );
  DFF ram_reg_1096__2_ ( .D(n11851), .CP(wclk), .Q(ram[7610]) );
  DFF ram_reg_1096__1_ ( .D(n11850), .CP(wclk), .Q(ram[7609]) );
  DFF ram_reg_1096__0_ ( .D(n11849), .CP(wclk), .Q(ram[7608]) );
  DFF ram_reg_1100__7_ ( .D(n11824), .CP(wclk), .Q(ram[7583]) );
  DFF ram_reg_1100__6_ ( .D(n11823), .CP(wclk), .Q(ram[7582]) );
  DFF ram_reg_1100__5_ ( .D(n11822), .CP(wclk), .Q(ram[7581]) );
  DFF ram_reg_1100__4_ ( .D(n11821), .CP(wclk), .Q(ram[7580]) );
  DFF ram_reg_1100__3_ ( .D(n11820), .CP(wclk), .Q(ram[7579]) );
  DFF ram_reg_1100__2_ ( .D(n11819), .CP(wclk), .Q(ram[7578]) );
  DFF ram_reg_1100__1_ ( .D(n11818), .CP(wclk), .Q(ram[7577]) );
  DFF ram_reg_1100__0_ ( .D(n11817), .CP(wclk), .Q(ram[7576]) );
  DFF ram_reg_1104__7_ ( .D(n11792), .CP(wclk), .Q(ram[7551]) );
  DFF ram_reg_1104__6_ ( .D(n11791), .CP(wclk), .Q(ram[7550]) );
  DFF ram_reg_1104__5_ ( .D(n11790), .CP(wclk), .Q(ram[7549]) );
  DFF ram_reg_1104__4_ ( .D(n11789), .CP(wclk), .Q(ram[7548]) );
  DFF ram_reg_1104__3_ ( .D(n11788), .CP(wclk), .Q(ram[7547]) );
  DFF ram_reg_1104__2_ ( .D(n11787), .CP(wclk), .Q(ram[7546]) );
  DFF ram_reg_1104__1_ ( .D(n11786), .CP(wclk), .Q(ram[7545]) );
  DFF ram_reg_1104__0_ ( .D(n11785), .CP(wclk), .Q(ram[7544]) );
  DFF ram_reg_1108__7_ ( .D(n11760), .CP(wclk), .Q(ram[7519]) );
  DFF ram_reg_1108__6_ ( .D(n11759), .CP(wclk), .Q(ram[7518]) );
  DFF ram_reg_1108__5_ ( .D(n11758), .CP(wclk), .Q(ram[7517]) );
  DFF ram_reg_1108__4_ ( .D(n11757), .CP(wclk), .Q(ram[7516]) );
  DFF ram_reg_1108__3_ ( .D(n11756), .CP(wclk), .Q(ram[7515]) );
  DFF ram_reg_1108__2_ ( .D(n11755), .CP(wclk), .Q(ram[7514]) );
  DFF ram_reg_1108__1_ ( .D(n11754), .CP(wclk), .Q(ram[7513]) );
  DFF ram_reg_1108__0_ ( .D(n11753), .CP(wclk), .Q(ram[7512]) );
  DFF ram_reg_1112__7_ ( .D(n11728), .CP(wclk), .Q(ram[7487]) );
  DFF ram_reg_1112__6_ ( .D(n11727), .CP(wclk), .Q(ram[7486]) );
  DFF ram_reg_1112__5_ ( .D(n11726), .CP(wclk), .Q(ram[7485]) );
  DFF ram_reg_1112__4_ ( .D(n11725), .CP(wclk), .Q(ram[7484]) );
  DFF ram_reg_1112__3_ ( .D(n11724), .CP(wclk), .Q(ram[7483]) );
  DFF ram_reg_1112__2_ ( .D(n11723), .CP(wclk), .Q(ram[7482]) );
  DFF ram_reg_1112__1_ ( .D(n11722), .CP(wclk), .Q(ram[7481]) );
  DFF ram_reg_1112__0_ ( .D(n11721), .CP(wclk), .Q(ram[7480]) );
  DFF ram_reg_1116__7_ ( .D(n11696), .CP(wclk), .Q(ram[7455]) );
  DFF ram_reg_1116__6_ ( .D(n11695), .CP(wclk), .Q(ram[7454]) );
  DFF ram_reg_1116__5_ ( .D(n11694), .CP(wclk), .Q(ram[7453]) );
  DFF ram_reg_1116__4_ ( .D(n11693), .CP(wclk), .Q(ram[7452]) );
  DFF ram_reg_1116__3_ ( .D(n11692), .CP(wclk), .Q(ram[7451]) );
  DFF ram_reg_1116__2_ ( .D(n11691), .CP(wclk), .Q(ram[7450]) );
  DFF ram_reg_1116__1_ ( .D(n11690), .CP(wclk), .Q(ram[7449]) );
  DFF ram_reg_1116__0_ ( .D(n11689), .CP(wclk), .Q(ram[7448]) );
  DFF ram_reg_1120__7_ ( .D(n11664), .CP(wclk), .Q(ram[7423]) );
  DFF ram_reg_1120__6_ ( .D(n11663), .CP(wclk), .Q(ram[7422]) );
  DFF ram_reg_1120__5_ ( .D(n11662), .CP(wclk), .Q(ram[7421]) );
  DFF ram_reg_1120__4_ ( .D(n11661), .CP(wclk), .Q(ram[7420]) );
  DFF ram_reg_1120__3_ ( .D(n11660), .CP(wclk), .Q(ram[7419]) );
  DFF ram_reg_1120__2_ ( .D(n11659), .CP(wclk), .Q(ram[7418]) );
  DFF ram_reg_1120__1_ ( .D(n11658), .CP(wclk), .Q(ram[7417]) );
  DFF ram_reg_1120__0_ ( .D(n11657), .CP(wclk), .Q(ram[7416]) );
  DFF ram_reg_1124__7_ ( .D(n11632), .CP(wclk), .Q(ram[7391]) );
  DFF ram_reg_1124__6_ ( .D(n11631), .CP(wclk), .Q(ram[7390]) );
  DFF ram_reg_1124__5_ ( .D(n11630), .CP(wclk), .Q(ram[7389]) );
  DFF ram_reg_1124__4_ ( .D(n11629), .CP(wclk), .Q(ram[7388]) );
  DFF ram_reg_1124__3_ ( .D(n11628), .CP(wclk), .Q(ram[7387]) );
  DFF ram_reg_1124__2_ ( .D(n11627), .CP(wclk), .Q(ram[7386]) );
  DFF ram_reg_1124__1_ ( .D(n11626), .CP(wclk), .Q(ram[7385]) );
  DFF ram_reg_1124__0_ ( .D(n11625), .CP(wclk), .Q(ram[7384]) );
  DFF ram_reg_1128__7_ ( .D(n11600), .CP(wclk), .Q(ram[7359]) );
  DFF ram_reg_1128__6_ ( .D(n11599), .CP(wclk), .Q(ram[7358]) );
  DFF ram_reg_1128__5_ ( .D(n11598), .CP(wclk), .Q(ram[7357]) );
  DFF ram_reg_1128__4_ ( .D(n11597), .CP(wclk), .Q(ram[7356]) );
  DFF ram_reg_1128__3_ ( .D(n11596), .CP(wclk), .Q(ram[7355]) );
  DFF ram_reg_1128__2_ ( .D(n11595), .CP(wclk), .Q(ram[7354]) );
  DFF ram_reg_1128__1_ ( .D(n11594), .CP(wclk), .Q(ram[7353]) );
  DFF ram_reg_1128__0_ ( .D(n11593), .CP(wclk), .Q(ram[7352]) );
  DFF ram_reg_1132__7_ ( .D(n11568), .CP(wclk), .Q(ram[7327]) );
  DFF ram_reg_1132__6_ ( .D(n11567), .CP(wclk), .Q(ram[7326]) );
  DFF ram_reg_1132__5_ ( .D(n11566), .CP(wclk), .Q(ram[7325]) );
  DFF ram_reg_1132__4_ ( .D(n11565), .CP(wclk), .Q(ram[7324]) );
  DFF ram_reg_1132__3_ ( .D(n11564), .CP(wclk), .Q(ram[7323]) );
  DFF ram_reg_1132__2_ ( .D(n11563), .CP(wclk), .Q(ram[7322]) );
  DFF ram_reg_1132__1_ ( .D(n11562), .CP(wclk), .Q(ram[7321]) );
  DFF ram_reg_1132__0_ ( .D(n11561), .CP(wclk), .Q(ram[7320]) );
  DFF ram_reg_1136__7_ ( .D(n11536), .CP(wclk), .Q(ram[7295]) );
  DFF ram_reg_1136__6_ ( .D(n11535), .CP(wclk), .Q(ram[7294]) );
  DFF ram_reg_1136__5_ ( .D(n11534), .CP(wclk), .Q(ram[7293]) );
  DFF ram_reg_1136__4_ ( .D(n11533), .CP(wclk), .Q(ram[7292]) );
  DFF ram_reg_1136__3_ ( .D(n11532), .CP(wclk), .Q(ram[7291]) );
  DFF ram_reg_1136__2_ ( .D(n11531), .CP(wclk), .Q(ram[7290]) );
  DFF ram_reg_1136__1_ ( .D(n11530), .CP(wclk), .Q(ram[7289]) );
  DFF ram_reg_1136__0_ ( .D(n11529), .CP(wclk), .Q(ram[7288]) );
  DFF ram_reg_1140__7_ ( .D(n11504), .CP(wclk), .Q(ram[7263]) );
  DFF ram_reg_1140__6_ ( .D(n11503), .CP(wclk), .Q(ram[7262]) );
  DFF ram_reg_1140__5_ ( .D(n11502), .CP(wclk), .Q(ram[7261]) );
  DFF ram_reg_1140__4_ ( .D(n11501), .CP(wclk), .Q(ram[7260]) );
  DFF ram_reg_1140__3_ ( .D(n11500), .CP(wclk), .Q(ram[7259]) );
  DFF ram_reg_1140__2_ ( .D(n11499), .CP(wclk), .Q(ram[7258]) );
  DFF ram_reg_1140__1_ ( .D(n11498), .CP(wclk), .Q(ram[7257]) );
  DFF ram_reg_1140__0_ ( .D(n11497), .CP(wclk), .Q(ram[7256]) );
  DFF ram_reg_1144__7_ ( .D(n11472), .CP(wclk), .Q(ram[7231]) );
  DFF ram_reg_1144__6_ ( .D(n11471), .CP(wclk), .Q(ram[7230]) );
  DFF ram_reg_1144__5_ ( .D(n11470), .CP(wclk), .Q(ram[7229]) );
  DFF ram_reg_1144__4_ ( .D(n11469), .CP(wclk), .Q(ram[7228]) );
  DFF ram_reg_1144__3_ ( .D(n11468), .CP(wclk), .Q(ram[7227]) );
  DFF ram_reg_1144__2_ ( .D(n11467), .CP(wclk), .Q(ram[7226]) );
  DFF ram_reg_1144__1_ ( .D(n11466), .CP(wclk), .Q(ram[7225]) );
  DFF ram_reg_1144__0_ ( .D(n11465), .CP(wclk), .Q(ram[7224]) );
  DFF ram_reg_1148__7_ ( .D(n11440), .CP(wclk), .Q(ram[7199]) );
  DFF ram_reg_1148__6_ ( .D(n11439), .CP(wclk), .Q(ram[7198]) );
  DFF ram_reg_1148__5_ ( .D(n11438), .CP(wclk), .Q(ram[7197]) );
  DFF ram_reg_1148__4_ ( .D(n11437), .CP(wclk), .Q(ram[7196]) );
  DFF ram_reg_1148__3_ ( .D(n11436), .CP(wclk), .Q(ram[7195]) );
  DFF ram_reg_1148__2_ ( .D(n11435), .CP(wclk), .Q(ram[7194]) );
  DFF ram_reg_1148__1_ ( .D(n11434), .CP(wclk), .Q(ram[7193]) );
  DFF ram_reg_1148__0_ ( .D(n11433), .CP(wclk), .Q(ram[7192]) );
  DFF ram_reg_1156__7_ ( .D(n11376), .CP(wclk), .Q(ram[7135]) );
  DFF ram_reg_1156__6_ ( .D(n11375), .CP(wclk), .Q(ram[7134]) );
  DFF ram_reg_1156__5_ ( .D(n11374), .CP(wclk), .Q(ram[7133]) );
  DFF ram_reg_1156__4_ ( .D(n11373), .CP(wclk), .Q(ram[7132]) );
  DFF ram_reg_1156__3_ ( .D(n11372), .CP(wclk), .Q(ram[7131]) );
  DFF ram_reg_1156__2_ ( .D(n11371), .CP(wclk), .Q(ram[7130]) );
  DFF ram_reg_1156__1_ ( .D(n11370), .CP(wclk), .Q(ram[7129]) );
  DFF ram_reg_1156__0_ ( .D(n11369), .CP(wclk), .Q(ram[7128]) );
  DFF ram_reg_1168__7_ ( .D(n11280), .CP(wclk), .Q(ram[7039]) );
  DFF ram_reg_1168__6_ ( .D(n11279), .CP(wclk), .Q(ram[7038]) );
  DFF ram_reg_1168__5_ ( .D(n11278), .CP(wclk), .Q(ram[7037]) );
  DFF ram_reg_1168__4_ ( .D(n11277), .CP(wclk), .Q(ram[7036]) );
  DFF ram_reg_1168__3_ ( .D(n11276), .CP(wclk), .Q(ram[7035]) );
  DFF ram_reg_1168__2_ ( .D(n11275), .CP(wclk), .Q(ram[7034]) );
  DFF ram_reg_1168__1_ ( .D(n11274), .CP(wclk), .Q(ram[7033]) );
  DFF ram_reg_1168__0_ ( .D(n11273), .CP(wclk), .Q(ram[7032]) );
  DFF ram_reg_1172__7_ ( .D(n11248), .CP(wclk), .Q(ram[7007]) );
  DFF ram_reg_1172__6_ ( .D(n11247), .CP(wclk), .Q(ram[7006]) );
  DFF ram_reg_1172__5_ ( .D(n11246), .CP(wclk), .Q(ram[7005]) );
  DFF ram_reg_1172__4_ ( .D(n11245), .CP(wclk), .Q(ram[7004]) );
  DFF ram_reg_1172__3_ ( .D(n11244), .CP(wclk), .Q(ram[7003]) );
  DFF ram_reg_1172__2_ ( .D(n11243), .CP(wclk), .Q(ram[7002]) );
  DFF ram_reg_1172__1_ ( .D(n11242), .CP(wclk), .Q(ram[7001]) );
  DFF ram_reg_1172__0_ ( .D(n11241), .CP(wclk), .Q(ram[7000]) );
  DFF ram_reg_1188__7_ ( .D(n11120), .CP(wclk), .Q(ram[6879]) );
  DFF ram_reg_1188__6_ ( .D(n11119), .CP(wclk), .Q(ram[6878]) );
  DFF ram_reg_1188__5_ ( .D(n11118), .CP(wclk), .Q(ram[6877]) );
  DFF ram_reg_1188__4_ ( .D(n11117), .CP(wclk), .Q(ram[6876]) );
  DFF ram_reg_1188__3_ ( .D(n11116), .CP(wclk), .Q(ram[6875]) );
  DFF ram_reg_1188__2_ ( .D(n11115), .CP(wclk), .Q(ram[6874]) );
  DFF ram_reg_1188__1_ ( .D(n11114), .CP(wclk), .Q(ram[6873]) );
  DFF ram_reg_1188__0_ ( .D(n11113), .CP(wclk), .Q(ram[6872]) );
  DFF ram_reg_1204__7_ ( .D(n10992), .CP(wclk), .Q(ram[6751]) );
  DFF ram_reg_1204__6_ ( .D(n10991), .CP(wclk), .Q(ram[6750]) );
  DFF ram_reg_1204__5_ ( .D(n10990), .CP(wclk), .Q(ram[6749]) );
  DFF ram_reg_1204__4_ ( .D(n10989), .CP(wclk), .Q(ram[6748]) );
  DFF ram_reg_1204__3_ ( .D(n10988), .CP(wclk), .Q(ram[6747]) );
  DFF ram_reg_1204__2_ ( .D(n10987), .CP(wclk), .Q(ram[6746]) );
  DFF ram_reg_1204__1_ ( .D(n10986), .CP(wclk), .Q(ram[6745]) );
  DFF ram_reg_1204__0_ ( .D(n10985), .CP(wclk), .Q(ram[6744]) );
  DFF ram_reg_1216__7_ ( .D(n10896), .CP(wclk), .Q(ram[6655]) );
  DFF ram_reg_1216__6_ ( .D(n10895), .CP(wclk), .Q(ram[6654]) );
  DFF ram_reg_1216__5_ ( .D(n10894), .CP(wclk), .Q(ram[6653]) );
  DFF ram_reg_1216__4_ ( .D(n10893), .CP(wclk), .Q(ram[6652]) );
  DFF ram_reg_1216__3_ ( .D(n10892), .CP(wclk), .Q(ram[6651]) );
  DFF ram_reg_1216__2_ ( .D(n10891), .CP(wclk), .Q(ram[6650]) );
  DFF ram_reg_1216__1_ ( .D(n10890), .CP(wclk), .Q(ram[6649]) );
  DFF ram_reg_1216__0_ ( .D(n10889), .CP(wclk), .Q(ram[6648]) );
  DFF ram_reg_1220__7_ ( .D(n10864), .CP(wclk), .Q(ram[6623]) );
  DFF ram_reg_1220__6_ ( .D(n10863), .CP(wclk), .Q(ram[6622]) );
  DFF ram_reg_1220__5_ ( .D(n10862), .CP(wclk), .Q(ram[6621]) );
  DFF ram_reg_1220__4_ ( .D(n10861), .CP(wclk), .Q(ram[6620]) );
  DFF ram_reg_1220__3_ ( .D(n10860), .CP(wclk), .Q(ram[6619]) );
  DFF ram_reg_1220__2_ ( .D(n10859), .CP(wclk), .Q(ram[6618]) );
  DFF ram_reg_1220__1_ ( .D(n10858), .CP(wclk), .Q(ram[6617]) );
  DFF ram_reg_1220__0_ ( .D(n10857), .CP(wclk), .Q(ram[6616]) );
  DFF ram_reg_1232__7_ ( .D(n10768), .CP(wclk), .Q(ram[6527]) );
  DFF ram_reg_1232__6_ ( .D(n10767), .CP(wclk), .Q(ram[6526]) );
  DFF ram_reg_1232__5_ ( .D(n10766), .CP(wclk), .Q(ram[6525]) );
  DFF ram_reg_1232__4_ ( .D(n10765), .CP(wclk), .Q(ram[6524]) );
  DFF ram_reg_1232__3_ ( .D(n10764), .CP(wclk), .Q(ram[6523]) );
  DFF ram_reg_1232__2_ ( .D(n10763), .CP(wclk), .Q(ram[6522]) );
  DFF ram_reg_1232__1_ ( .D(n10762), .CP(wclk), .Q(ram[6521]) );
  DFF ram_reg_1232__0_ ( .D(n10761), .CP(wclk), .Q(ram[6520]) );
  DFF ram_reg_1236__7_ ( .D(n10736), .CP(wclk), .Q(ram[6495]) );
  DFF ram_reg_1236__6_ ( .D(n10735), .CP(wclk), .Q(ram[6494]) );
  DFF ram_reg_1236__5_ ( .D(n10734), .CP(wclk), .Q(ram[6493]) );
  DFF ram_reg_1236__4_ ( .D(n10733), .CP(wclk), .Q(ram[6492]) );
  DFF ram_reg_1236__3_ ( .D(n10732), .CP(wclk), .Q(ram[6491]) );
  DFF ram_reg_1236__2_ ( .D(n10731), .CP(wclk), .Q(ram[6490]) );
  DFF ram_reg_1236__1_ ( .D(n10730), .CP(wclk), .Q(ram[6489]) );
  DFF ram_reg_1236__0_ ( .D(n10729), .CP(wclk), .Q(ram[6488]) );
  DFF ram_reg_1244__7_ ( .D(n10672), .CP(wclk), .Q(ram[6431]) );
  DFF ram_reg_1244__6_ ( .D(n10671), .CP(wclk), .Q(ram[6430]) );
  DFF ram_reg_1244__5_ ( .D(n10670), .CP(wclk), .Q(ram[6429]) );
  DFF ram_reg_1244__4_ ( .D(n10669), .CP(wclk), .Q(ram[6428]) );
  DFF ram_reg_1244__3_ ( .D(n10668), .CP(wclk), .Q(ram[6427]) );
  DFF ram_reg_1244__2_ ( .D(n10667), .CP(wclk), .Q(ram[6426]) );
  DFF ram_reg_1244__1_ ( .D(n10666), .CP(wclk), .Q(ram[6425]) );
  DFF ram_reg_1244__0_ ( .D(n10665), .CP(wclk), .Q(ram[6424]) );
  DFF ram_reg_1252__7_ ( .D(n10608), .CP(wclk), .Q(ram[6367]) );
  DFF ram_reg_1252__6_ ( .D(n10607), .CP(wclk), .Q(ram[6366]) );
  DFF ram_reg_1252__5_ ( .D(n10606), .CP(wclk), .Q(ram[6365]) );
  DFF ram_reg_1252__4_ ( .D(n10605), .CP(wclk), .Q(ram[6364]) );
  DFF ram_reg_1252__3_ ( .D(n10604), .CP(wclk), .Q(ram[6363]) );
  DFF ram_reg_1252__2_ ( .D(n10603), .CP(wclk), .Q(ram[6362]) );
  DFF ram_reg_1252__1_ ( .D(n10602), .CP(wclk), .Q(ram[6361]) );
  DFF ram_reg_1252__0_ ( .D(n10601), .CP(wclk), .Q(ram[6360]) );
  DFF ram_reg_1268__7_ ( .D(n10480), .CP(wclk), .Q(ram[6239]) );
  DFF ram_reg_1268__6_ ( .D(n10479), .CP(wclk), .Q(ram[6238]) );
  DFF ram_reg_1268__5_ ( .D(n10478), .CP(wclk), .Q(ram[6237]) );
  DFF ram_reg_1268__4_ ( .D(n10477), .CP(wclk), .Q(ram[6236]) );
  DFF ram_reg_1268__3_ ( .D(n10476), .CP(wclk), .Q(ram[6235]) );
  DFF ram_reg_1268__2_ ( .D(n10475), .CP(wclk), .Q(ram[6234]) );
  DFF ram_reg_1268__1_ ( .D(n10474), .CP(wclk), .Q(ram[6233]) );
  DFF ram_reg_1268__0_ ( .D(n10473), .CP(wclk), .Q(ram[6232]) );
  DFF ram_reg_1280__7_ ( .D(n10384), .CP(wclk), .Q(ram[6143]) );
  DFF ram_reg_1280__6_ ( .D(n10383), .CP(wclk), .Q(ram[6142]) );
  DFF ram_reg_1280__5_ ( .D(n10382), .CP(wclk), .Q(ram[6141]) );
  DFF ram_reg_1280__4_ ( .D(n10381), .CP(wclk), .Q(ram[6140]) );
  DFF ram_reg_1280__3_ ( .D(n10380), .CP(wclk), .Q(ram[6139]) );
  DFF ram_reg_1280__2_ ( .D(n10379), .CP(wclk), .Q(ram[6138]) );
  DFF ram_reg_1280__1_ ( .D(n10378), .CP(wclk), .Q(ram[6137]) );
  DFF ram_reg_1280__0_ ( .D(n10377), .CP(wclk), .Q(ram[6136]) );
  DFF ram_reg_1284__7_ ( .D(n10352), .CP(wclk), .Q(ram[6111]) );
  DFF ram_reg_1284__6_ ( .D(n10351), .CP(wclk), .Q(ram[6110]) );
  DFF ram_reg_1284__5_ ( .D(n10350), .CP(wclk), .Q(ram[6109]) );
  DFF ram_reg_1284__4_ ( .D(n10349), .CP(wclk), .Q(ram[6108]) );
  DFF ram_reg_1284__3_ ( .D(n10348), .CP(wclk), .Q(ram[6107]) );
  DFF ram_reg_1284__2_ ( .D(n10347), .CP(wclk), .Q(ram[6106]) );
  DFF ram_reg_1284__1_ ( .D(n10346), .CP(wclk), .Q(ram[6105]) );
  DFF ram_reg_1284__0_ ( .D(n10345), .CP(wclk), .Q(ram[6104]) );
  DFF ram_reg_1296__7_ ( .D(n10256), .CP(wclk), .Q(ram[6015]) );
  DFF ram_reg_1296__6_ ( .D(n10255), .CP(wclk), .Q(ram[6014]) );
  DFF ram_reg_1296__5_ ( .D(n10254), .CP(wclk), .Q(ram[6013]) );
  DFF ram_reg_1296__4_ ( .D(n10253), .CP(wclk), .Q(ram[6012]) );
  DFF ram_reg_1296__3_ ( .D(n10252), .CP(wclk), .Q(ram[6011]) );
  DFF ram_reg_1296__2_ ( .D(n10251), .CP(wclk), .Q(ram[6010]) );
  DFF ram_reg_1296__1_ ( .D(n10250), .CP(wclk), .Q(ram[6009]) );
  DFF ram_reg_1296__0_ ( .D(n10249), .CP(wclk), .Q(ram[6008]) );
  DFF ram_reg_1300__7_ ( .D(n10224), .CP(wclk), .Q(ram[5983]) );
  DFF ram_reg_1300__6_ ( .D(n10223), .CP(wclk), .Q(ram[5982]) );
  DFF ram_reg_1300__5_ ( .D(n10222), .CP(wclk), .Q(ram[5981]) );
  DFF ram_reg_1300__4_ ( .D(n10221), .CP(wclk), .Q(ram[5980]) );
  DFF ram_reg_1300__3_ ( .D(n10220), .CP(wclk), .Q(ram[5979]) );
  DFF ram_reg_1300__2_ ( .D(n10219), .CP(wclk), .Q(ram[5978]) );
  DFF ram_reg_1300__1_ ( .D(n10218), .CP(wclk), .Q(ram[5977]) );
  DFF ram_reg_1300__0_ ( .D(n10217), .CP(wclk), .Q(ram[5976]) );
  DFF ram_reg_1316__7_ ( .D(n10096), .CP(wclk), .Q(ram[5855]) );
  DFF ram_reg_1316__6_ ( .D(n10095), .CP(wclk), .Q(ram[5854]) );
  DFF ram_reg_1316__5_ ( .D(n10094), .CP(wclk), .Q(ram[5853]) );
  DFF ram_reg_1316__4_ ( .D(n10093), .CP(wclk), .Q(ram[5852]) );
  DFF ram_reg_1316__3_ ( .D(n10092), .CP(wclk), .Q(ram[5851]) );
  DFF ram_reg_1316__2_ ( .D(n10091), .CP(wclk), .Q(ram[5850]) );
  DFF ram_reg_1316__1_ ( .D(n10090), .CP(wclk), .Q(ram[5849]) );
  DFF ram_reg_1316__0_ ( .D(n10089), .CP(wclk), .Q(ram[5848]) );
  DFF ram_reg_1332__7_ ( .D(n9968), .CP(wclk), .Q(ram[5727]) );
  DFF ram_reg_1332__6_ ( .D(n9967), .CP(wclk), .Q(ram[5726]) );
  DFF ram_reg_1332__5_ ( .D(n9966), .CP(wclk), .Q(ram[5725]) );
  DFF ram_reg_1332__4_ ( .D(n9965), .CP(wclk), .Q(ram[5724]) );
  DFF ram_reg_1332__3_ ( .D(n9964), .CP(wclk), .Q(ram[5723]) );
  DFF ram_reg_1332__2_ ( .D(n9963), .CP(wclk), .Q(ram[5722]) );
  DFF ram_reg_1332__1_ ( .D(n9962), .CP(wclk), .Q(ram[5721]) );
  DFF ram_reg_1332__0_ ( .D(n9961), .CP(wclk), .Q(ram[5720]) );
  DFF ram_reg_1344__7_ ( .D(n9872), .CP(wclk), .Q(ram[5631]) );
  DFF ram_reg_1344__6_ ( .D(n9871), .CP(wclk), .Q(ram[5630]) );
  DFF ram_reg_1344__5_ ( .D(n9870), .CP(wclk), .Q(ram[5629]) );
  DFF ram_reg_1344__4_ ( .D(n9869), .CP(wclk), .Q(ram[5628]) );
  DFF ram_reg_1344__3_ ( .D(n9868), .CP(wclk), .Q(ram[5627]) );
  DFF ram_reg_1344__2_ ( .D(n9867), .CP(wclk), .Q(ram[5626]) );
  DFF ram_reg_1344__1_ ( .D(n9866), .CP(wclk), .Q(ram[5625]) );
  DFF ram_reg_1344__0_ ( .D(n9865), .CP(wclk), .Q(ram[5624]) );
  DFF ram_reg_1348__7_ ( .D(n9840), .CP(wclk), .Q(ram[5599]) );
  DFF ram_reg_1348__6_ ( .D(n9839), .CP(wclk), .Q(ram[5598]) );
  DFF ram_reg_1348__5_ ( .D(n9838), .CP(wclk), .Q(ram[5597]) );
  DFF ram_reg_1348__4_ ( .D(n9837), .CP(wclk), .Q(ram[5596]) );
  DFF ram_reg_1348__3_ ( .D(n9836), .CP(wclk), .Q(ram[5595]) );
  DFF ram_reg_1348__2_ ( .D(n9835), .CP(wclk), .Q(ram[5594]) );
  DFF ram_reg_1348__1_ ( .D(n9834), .CP(wclk), .Q(ram[5593]) );
  DFF ram_reg_1348__0_ ( .D(n9833), .CP(wclk), .Q(ram[5592]) );
  DFF ram_reg_1356__7_ ( .D(n9776), .CP(wclk), .Q(ram[5535]) );
  DFF ram_reg_1356__6_ ( .D(n9775), .CP(wclk), .Q(ram[5534]) );
  DFF ram_reg_1356__5_ ( .D(n9774), .CP(wclk), .Q(ram[5533]) );
  DFF ram_reg_1356__4_ ( .D(n9773), .CP(wclk), .Q(ram[5532]) );
  DFF ram_reg_1356__3_ ( .D(n9772), .CP(wclk), .Q(ram[5531]) );
  DFF ram_reg_1356__2_ ( .D(n9771), .CP(wclk), .Q(ram[5530]) );
  DFF ram_reg_1356__1_ ( .D(n9770), .CP(wclk), .Q(ram[5529]) );
  DFF ram_reg_1356__0_ ( .D(n9769), .CP(wclk), .Q(ram[5528]) );
  DFF ram_reg_1360__7_ ( .D(n9744), .CP(wclk), .Q(ram[5503]) );
  DFF ram_reg_1360__6_ ( .D(n9743), .CP(wclk), .Q(ram[5502]) );
  DFF ram_reg_1360__5_ ( .D(n9742), .CP(wclk), .Q(ram[5501]) );
  DFF ram_reg_1360__4_ ( .D(n9741), .CP(wclk), .Q(ram[5500]) );
  DFF ram_reg_1360__3_ ( .D(n9740), .CP(wclk), .Q(ram[5499]) );
  DFF ram_reg_1360__2_ ( .D(n9739), .CP(wclk), .Q(ram[5498]) );
  DFF ram_reg_1360__1_ ( .D(n9738), .CP(wclk), .Q(ram[5497]) );
  DFF ram_reg_1360__0_ ( .D(n9737), .CP(wclk), .Q(ram[5496]) );
  DFF ram_reg_1364__7_ ( .D(n9712), .CP(wclk), .Q(ram[5471]) );
  DFF ram_reg_1364__6_ ( .D(n9711), .CP(wclk), .Q(ram[5470]) );
  DFF ram_reg_1364__5_ ( .D(n9710), .CP(wclk), .Q(ram[5469]) );
  DFF ram_reg_1364__4_ ( .D(n9709), .CP(wclk), .Q(ram[5468]) );
  DFF ram_reg_1364__3_ ( .D(n9708), .CP(wclk), .Q(ram[5467]) );
  DFF ram_reg_1364__2_ ( .D(n9707), .CP(wclk), .Q(ram[5466]) );
  DFF ram_reg_1364__1_ ( .D(n9706), .CP(wclk), .Q(ram[5465]) );
  DFF ram_reg_1364__0_ ( .D(n9705), .CP(wclk), .Q(ram[5464]) );
  DFF ram_reg_1368__7_ ( .D(n9680), .CP(wclk), .Q(ram[5439]) );
  DFF ram_reg_1368__6_ ( .D(n9679), .CP(wclk), .Q(ram[5438]) );
  DFF ram_reg_1368__5_ ( .D(n9678), .CP(wclk), .Q(ram[5437]) );
  DFF ram_reg_1368__4_ ( .D(n9677), .CP(wclk), .Q(ram[5436]) );
  DFF ram_reg_1368__3_ ( .D(n9676), .CP(wclk), .Q(ram[5435]) );
  DFF ram_reg_1368__2_ ( .D(n9675), .CP(wclk), .Q(ram[5434]) );
  DFF ram_reg_1368__1_ ( .D(n9674), .CP(wclk), .Q(ram[5433]) );
  DFF ram_reg_1368__0_ ( .D(n9673), .CP(wclk), .Q(ram[5432]) );
  DFF ram_reg_1372__7_ ( .D(n9648), .CP(wclk), .Q(ram[5407]) );
  DFF ram_reg_1372__6_ ( .D(n9647), .CP(wclk), .Q(ram[5406]) );
  DFF ram_reg_1372__5_ ( .D(n9646), .CP(wclk), .Q(ram[5405]) );
  DFF ram_reg_1372__4_ ( .D(n9645), .CP(wclk), .Q(ram[5404]) );
  DFF ram_reg_1372__3_ ( .D(n9644), .CP(wclk), .Q(ram[5403]) );
  DFF ram_reg_1372__2_ ( .D(n9643), .CP(wclk), .Q(ram[5402]) );
  DFF ram_reg_1372__1_ ( .D(n9642), .CP(wclk), .Q(ram[5401]) );
  DFF ram_reg_1372__0_ ( .D(n9641), .CP(wclk), .Q(ram[5400]) );
  DFF ram_reg_1376__7_ ( .D(n9616), .CP(wclk), .Q(ram[5375]) );
  DFF ram_reg_1376__6_ ( .D(n9615), .CP(wclk), .Q(ram[5374]) );
  DFF ram_reg_1376__5_ ( .D(n9614), .CP(wclk), .Q(ram[5373]) );
  DFF ram_reg_1376__4_ ( .D(n9613), .CP(wclk), .Q(ram[5372]) );
  DFF ram_reg_1376__3_ ( .D(n9612), .CP(wclk), .Q(ram[5371]) );
  DFF ram_reg_1376__2_ ( .D(n9611), .CP(wclk), .Q(ram[5370]) );
  DFF ram_reg_1376__1_ ( .D(n9610), .CP(wclk), .Q(ram[5369]) );
  DFF ram_reg_1376__0_ ( .D(n9609), .CP(wclk), .Q(ram[5368]) );
  DFF ram_reg_1380__7_ ( .D(n9584), .CP(wclk), .Q(ram[5343]) );
  DFF ram_reg_1380__6_ ( .D(n9583), .CP(wclk), .Q(ram[5342]) );
  DFF ram_reg_1380__5_ ( .D(n9582), .CP(wclk), .Q(ram[5341]) );
  DFF ram_reg_1380__4_ ( .D(n9581), .CP(wclk), .Q(ram[5340]) );
  DFF ram_reg_1380__3_ ( .D(n9580), .CP(wclk), .Q(ram[5339]) );
  DFF ram_reg_1380__2_ ( .D(n9579), .CP(wclk), .Q(ram[5338]) );
  DFF ram_reg_1380__1_ ( .D(n9578), .CP(wclk), .Q(ram[5337]) );
  DFF ram_reg_1380__0_ ( .D(n9577), .CP(wclk), .Q(ram[5336]) );
  DFF ram_reg_1392__7_ ( .D(n9488), .CP(wclk), .Q(ram[5247]) );
  DFF ram_reg_1392__6_ ( .D(n9487), .CP(wclk), .Q(ram[5246]) );
  DFF ram_reg_1392__5_ ( .D(n9486), .CP(wclk), .Q(ram[5245]) );
  DFF ram_reg_1392__4_ ( .D(n9485), .CP(wclk), .Q(ram[5244]) );
  DFF ram_reg_1392__3_ ( .D(n9484), .CP(wclk), .Q(ram[5243]) );
  DFF ram_reg_1392__2_ ( .D(n9483), .CP(wclk), .Q(ram[5242]) );
  DFF ram_reg_1392__1_ ( .D(n9482), .CP(wclk), .Q(ram[5241]) );
  DFF ram_reg_1392__0_ ( .D(n9481), .CP(wclk), .Q(ram[5240]) );
  DFF ram_reg_1396__7_ ( .D(n9456), .CP(wclk), .Q(ram[5215]) );
  DFF ram_reg_1396__6_ ( .D(n9455), .CP(wclk), .Q(ram[5214]) );
  DFF ram_reg_1396__5_ ( .D(n9454), .CP(wclk), .Q(ram[5213]) );
  DFF ram_reg_1396__4_ ( .D(n9453), .CP(wclk), .Q(ram[5212]) );
  DFF ram_reg_1396__3_ ( .D(n9452), .CP(wclk), .Q(ram[5211]) );
  DFF ram_reg_1396__2_ ( .D(n9451), .CP(wclk), .Q(ram[5210]) );
  DFF ram_reg_1396__1_ ( .D(n9450), .CP(wclk), .Q(ram[5209]) );
  DFF ram_reg_1396__0_ ( .D(n9449), .CP(wclk), .Q(ram[5208]) );
  DFF ram_reg_1428__7_ ( .D(n9200), .CP(wclk), .Q(ram[4959]) );
  DFF ram_reg_1428__6_ ( .D(n9199), .CP(wclk), .Q(ram[4958]) );
  DFF ram_reg_1428__5_ ( .D(n9198), .CP(wclk), .Q(ram[4957]) );
  DFF ram_reg_1428__4_ ( .D(n9197), .CP(wclk), .Q(ram[4956]) );
  DFF ram_reg_1428__3_ ( .D(n9196), .CP(wclk), .Q(ram[4955]) );
  DFF ram_reg_1428__2_ ( .D(n9195), .CP(wclk), .Q(ram[4954]) );
  DFF ram_reg_1428__1_ ( .D(n9194), .CP(wclk), .Q(ram[4953]) );
  DFF ram_reg_1428__0_ ( .D(n9193), .CP(wclk), .Q(ram[4952]) );
  DFF ram_reg_1476__7_ ( .D(n8816), .CP(wclk), .Q(ram[4575]) );
  DFF ram_reg_1476__6_ ( .D(n8815), .CP(wclk), .Q(ram[4574]) );
  DFF ram_reg_1476__5_ ( .D(n8814), .CP(wclk), .Q(ram[4573]) );
  DFF ram_reg_1476__4_ ( .D(n8813), .CP(wclk), .Q(ram[4572]) );
  DFF ram_reg_1476__3_ ( .D(n8812), .CP(wclk), .Q(ram[4571]) );
  DFF ram_reg_1476__2_ ( .D(n8811), .CP(wclk), .Q(ram[4570]) );
  DFF ram_reg_1476__1_ ( .D(n8810), .CP(wclk), .Q(ram[4569]) );
  DFF ram_reg_1476__0_ ( .D(n8809), .CP(wclk), .Q(ram[4568]) );
  DFF ram_reg_1492__7_ ( .D(n8688), .CP(wclk), .Q(ram[4447]) );
  DFF ram_reg_1492__6_ ( .D(n8687), .CP(wclk), .Q(ram[4446]) );
  DFF ram_reg_1492__5_ ( .D(n8686), .CP(wclk), .Q(ram[4445]) );
  DFF ram_reg_1492__4_ ( .D(n8685), .CP(wclk), .Q(ram[4444]) );
  DFF ram_reg_1492__3_ ( .D(n8684), .CP(wclk), .Q(ram[4443]) );
  DFF ram_reg_1492__2_ ( .D(n8683), .CP(wclk), .Q(ram[4442]) );
  DFF ram_reg_1492__1_ ( .D(n8682), .CP(wclk), .Q(ram[4441]) );
  DFF ram_reg_1492__0_ ( .D(n8681), .CP(wclk), .Q(ram[4440]) );
  DFF ram_reg_1536__7_ ( .D(n8336), .CP(wclk), .Q(ram[4095]) );
  DFF ram_reg_1536__6_ ( .D(n8335), .CP(wclk), .Q(ram[4094]) );
  DFF ram_reg_1536__5_ ( .D(n8334), .CP(wclk), .Q(ram[4093]) );
  DFF ram_reg_1536__4_ ( .D(n8333), .CP(wclk), .Q(ram[4092]) );
  DFF ram_reg_1536__3_ ( .D(n8332), .CP(wclk), .Q(ram[4091]) );
  DFF ram_reg_1536__2_ ( .D(n8331), .CP(wclk), .Q(ram[4090]) );
  DFF ram_reg_1536__1_ ( .D(n8330), .CP(wclk), .Q(ram[4089]) );
  DFF ram_reg_1536__0_ ( .D(n8329), .CP(wclk), .Q(ram[4088]) );
  DFF ram_reg_1540__7_ ( .D(n8304), .CP(wclk), .Q(ram[4063]) );
  DFF ram_reg_1540__6_ ( .D(n8303), .CP(wclk), .Q(ram[4062]) );
  DFF ram_reg_1540__5_ ( .D(n8302), .CP(wclk), .Q(ram[4061]) );
  DFF ram_reg_1540__4_ ( .D(n8301), .CP(wclk), .Q(ram[4060]) );
  DFF ram_reg_1540__3_ ( .D(n8300), .CP(wclk), .Q(ram[4059]) );
  DFF ram_reg_1540__2_ ( .D(n8299), .CP(wclk), .Q(ram[4058]) );
  DFF ram_reg_1540__1_ ( .D(n8298), .CP(wclk), .Q(ram[4057]) );
  DFF ram_reg_1540__0_ ( .D(n8297), .CP(wclk), .Q(ram[4056]) );
  DFF ram_reg_1548__7_ ( .D(n8240), .CP(wclk), .Q(ram[3999]) );
  DFF ram_reg_1548__6_ ( .D(n8239), .CP(wclk), .Q(ram[3998]) );
  DFF ram_reg_1548__5_ ( .D(n8238), .CP(wclk), .Q(ram[3997]) );
  DFF ram_reg_1548__4_ ( .D(n8237), .CP(wclk), .Q(ram[3996]) );
  DFF ram_reg_1548__3_ ( .D(n8236), .CP(wclk), .Q(ram[3995]) );
  DFF ram_reg_1548__2_ ( .D(n8235), .CP(wclk), .Q(ram[3994]) );
  DFF ram_reg_1548__1_ ( .D(n8234), .CP(wclk), .Q(ram[3993]) );
  DFF ram_reg_1548__0_ ( .D(n8233), .CP(wclk), .Q(ram[3992]) );
  DFF ram_reg_1552__7_ ( .D(n8208), .CP(wclk), .Q(ram[3967]) );
  DFF ram_reg_1552__6_ ( .D(n8207), .CP(wclk), .Q(ram[3966]) );
  DFF ram_reg_1552__5_ ( .D(n8206), .CP(wclk), .Q(ram[3965]) );
  DFF ram_reg_1552__4_ ( .D(n8205), .CP(wclk), .Q(ram[3964]) );
  DFF ram_reg_1552__3_ ( .D(n8204), .CP(wclk), .Q(ram[3963]) );
  DFF ram_reg_1552__2_ ( .D(n8203), .CP(wclk), .Q(ram[3962]) );
  DFF ram_reg_1552__1_ ( .D(n8202), .CP(wclk), .Q(ram[3961]) );
  DFF ram_reg_1552__0_ ( .D(n8201), .CP(wclk), .Q(ram[3960]) );
  DFF ram_reg_1556__7_ ( .D(n8176), .CP(wclk), .Q(ram[3935]) );
  DFF ram_reg_1556__6_ ( .D(n8175), .CP(wclk), .Q(ram[3934]) );
  DFF ram_reg_1556__5_ ( .D(n8174), .CP(wclk), .Q(ram[3933]) );
  DFF ram_reg_1556__4_ ( .D(n8173), .CP(wclk), .Q(ram[3932]) );
  DFF ram_reg_1556__3_ ( .D(n8172), .CP(wclk), .Q(ram[3931]) );
  DFF ram_reg_1556__2_ ( .D(n8171), .CP(wclk), .Q(ram[3930]) );
  DFF ram_reg_1556__1_ ( .D(n8170), .CP(wclk), .Q(ram[3929]) );
  DFF ram_reg_1556__0_ ( .D(n8169), .CP(wclk), .Q(ram[3928]) );
  DFF ram_reg_1560__7_ ( .D(n8144), .CP(wclk), .Q(ram[3903]) );
  DFF ram_reg_1560__6_ ( .D(n8143), .CP(wclk), .Q(ram[3902]) );
  DFF ram_reg_1560__5_ ( .D(n8142), .CP(wclk), .Q(ram[3901]) );
  DFF ram_reg_1560__4_ ( .D(n8141), .CP(wclk), .Q(ram[3900]) );
  DFF ram_reg_1560__3_ ( .D(n8140), .CP(wclk), .Q(ram[3899]) );
  DFF ram_reg_1560__2_ ( .D(n8139), .CP(wclk), .Q(ram[3898]) );
  DFF ram_reg_1560__1_ ( .D(n8138), .CP(wclk), .Q(ram[3897]) );
  DFF ram_reg_1560__0_ ( .D(n8137), .CP(wclk), .Q(ram[3896]) );
  DFF ram_reg_1564__7_ ( .D(n8112), .CP(wclk), .Q(ram[3871]) );
  DFF ram_reg_1564__6_ ( .D(n8111), .CP(wclk), .Q(ram[3870]) );
  DFF ram_reg_1564__5_ ( .D(n8110), .CP(wclk), .Q(ram[3869]) );
  DFF ram_reg_1564__4_ ( .D(n8109), .CP(wclk), .Q(ram[3868]) );
  DFF ram_reg_1564__3_ ( .D(n8108), .CP(wclk), .Q(ram[3867]) );
  DFF ram_reg_1564__2_ ( .D(n8107), .CP(wclk), .Q(ram[3866]) );
  DFF ram_reg_1564__1_ ( .D(n8106), .CP(wclk), .Q(ram[3865]) );
  DFF ram_reg_1564__0_ ( .D(n8105), .CP(wclk), .Q(ram[3864]) );
  DFF ram_reg_1568__7_ ( .D(n8080), .CP(wclk), .Q(ram[3839]) );
  DFF ram_reg_1568__6_ ( .D(n8079), .CP(wclk), .Q(ram[3838]) );
  DFF ram_reg_1568__5_ ( .D(n8078), .CP(wclk), .Q(ram[3837]) );
  DFF ram_reg_1568__4_ ( .D(n8077), .CP(wclk), .Q(ram[3836]) );
  DFF ram_reg_1568__3_ ( .D(n8076), .CP(wclk), .Q(ram[3835]) );
  DFF ram_reg_1568__2_ ( .D(n8075), .CP(wclk), .Q(ram[3834]) );
  DFF ram_reg_1568__1_ ( .D(n8074), .CP(wclk), .Q(ram[3833]) );
  DFF ram_reg_1568__0_ ( .D(n8073), .CP(wclk), .Q(ram[3832]) );
  DFF ram_reg_1572__7_ ( .D(n8048), .CP(wclk), .Q(ram[3807]) );
  DFF ram_reg_1572__6_ ( .D(n8047), .CP(wclk), .Q(ram[3806]) );
  DFF ram_reg_1572__5_ ( .D(n8046), .CP(wclk), .Q(ram[3805]) );
  DFF ram_reg_1572__4_ ( .D(n8045), .CP(wclk), .Q(ram[3804]) );
  DFF ram_reg_1572__3_ ( .D(n8044), .CP(wclk), .Q(ram[3803]) );
  DFF ram_reg_1572__2_ ( .D(n8043), .CP(wclk), .Q(ram[3802]) );
  DFF ram_reg_1572__1_ ( .D(n8042), .CP(wclk), .Q(ram[3801]) );
  DFF ram_reg_1572__0_ ( .D(n8041), .CP(wclk), .Q(ram[3800]) );
  DFF ram_reg_1584__7_ ( .D(n7952), .CP(wclk), .Q(ram[3711]) );
  DFF ram_reg_1584__6_ ( .D(n7951), .CP(wclk), .Q(ram[3710]) );
  DFF ram_reg_1584__5_ ( .D(n7950), .CP(wclk), .Q(ram[3709]) );
  DFF ram_reg_1584__4_ ( .D(n7949), .CP(wclk), .Q(ram[3708]) );
  DFF ram_reg_1584__3_ ( .D(n7948), .CP(wclk), .Q(ram[3707]) );
  DFF ram_reg_1584__2_ ( .D(n7947), .CP(wclk), .Q(ram[3706]) );
  DFF ram_reg_1584__1_ ( .D(n7946), .CP(wclk), .Q(ram[3705]) );
  DFF ram_reg_1584__0_ ( .D(n7945), .CP(wclk), .Q(ram[3704]) );
  DFF ram_reg_1588__7_ ( .D(n7920), .CP(wclk), .Q(ram[3679]) );
  DFF ram_reg_1588__6_ ( .D(n7919), .CP(wclk), .Q(ram[3678]) );
  DFF ram_reg_1588__5_ ( .D(n7918), .CP(wclk), .Q(ram[3677]) );
  DFF ram_reg_1588__4_ ( .D(n7917), .CP(wclk), .Q(ram[3676]) );
  DFF ram_reg_1588__3_ ( .D(n7916), .CP(wclk), .Q(ram[3675]) );
  DFF ram_reg_1588__2_ ( .D(n7915), .CP(wclk), .Q(ram[3674]) );
  DFF ram_reg_1588__1_ ( .D(n7914), .CP(wclk), .Q(ram[3673]) );
  DFF ram_reg_1588__0_ ( .D(n7913), .CP(wclk), .Q(ram[3672]) );
  DFF ram_reg_1600__7_ ( .D(n7824), .CP(wclk), .Q(ram[3583]) );
  DFF ram_reg_1600__6_ ( .D(n7823), .CP(wclk), .Q(ram[3582]) );
  DFF ram_reg_1600__5_ ( .D(n7822), .CP(wclk), .Q(ram[3581]) );
  DFF ram_reg_1600__4_ ( .D(n7821), .CP(wclk), .Q(ram[3580]) );
  DFF ram_reg_1600__3_ ( .D(n7820), .CP(wclk), .Q(ram[3579]) );
  DFF ram_reg_1600__2_ ( .D(n7819), .CP(wclk), .Q(ram[3578]) );
  DFF ram_reg_1600__1_ ( .D(n7818), .CP(wclk), .Q(ram[3577]) );
  DFF ram_reg_1600__0_ ( .D(n7817), .CP(wclk), .Q(ram[3576]) );
  DFF ram_reg_1604__7_ ( .D(n7792), .CP(wclk), .Q(ram[3551]) );
  DFF ram_reg_1604__6_ ( .D(n7791), .CP(wclk), .Q(ram[3550]) );
  DFF ram_reg_1604__5_ ( .D(n7790), .CP(wclk), .Q(ram[3549]) );
  DFF ram_reg_1604__4_ ( .D(n7789), .CP(wclk), .Q(ram[3548]) );
  DFF ram_reg_1604__3_ ( .D(n7788), .CP(wclk), .Q(ram[3547]) );
  DFF ram_reg_1604__2_ ( .D(n7787), .CP(wclk), .Q(ram[3546]) );
  DFF ram_reg_1604__1_ ( .D(n7786), .CP(wclk), .Q(ram[3545]) );
  DFF ram_reg_1604__0_ ( .D(n7785), .CP(wclk), .Q(ram[3544]) );
  DFF ram_reg_1608__7_ ( .D(n7760), .CP(wclk), .Q(ram[3519]) );
  DFF ram_reg_1608__6_ ( .D(n7759), .CP(wclk), .Q(ram[3518]) );
  DFF ram_reg_1608__5_ ( .D(n7758), .CP(wclk), .Q(ram[3517]) );
  DFF ram_reg_1608__4_ ( .D(n7757), .CP(wclk), .Q(ram[3516]) );
  DFF ram_reg_1608__3_ ( .D(n7756), .CP(wclk), .Q(ram[3515]) );
  DFF ram_reg_1608__2_ ( .D(n7755), .CP(wclk), .Q(ram[3514]) );
  DFF ram_reg_1608__1_ ( .D(n7754), .CP(wclk), .Q(ram[3513]) );
  DFF ram_reg_1608__0_ ( .D(n7753), .CP(wclk), .Q(ram[3512]) );
  DFF ram_reg_1612__7_ ( .D(n7728), .CP(wclk), .Q(ram[3487]) );
  DFF ram_reg_1612__6_ ( .D(n7727), .CP(wclk), .Q(ram[3486]) );
  DFF ram_reg_1612__5_ ( .D(n7726), .CP(wclk), .Q(ram[3485]) );
  DFF ram_reg_1612__4_ ( .D(n7725), .CP(wclk), .Q(ram[3484]) );
  DFF ram_reg_1612__3_ ( .D(n7724), .CP(wclk), .Q(ram[3483]) );
  DFF ram_reg_1612__2_ ( .D(n7723), .CP(wclk), .Q(ram[3482]) );
  DFF ram_reg_1612__1_ ( .D(n7722), .CP(wclk), .Q(ram[3481]) );
  DFF ram_reg_1612__0_ ( .D(n7721), .CP(wclk), .Q(ram[3480]) );
  DFF ram_reg_1616__7_ ( .D(n7696), .CP(wclk), .Q(ram[3455]) );
  DFF ram_reg_1616__6_ ( .D(n7695), .CP(wclk), .Q(ram[3454]) );
  DFF ram_reg_1616__5_ ( .D(n7694), .CP(wclk), .Q(ram[3453]) );
  DFF ram_reg_1616__4_ ( .D(n7693), .CP(wclk), .Q(ram[3452]) );
  DFF ram_reg_1616__3_ ( .D(n7692), .CP(wclk), .Q(ram[3451]) );
  DFF ram_reg_1616__2_ ( .D(n7691), .CP(wclk), .Q(ram[3450]) );
  DFF ram_reg_1616__1_ ( .D(n7690), .CP(wclk), .Q(ram[3449]) );
  DFF ram_reg_1616__0_ ( .D(n7689), .CP(wclk), .Q(ram[3448]) );
  DFF ram_reg_1620__7_ ( .D(n7664), .CP(wclk), .Q(ram[3423]) );
  DFF ram_reg_1620__6_ ( .D(n7663), .CP(wclk), .Q(ram[3422]) );
  DFF ram_reg_1620__5_ ( .D(n7662), .CP(wclk), .Q(ram[3421]) );
  DFF ram_reg_1620__4_ ( .D(n7661), .CP(wclk), .Q(ram[3420]) );
  DFF ram_reg_1620__3_ ( .D(n7660), .CP(wclk), .Q(ram[3419]) );
  DFF ram_reg_1620__2_ ( .D(n7659), .CP(wclk), .Q(ram[3418]) );
  DFF ram_reg_1620__1_ ( .D(n7658), .CP(wclk), .Q(ram[3417]) );
  DFF ram_reg_1620__0_ ( .D(n7657), .CP(wclk), .Q(ram[3416]) );
  DFF ram_reg_1624__7_ ( .D(n7632), .CP(wclk), .Q(ram[3391]) );
  DFF ram_reg_1624__6_ ( .D(n7631), .CP(wclk), .Q(ram[3390]) );
  DFF ram_reg_1624__5_ ( .D(n7630), .CP(wclk), .Q(ram[3389]) );
  DFF ram_reg_1624__4_ ( .D(n7629), .CP(wclk), .Q(ram[3388]) );
  DFF ram_reg_1624__3_ ( .D(n7628), .CP(wclk), .Q(ram[3387]) );
  DFF ram_reg_1624__2_ ( .D(n7627), .CP(wclk), .Q(ram[3386]) );
  DFF ram_reg_1624__1_ ( .D(n7626), .CP(wclk), .Q(ram[3385]) );
  DFF ram_reg_1624__0_ ( .D(n7625), .CP(wclk), .Q(ram[3384]) );
  DFF ram_reg_1628__7_ ( .D(n7600), .CP(wclk), .Q(ram[3359]) );
  DFF ram_reg_1628__6_ ( .D(n7599), .CP(wclk), .Q(ram[3358]) );
  DFF ram_reg_1628__5_ ( .D(n7598), .CP(wclk), .Q(ram[3357]) );
  DFF ram_reg_1628__4_ ( .D(n7597), .CP(wclk), .Q(ram[3356]) );
  DFF ram_reg_1628__3_ ( .D(n7596), .CP(wclk), .Q(ram[3355]) );
  DFF ram_reg_1628__2_ ( .D(n7595), .CP(wclk), .Q(ram[3354]) );
  DFF ram_reg_1628__1_ ( .D(n7594), .CP(wclk), .Q(ram[3353]) );
  DFF ram_reg_1628__0_ ( .D(n7593), .CP(wclk), .Q(ram[3352]) );
  DFF ram_reg_1632__7_ ( .D(n7568), .CP(wclk), .Q(ram[3327]) );
  DFF ram_reg_1632__6_ ( .D(n7567), .CP(wclk), .Q(ram[3326]) );
  DFF ram_reg_1632__5_ ( .D(n7566), .CP(wclk), .Q(ram[3325]) );
  DFF ram_reg_1632__4_ ( .D(n7565), .CP(wclk), .Q(ram[3324]) );
  DFF ram_reg_1632__3_ ( .D(n7564), .CP(wclk), .Q(ram[3323]) );
  DFF ram_reg_1632__2_ ( .D(n7563), .CP(wclk), .Q(ram[3322]) );
  DFF ram_reg_1632__1_ ( .D(n7562), .CP(wclk), .Q(ram[3321]) );
  DFF ram_reg_1632__0_ ( .D(n7561), .CP(wclk), .Q(ram[3320]) );
  DFF ram_reg_1636__7_ ( .D(n7536), .CP(wclk), .Q(ram[3295]) );
  DFF ram_reg_1636__6_ ( .D(n7535), .CP(wclk), .Q(ram[3294]) );
  DFF ram_reg_1636__5_ ( .D(n7534), .CP(wclk), .Q(ram[3293]) );
  DFF ram_reg_1636__4_ ( .D(n7533), .CP(wclk), .Q(ram[3292]) );
  DFF ram_reg_1636__3_ ( .D(n7532), .CP(wclk), .Q(ram[3291]) );
  DFF ram_reg_1636__2_ ( .D(n7531), .CP(wclk), .Q(ram[3290]) );
  DFF ram_reg_1636__1_ ( .D(n7530), .CP(wclk), .Q(ram[3289]) );
  DFF ram_reg_1636__0_ ( .D(n7529), .CP(wclk), .Q(ram[3288]) );
  DFF ram_reg_1640__7_ ( .D(n7504), .CP(wclk), .Q(ram[3263]) );
  DFF ram_reg_1640__6_ ( .D(n7503), .CP(wclk), .Q(ram[3262]) );
  DFF ram_reg_1640__5_ ( .D(n7502), .CP(wclk), .Q(ram[3261]) );
  DFF ram_reg_1640__4_ ( .D(n7501), .CP(wclk), .Q(ram[3260]) );
  DFF ram_reg_1640__3_ ( .D(n7500), .CP(wclk), .Q(ram[3259]) );
  DFF ram_reg_1640__2_ ( .D(n7499), .CP(wclk), .Q(ram[3258]) );
  DFF ram_reg_1640__1_ ( .D(n7498), .CP(wclk), .Q(ram[3257]) );
  DFF ram_reg_1640__0_ ( .D(n7497), .CP(wclk), .Q(ram[3256]) );
  DFF ram_reg_1644__7_ ( .D(n7472), .CP(wclk), .Q(ram[3231]) );
  DFF ram_reg_1644__6_ ( .D(n7471), .CP(wclk), .Q(ram[3230]) );
  DFF ram_reg_1644__5_ ( .D(n7470), .CP(wclk), .Q(ram[3229]) );
  DFF ram_reg_1644__4_ ( .D(n7469), .CP(wclk), .Q(ram[3228]) );
  DFF ram_reg_1644__3_ ( .D(n7468), .CP(wclk), .Q(ram[3227]) );
  DFF ram_reg_1644__2_ ( .D(n7467), .CP(wclk), .Q(ram[3226]) );
  DFF ram_reg_1644__1_ ( .D(n7466), .CP(wclk), .Q(ram[3225]) );
  DFF ram_reg_1644__0_ ( .D(n7465), .CP(wclk), .Q(ram[3224]) );
  DFF ram_reg_1648__7_ ( .D(n7440), .CP(wclk), .Q(ram[3199]) );
  DFF ram_reg_1648__6_ ( .D(n7439), .CP(wclk), .Q(ram[3198]) );
  DFF ram_reg_1648__5_ ( .D(n7438), .CP(wclk), .Q(ram[3197]) );
  DFF ram_reg_1648__4_ ( .D(n7437), .CP(wclk), .Q(ram[3196]) );
  DFF ram_reg_1648__3_ ( .D(n7436), .CP(wclk), .Q(ram[3195]) );
  DFF ram_reg_1648__2_ ( .D(n7435), .CP(wclk), .Q(ram[3194]) );
  DFF ram_reg_1648__1_ ( .D(n7434), .CP(wclk), .Q(ram[3193]) );
  DFF ram_reg_1648__0_ ( .D(n7433), .CP(wclk), .Q(ram[3192]) );
  DFF ram_reg_1652__7_ ( .D(n7408), .CP(wclk), .Q(ram[3167]) );
  DFF ram_reg_1652__6_ ( .D(n7407), .CP(wclk), .Q(ram[3166]) );
  DFF ram_reg_1652__5_ ( .D(n7406), .CP(wclk), .Q(ram[3165]) );
  DFF ram_reg_1652__4_ ( .D(n7405), .CP(wclk), .Q(ram[3164]) );
  DFF ram_reg_1652__3_ ( .D(n7404), .CP(wclk), .Q(ram[3163]) );
  DFF ram_reg_1652__2_ ( .D(n7403), .CP(wclk), .Q(ram[3162]) );
  DFF ram_reg_1652__1_ ( .D(n7402), .CP(wclk), .Q(ram[3161]) );
  DFF ram_reg_1652__0_ ( .D(n7401), .CP(wclk), .Q(ram[3160]) );
  DFF ram_reg_1656__7_ ( .D(n7376), .CP(wclk), .Q(ram[3135]) );
  DFF ram_reg_1656__6_ ( .D(n7375), .CP(wclk), .Q(ram[3134]) );
  DFF ram_reg_1656__5_ ( .D(n7374), .CP(wclk), .Q(ram[3133]) );
  DFF ram_reg_1656__4_ ( .D(n7373), .CP(wclk), .Q(ram[3132]) );
  DFF ram_reg_1656__3_ ( .D(n7372), .CP(wclk), .Q(ram[3131]) );
  DFF ram_reg_1656__2_ ( .D(n7371), .CP(wclk), .Q(ram[3130]) );
  DFF ram_reg_1656__1_ ( .D(n7370), .CP(wclk), .Q(ram[3129]) );
  DFF ram_reg_1656__0_ ( .D(n7369), .CP(wclk), .Q(ram[3128]) );
  DFF ram_reg_1660__7_ ( .D(n7344), .CP(wclk), .Q(ram[3103]) );
  DFF ram_reg_1660__6_ ( .D(n7343), .CP(wclk), .Q(ram[3102]) );
  DFF ram_reg_1660__5_ ( .D(n7342), .CP(wclk), .Q(ram[3101]) );
  DFF ram_reg_1660__4_ ( .D(n7341), .CP(wclk), .Q(ram[3100]) );
  DFF ram_reg_1660__3_ ( .D(n7340), .CP(wclk), .Q(ram[3099]) );
  DFF ram_reg_1660__2_ ( .D(n7339), .CP(wclk), .Q(ram[3098]) );
  DFF ram_reg_1660__1_ ( .D(n7338), .CP(wclk), .Q(ram[3097]) );
  DFF ram_reg_1660__0_ ( .D(n7337), .CP(wclk), .Q(ram[3096]) );
  DFF ram_reg_1668__7_ ( .D(n7280), .CP(wclk), .Q(ram[3039]) );
  DFF ram_reg_1668__6_ ( .D(n7279), .CP(wclk), .Q(ram[3038]) );
  DFF ram_reg_1668__5_ ( .D(n7278), .CP(wclk), .Q(ram[3037]) );
  DFF ram_reg_1668__4_ ( .D(n7277), .CP(wclk), .Q(ram[3036]) );
  DFF ram_reg_1668__3_ ( .D(n7276), .CP(wclk), .Q(ram[3035]) );
  DFF ram_reg_1668__2_ ( .D(n7275), .CP(wclk), .Q(ram[3034]) );
  DFF ram_reg_1668__1_ ( .D(n7274), .CP(wclk), .Q(ram[3033]) );
  DFF ram_reg_1668__0_ ( .D(n7273), .CP(wclk), .Q(ram[3032]) );
  DFF ram_reg_1680__7_ ( .D(n7184), .CP(wclk), .Q(ram[2943]) );
  DFF ram_reg_1680__6_ ( .D(n7183), .CP(wclk), .Q(ram[2942]) );
  DFF ram_reg_1680__5_ ( .D(n7182), .CP(wclk), .Q(ram[2941]) );
  DFF ram_reg_1680__4_ ( .D(n7181), .CP(wclk), .Q(ram[2940]) );
  DFF ram_reg_1680__3_ ( .D(n7180), .CP(wclk), .Q(ram[2939]) );
  DFF ram_reg_1680__2_ ( .D(n7179), .CP(wclk), .Q(ram[2938]) );
  DFF ram_reg_1680__1_ ( .D(n7178), .CP(wclk), .Q(ram[2937]) );
  DFF ram_reg_1680__0_ ( .D(n7177), .CP(wclk), .Q(ram[2936]) );
  DFF ram_reg_1684__7_ ( .D(n7152), .CP(wclk), .Q(ram[2911]) );
  DFF ram_reg_1684__6_ ( .D(n7151), .CP(wclk), .Q(ram[2910]) );
  DFF ram_reg_1684__5_ ( .D(n7150), .CP(wclk), .Q(ram[2909]) );
  DFF ram_reg_1684__4_ ( .D(n7149), .CP(wclk), .Q(ram[2908]) );
  DFF ram_reg_1684__3_ ( .D(n7148), .CP(wclk), .Q(ram[2907]) );
  DFF ram_reg_1684__2_ ( .D(n7147), .CP(wclk), .Q(ram[2906]) );
  DFF ram_reg_1684__1_ ( .D(n7146), .CP(wclk), .Q(ram[2905]) );
  DFF ram_reg_1684__0_ ( .D(n7145), .CP(wclk), .Q(ram[2904]) );
  DFF ram_reg_1700__7_ ( .D(n7024), .CP(wclk), .Q(ram[2783]) );
  DFF ram_reg_1700__6_ ( .D(n7023), .CP(wclk), .Q(ram[2782]) );
  DFF ram_reg_1700__5_ ( .D(n7022), .CP(wclk), .Q(ram[2781]) );
  DFF ram_reg_1700__4_ ( .D(n7021), .CP(wclk), .Q(ram[2780]) );
  DFF ram_reg_1700__3_ ( .D(n7020), .CP(wclk), .Q(ram[2779]) );
  DFF ram_reg_1700__2_ ( .D(n7019), .CP(wclk), .Q(ram[2778]) );
  DFF ram_reg_1700__1_ ( .D(n7018), .CP(wclk), .Q(ram[2777]) );
  DFF ram_reg_1700__0_ ( .D(n7017), .CP(wclk), .Q(ram[2776]) );
  DFF ram_reg_1716__7_ ( .D(n6896), .CP(wclk), .Q(ram[2655]) );
  DFF ram_reg_1716__6_ ( .D(n6895), .CP(wclk), .Q(ram[2654]) );
  DFF ram_reg_1716__5_ ( .D(n6894), .CP(wclk), .Q(ram[2653]) );
  DFF ram_reg_1716__4_ ( .D(n6893), .CP(wclk), .Q(ram[2652]) );
  DFF ram_reg_1716__3_ ( .D(n6892), .CP(wclk), .Q(ram[2651]) );
  DFF ram_reg_1716__2_ ( .D(n6891), .CP(wclk), .Q(ram[2650]) );
  DFF ram_reg_1716__1_ ( .D(n6890), .CP(wclk), .Q(ram[2649]) );
  DFF ram_reg_1716__0_ ( .D(n6889), .CP(wclk), .Q(ram[2648]) );
  DFF ram_reg_1728__7_ ( .D(n6800), .CP(wclk), .Q(ram[2559]) );
  DFF ram_reg_1728__6_ ( .D(n6799), .CP(wclk), .Q(ram[2558]) );
  DFF ram_reg_1728__5_ ( .D(n6798), .CP(wclk), .Q(ram[2557]) );
  DFF ram_reg_1728__4_ ( .D(n6797), .CP(wclk), .Q(ram[2556]) );
  DFF ram_reg_1728__3_ ( .D(n6796), .CP(wclk), .Q(ram[2555]) );
  DFF ram_reg_1728__2_ ( .D(n6795), .CP(wclk), .Q(ram[2554]) );
  DFF ram_reg_1728__1_ ( .D(n6794), .CP(wclk), .Q(ram[2553]) );
  DFF ram_reg_1728__0_ ( .D(n6793), .CP(wclk), .Q(ram[2552]) );
  DFF ram_reg_1732__7_ ( .D(n6768), .CP(wclk), .Q(ram[2527]) );
  DFF ram_reg_1732__6_ ( .D(n6767), .CP(wclk), .Q(ram[2526]) );
  DFF ram_reg_1732__5_ ( .D(n6766), .CP(wclk), .Q(ram[2525]) );
  DFF ram_reg_1732__4_ ( .D(n6765), .CP(wclk), .Q(ram[2524]) );
  DFF ram_reg_1732__3_ ( .D(n6764), .CP(wclk), .Q(ram[2523]) );
  DFF ram_reg_1732__2_ ( .D(n6763), .CP(wclk), .Q(ram[2522]) );
  DFF ram_reg_1732__1_ ( .D(n6762), .CP(wclk), .Q(ram[2521]) );
  DFF ram_reg_1732__0_ ( .D(n6761), .CP(wclk), .Q(ram[2520]) );
  DFF ram_reg_1744__7_ ( .D(n6672), .CP(wclk), .Q(ram[2431]) );
  DFF ram_reg_1744__6_ ( .D(n6671), .CP(wclk), .Q(ram[2430]) );
  DFF ram_reg_1744__5_ ( .D(n6670), .CP(wclk), .Q(ram[2429]) );
  DFF ram_reg_1744__4_ ( .D(n6669), .CP(wclk), .Q(ram[2428]) );
  DFF ram_reg_1744__3_ ( .D(n6668), .CP(wclk), .Q(ram[2427]) );
  DFF ram_reg_1744__2_ ( .D(n6667), .CP(wclk), .Q(ram[2426]) );
  DFF ram_reg_1744__1_ ( .D(n6666), .CP(wclk), .Q(ram[2425]) );
  DFF ram_reg_1744__0_ ( .D(n6665), .CP(wclk), .Q(ram[2424]) );
  DFF ram_reg_1748__7_ ( .D(n6640), .CP(wclk), .Q(ram[2399]) );
  DFF ram_reg_1748__6_ ( .D(n6639), .CP(wclk), .Q(ram[2398]) );
  DFF ram_reg_1748__5_ ( .D(n6638), .CP(wclk), .Q(ram[2397]) );
  DFF ram_reg_1748__4_ ( .D(n6637), .CP(wclk), .Q(ram[2396]) );
  DFF ram_reg_1748__3_ ( .D(n6636), .CP(wclk), .Q(ram[2395]) );
  DFF ram_reg_1748__2_ ( .D(n6635), .CP(wclk), .Q(ram[2394]) );
  DFF ram_reg_1748__1_ ( .D(n6634), .CP(wclk), .Q(ram[2393]) );
  DFF ram_reg_1748__0_ ( .D(n6633), .CP(wclk), .Q(ram[2392]) );
  DFF ram_reg_1756__7_ ( .D(n6576), .CP(wclk), .Q(ram[2335]) );
  DFF ram_reg_1756__6_ ( .D(n6575), .CP(wclk), .Q(ram[2334]) );
  DFF ram_reg_1756__5_ ( .D(n6574), .CP(wclk), .Q(ram[2333]) );
  DFF ram_reg_1756__4_ ( .D(n6573), .CP(wclk), .Q(ram[2332]) );
  DFF ram_reg_1756__3_ ( .D(n6572), .CP(wclk), .Q(ram[2331]) );
  DFF ram_reg_1756__2_ ( .D(n6571), .CP(wclk), .Q(ram[2330]) );
  DFF ram_reg_1756__1_ ( .D(n6570), .CP(wclk), .Q(ram[2329]) );
  DFF ram_reg_1756__0_ ( .D(n6569), .CP(wclk), .Q(ram[2328]) );
  DFF ram_reg_1764__7_ ( .D(n6512), .CP(wclk), .Q(ram[2271]) );
  DFF ram_reg_1764__6_ ( .D(n6511), .CP(wclk), .Q(ram[2270]) );
  DFF ram_reg_1764__5_ ( .D(n6510), .CP(wclk), .Q(ram[2269]) );
  DFF ram_reg_1764__4_ ( .D(n6509), .CP(wclk), .Q(ram[2268]) );
  DFF ram_reg_1764__3_ ( .D(n6508), .CP(wclk), .Q(ram[2267]) );
  DFF ram_reg_1764__2_ ( .D(n6507), .CP(wclk), .Q(ram[2266]) );
  DFF ram_reg_1764__1_ ( .D(n6506), .CP(wclk), .Q(ram[2265]) );
  DFF ram_reg_1764__0_ ( .D(n6505), .CP(wclk), .Q(ram[2264]) );
  DFF ram_reg_1780__7_ ( .D(n6384), .CP(wclk), .Q(ram[2143]) );
  DFF ram_reg_1780__6_ ( .D(n6383), .CP(wclk), .Q(ram[2142]) );
  DFF ram_reg_1780__5_ ( .D(n6382), .CP(wclk), .Q(ram[2141]) );
  DFF ram_reg_1780__4_ ( .D(n6381), .CP(wclk), .Q(ram[2140]) );
  DFF ram_reg_1780__3_ ( .D(n6380), .CP(wclk), .Q(ram[2139]) );
  DFF ram_reg_1780__2_ ( .D(n6379), .CP(wclk), .Q(ram[2138]) );
  DFF ram_reg_1780__1_ ( .D(n6378), .CP(wclk), .Q(ram[2137]) );
  DFF ram_reg_1780__0_ ( .D(n6377), .CP(wclk), .Q(ram[2136]) );
  DFF ram_reg_1792__7_ ( .D(n6288), .CP(wclk), .Q(ram[2047]) );
  DFF ram_reg_1792__6_ ( .D(n6287), .CP(wclk), .Q(ram[2046]) );
  DFF ram_reg_1792__5_ ( .D(n6286), .CP(wclk), .Q(ram[2045]) );
  DFF ram_reg_1792__4_ ( .D(n6285), .CP(wclk), .Q(ram[2044]) );
  DFF ram_reg_1792__3_ ( .D(n6284), .CP(wclk), .Q(ram[2043]) );
  DFF ram_reg_1792__2_ ( .D(n6283), .CP(wclk), .Q(ram[2042]) );
  DFF ram_reg_1792__1_ ( .D(n6282), .CP(wclk), .Q(ram[2041]) );
  DFF ram_reg_1792__0_ ( .D(n6281), .CP(wclk), .Q(ram[2040]) );
  DFF ram_reg_1796__7_ ( .D(n6256), .CP(wclk), .Q(ram[2015]) );
  DFF ram_reg_1796__6_ ( .D(n6255), .CP(wclk), .Q(ram[2014]) );
  DFF ram_reg_1796__5_ ( .D(n6254), .CP(wclk), .Q(ram[2013]) );
  DFF ram_reg_1796__4_ ( .D(n6253), .CP(wclk), .Q(ram[2012]) );
  DFF ram_reg_1796__3_ ( .D(n6252), .CP(wclk), .Q(ram[2011]) );
  DFF ram_reg_1796__2_ ( .D(n6251), .CP(wclk), .Q(ram[2010]) );
  DFF ram_reg_1796__1_ ( .D(n6250), .CP(wclk), .Q(ram[2009]) );
  DFF ram_reg_1796__0_ ( .D(n6249), .CP(wclk), .Q(ram[2008]) );
  DFF ram_reg_1804__7_ ( .D(n6192), .CP(wclk), .Q(ram[1951]) );
  DFF ram_reg_1804__6_ ( .D(n6191), .CP(wclk), .Q(ram[1950]) );
  DFF ram_reg_1804__5_ ( .D(n6190), .CP(wclk), .Q(ram[1949]) );
  DFF ram_reg_1804__4_ ( .D(n6189), .CP(wclk), .Q(ram[1948]) );
  DFF ram_reg_1804__3_ ( .D(n6188), .CP(wclk), .Q(ram[1947]) );
  DFF ram_reg_1804__2_ ( .D(n6187), .CP(wclk), .Q(ram[1946]) );
  DFF ram_reg_1804__1_ ( .D(n6186), .CP(wclk), .Q(ram[1945]) );
  DFF ram_reg_1804__0_ ( .D(n6185), .CP(wclk), .Q(ram[1944]) );
  DFF ram_reg_1808__7_ ( .D(n6160), .CP(wclk), .Q(ram[1919]) );
  DFF ram_reg_1808__6_ ( .D(n6159), .CP(wclk), .Q(ram[1918]) );
  DFF ram_reg_1808__5_ ( .D(n6158), .CP(wclk), .Q(ram[1917]) );
  DFF ram_reg_1808__4_ ( .D(n6157), .CP(wclk), .Q(ram[1916]) );
  DFF ram_reg_1808__3_ ( .D(n6156), .CP(wclk), .Q(ram[1915]) );
  DFF ram_reg_1808__2_ ( .D(n6155), .CP(wclk), .Q(ram[1914]) );
  DFF ram_reg_1808__1_ ( .D(n6154), .CP(wclk), .Q(ram[1913]) );
  DFF ram_reg_1808__0_ ( .D(n6153), .CP(wclk), .Q(ram[1912]) );
  DFF ram_reg_1812__7_ ( .D(n6128), .CP(wclk), .Q(ram[1887]) );
  DFF ram_reg_1812__6_ ( .D(n6127), .CP(wclk), .Q(ram[1886]) );
  DFF ram_reg_1812__5_ ( .D(n6126), .CP(wclk), .Q(ram[1885]) );
  DFF ram_reg_1812__4_ ( .D(n6125), .CP(wclk), .Q(ram[1884]) );
  DFF ram_reg_1812__3_ ( .D(n6124), .CP(wclk), .Q(ram[1883]) );
  DFF ram_reg_1812__2_ ( .D(n6123), .CP(wclk), .Q(ram[1882]) );
  DFF ram_reg_1812__1_ ( .D(n6122), .CP(wclk), .Q(ram[1881]) );
  DFF ram_reg_1812__0_ ( .D(n6121), .CP(wclk), .Q(ram[1880]) );
  DFF ram_reg_1816__7_ ( .D(n6096), .CP(wclk), .Q(ram[1855]) );
  DFF ram_reg_1816__6_ ( .D(n6095), .CP(wclk), .Q(ram[1854]) );
  DFF ram_reg_1816__5_ ( .D(n6094), .CP(wclk), .Q(ram[1853]) );
  DFF ram_reg_1816__4_ ( .D(n6093), .CP(wclk), .Q(ram[1852]) );
  DFF ram_reg_1816__3_ ( .D(n6092), .CP(wclk), .Q(ram[1851]) );
  DFF ram_reg_1816__2_ ( .D(n6091), .CP(wclk), .Q(ram[1850]) );
  DFF ram_reg_1816__1_ ( .D(n6090), .CP(wclk), .Q(ram[1849]) );
  DFF ram_reg_1816__0_ ( .D(n6089), .CP(wclk), .Q(ram[1848]) );
  DFF ram_reg_1820__7_ ( .D(n6064), .CP(wclk), .Q(ram[1823]) );
  DFF ram_reg_1820__6_ ( .D(n6063), .CP(wclk), .Q(ram[1822]) );
  DFF ram_reg_1820__5_ ( .D(n6062), .CP(wclk), .Q(ram[1821]) );
  DFF ram_reg_1820__4_ ( .D(n6061), .CP(wclk), .Q(ram[1820]) );
  DFF ram_reg_1820__3_ ( .D(n6060), .CP(wclk), .Q(ram[1819]) );
  DFF ram_reg_1820__2_ ( .D(n6059), .CP(wclk), .Q(ram[1818]) );
  DFF ram_reg_1820__1_ ( .D(n6058), .CP(wclk), .Q(ram[1817]) );
  DFF ram_reg_1820__0_ ( .D(n6057), .CP(wclk), .Q(ram[1816]) );
  DFF ram_reg_1824__7_ ( .D(n6032), .CP(wclk), .Q(ram[1791]) );
  DFF ram_reg_1824__6_ ( .D(n6031), .CP(wclk), .Q(ram[1790]) );
  DFF ram_reg_1824__5_ ( .D(n6030), .CP(wclk), .Q(ram[1789]) );
  DFF ram_reg_1824__4_ ( .D(n6029), .CP(wclk), .Q(ram[1788]) );
  DFF ram_reg_1824__3_ ( .D(n6028), .CP(wclk), .Q(ram[1787]) );
  DFF ram_reg_1824__2_ ( .D(n6027), .CP(wclk), .Q(ram[1786]) );
  DFF ram_reg_1824__1_ ( .D(n6026), .CP(wclk), .Q(ram[1785]) );
  DFF ram_reg_1824__0_ ( .D(n6025), .CP(wclk), .Q(ram[1784]) );
  DFF ram_reg_1828__7_ ( .D(n6000), .CP(wclk), .Q(ram[1759]) );
  DFF ram_reg_1828__6_ ( .D(n5999), .CP(wclk), .Q(ram[1758]) );
  DFF ram_reg_1828__5_ ( .D(n5998), .CP(wclk), .Q(ram[1757]) );
  DFF ram_reg_1828__4_ ( .D(n5997), .CP(wclk), .Q(ram[1756]) );
  DFF ram_reg_1828__3_ ( .D(n5996), .CP(wclk), .Q(ram[1755]) );
  DFF ram_reg_1828__2_ ( .D(n5995), .CP(wclk), .Q(ram[1754]) );
  DFF ram_reg_1828__1_ ( .D(n5994), .CP(wclk), .Q(ram[1753]) );
  DFF ram_reg_1828__0_ ( .D(n5993), .CP(wclk), .Q(ram[1752]) );
  DFF ram_reg_1840__7_ ( .D(n5904), .CP(wclk), .Q(ram[1663]) );
  DFF ram_reg_1840__6_ ( .D(n5903), .CP(wclk), .Q(ram[1662]) );
  DFF ram_reg_1840__5_ ( .D(n5902), .CP(wclk), .Q(ram[1661]) );
  DFF ram_reg_1840__4_ ( .D(n5901), .CP(wclk), .Q(ram[1660]) );
  DFF ram_reg_1840__3_ ( .D(n5900), .CP(wclk), .Q(ram[1659]) );
  DFF ram_reg_1840__2_ ( .D(n5899), .CP(wclk), .Q(ram[1658]) );
  DFF ram_reg_1840__1_ ( .D(n5898), .CP(wclk), .Q(ram[1657]) );
  DFF ram_reg_1840__0_ ( .D(n5897), .CP(wclk), .Q(ram[1656]) );
  DFF ram_reg_1844__7_ ( .D(n5872), .CP(wclk), .Q(ram[1631]) );
  DFF ram_reg_1844__6_ ( .D(n5871), .CP(wclk), .Q(ram[1630]) );
  DFF ram_reg_1844__5_ ( .D(n5870), .CP(wclk), .Q(ram[1629]) );
  DFF ram_reg_1844__4_ ( .D(n5869), .CP(wclk), .Q(ram[1628]) );
  DFF ram_reg_1844__3_ ( .D(n5868), .CP(wclk), .Q(ram[1627]) );
  DFF ram_reg_1844__2_ ( .D(n5867), .CP(wclk), .Q(ram[1626]) );
  DFF ram_reg_1844__1_ ( .D(n5866), .CP(wclk), .Q(ram[1625]) );
  DFF ram_reg_1844__0_ ( .D(n5865), .CP(wclk), .Q(ram[1624]) );
  DFF ram_reg_1856__7_ ( .D(n5776), .CP(wclk), .Q(ram[1535]) );
  DFF ram_reg_1856__6_ ( .D(n5775), .CP(wclk), .Q(ram[1534]) );
  DFF ram_reg_1856__5_ ( .D(n5774), .CP(wclk), .Q(ram[1533]) );
  DFF ram_reg_1856__4_ ( .D(n5773), .CP(wclk), .Q(ram[1532]) );
  DFF ram_reg_1856__3_ ( .D(n5772), .CP(wclk), .Q(ram[1531]) );
  DFF ram_reg_1856__2_ ( .D(n5771), .CP(wclk), .Q(ram[1530]) );
  DFF ram_reg_1856__1_ ( .D(n5770), .CP(wclk), .Q(ram[1529]) );
  DFF ram_reg_1856__0_ ( .D(n5769), .CP(wclk), .Q(ram[1528]) );
  DFF ram_reg_1860__7_ ( .D(n5744), .CP(wclk), .Q(ram[1503]) );
  DFF ram_reg_1860__6_ ( .D(n5743), .CP(wclk), .Q(ram[1502]) );
  DFF ram_reg_1860__5_ ( .D(n5742), .CP(wclk), .Q(ram[1501]) );
  DFF ram_reg_1860__4_ ( .D(n5741), .CP(wclk), .Q(ram[1500]) );
  DFF ram_reg_1860__3_ ( .D(n5740), .CP(wclk), .Q(ram[1499]) );
  DFF ram_reg_1860__2_ ( .D(n5739), .CP(wclk), .Q(ram[1498]) );
  DFF ram_reg_1860__1_ ( .D(n5738), .CP(wclk), .Q(ram[1497]) );
  DFF ram_reg_1860__0_ ( .D(n5737), .CP(wclk), .Q(ram[1496]) );
  DFF ram_reg_1864__7_ ( .D(n5712), .CP(wclk), .Q(ram[1471]) );
  DFF ram_reg_1864__6_ ( .D(n5711), .CP(wclk), .Q(ram[1470]) );
  DFF ram_reg_1864__5_ ( .D(n5710), .CP(wclk), .Q(ram[1469]) );
  DFF ram_reg_1864__4_ ( .D(n5709), .CP(wclk), .Q(ram[1468]) );
  DFF ram_reg_1864__3_ ( .D(n5708), .CP(wclk), .Q(ram[1467]) );
  DFF ram_reg_1864__2_ ( .D(n5707), .CP(wclk), .Q(ram[1466]) );
  DFF ram_reg_1864__1_ ( .D(n5706), .CP(wclk), .Q(ram[1465]) );
  DFF ram_reg_1864__0_ ( .D(n5705), .CP(wclk), .Q(ram[1464]) );
  DFF ram_reg_1868__7_ ( .D(n5680), .CP(wclk), .Q(ram[1439]) );
  DFF ram_reg_1868__6_ ( .D(n5679), .CP(wclk), .Q(ram[1438]) );
  DFF ram_reg_1868__5_ ( .D(n5678), .CP(wclk), .Q(ram[1437]) );
  DFF ram_reg_1868__4_ ( .D(n5677), .CP(wclk), .Q(ram[1436]) );
  DFF ram_reg_1868__3_ ( .D(n5676), .CP(wclk), .Q(ram[1435]) );
  DFF ram_reg_1868__2_ ( .D(n5675), .CP(wclk), .Q(ram[1434]) );
  DFF ram_reg_1868__1_ ( .D(n5674), .CP(wclk), .Q(ram[1433]) );
  DFF ram_reg_1868__0_ ( .D(n5673), .CP(wclk), .Q(ram[1432]) );
  DFF ram_reg_1872__7_ ( .D(n5648), .CP(wclk), .Q(ram[1407]) );
  DFF ram_reg_1872__6_ ( .D(n5647), .CP(wclk), .Q(ram[1406]) );
  DFF ram_reg_1872__5_ ( .D(n5646), .CP(wclk), .Q(ram[1405]) );
  DFF ram_reg_1872__4_ ( .D(n5645), .CP(wclk), .Q(ram[1404]) );
  DFF ram_reg_1872__3_ ( .D(n5644), .CP(wclk), .Q(ram[1403]) );
  DFF ram_reg_1872__2_ ( .D(n5643), .CP(wclk), .Q(ram[1402]) );
  DFF ram_reg_1872__1_ ( .D(n5642), .CP(wclk), .Q(ram[1401]) );
  DFF ram_reg_1872__0_ ( .D(n5641), .CP(wclk), .Q(ram[1400]) );
  DFF ram_reg_1876__7_ ( .D(n5616), .CP(wclk), .Q(ram[1375]) );
  DFF ram_reg_1876__6_ ( .D(n5615), .CP(wclk), .Q(ram[1374]) );
  DFF ram_reg_1876__5_ ( .D(n5614), .CP(wclk), .Q(ram[1373]) );
  DFF ram_reg_1876__4_ ( .D(n5613), .CP(wclk), .Q(ram[1372]) );
  DFF ram_reg_1876__3_ ( .D(n5612), .CP(wclk), .Q(ram[1371]) );
  DFF ram_reg_1876__2_ ( .D(n5611), .CP(wclk), .Q(ram[1370]) );
  DFF ram_reg_1876__1_ ( .D(n5610), .CP(wclk), .Q(ram[1369]) );
  DFF ram_reg_1876__0_ ( .D(n5609), .CP(wclk), .Q(ram[1368]) );
  DFF ram_reg_1880__7_ ( .D(n5584), .CP(wclk), .Q(ram[1343]) );
  DFF ram_reg_1880__6_ ( .D(n5583), .CP(wclk), .Q(ram[1342]) );
  DFF ram_reg_1880__5_ ( .D(n5582), .CP(wclk), .Q(ram[1341]) );
  DFF ram_reg_1880__4_ ( .D(n5581), .CP(wclk), .Q(ram[1340]) );
  DFF ram_reg_1880__3_ ( .D(n5580), .CP(wclk), .Q(ram[1339]) );
  DFF ram_reg_1880__2_ ( .D(n5579), .CP(wclk), .Q(ram[1338]) );
  DFF ram_reg_1880__1_ ( .D(n5578), .CP(wclk), .Q(ram[1337]) );
  DFF ram_reg_1880__0_ ( .D(n5577), .CP(wclk), .Q(ram[1336]) );
  DFF ram_reg_1884__7_ ( .D(n5552), .CP(wclk), .Q(ram[1311]) );
  DFF ram_reg_1884__6_ ( .D(n5551), .CP(wclk), .Q(ram[1310]) );
  DFF ram_reg_1884__5_ ( .D(n5550), .CP(wclk), .Q(ram[1309]) );
  DFF ram_reg_1884__4_ ( .D(n5549), .CP(wclk), .Q(ram[1308]) );
  DFF ram_reg_1884__3_ ( .D(n5548), .CP(wclk), .Q(ram[1307]) );
  DFF ram_reg_1884__2_ ( .D(n5547), .CP(wclk), .Q(ram[1306]) );
  DFF ram_reg_1884__1_ ( .D(n5546), .CP(wclk), .Q(ram[1305]) );
  DFF ram_reg_1884__0_ ( .D(n5545), .CP(wclk), .Q(ram[1304]) );
  DFF ram_reg_1888__7_ ( .D(n5520), .CP(wclk), .Q(ram[1279]) );
  DFF ram_reg_1888__6_ ( .D(n5519), .CP(wclk), .Q(ram[1278]) );
  DFF ram_reg_1888__5_ ( .D(n5518), .CP(wclk), .Q(ram[1277]) );
  DFF ram_reg_1888__4_ ( .D(n5517), .CP(wclk), .Q(ram[1276]) );
  DFF ram_reg_1888__3_ ( .D(n5516), .CP(wclk), .Q(ram[1275]) );
  DFF ram_reg_1888__2_ ( .D(n5515), .CP(wclk), .Q(ram[1274]) );
  DFF ram_reg_1888__1_ ( .D(n5514), .CP(wclk), .Q(ram[1273]) );
  DFF ram_reg_1888__0_ ( .D(n5513), .CP(wclk), .Q(ram[1272]) );
  DFF ram_reg_1892__7_ ( .D(n5488), .CP(wclk), .Q(ram[1247]) );
  DFF ram_reg_1892__6_ ( .D(n5487), .CP(wclk), .Q(ram[1246]) );
  DFF ram_reg_1892__5_ ( .D(n5486), .CP(wclk), .Q(ram[1245]) );
  DFF ram_reg_1892__4_ ( .D(n5485), .CP(wclk), .Q(ram[1244]) );
  DFF ram_reg_1892__3_ ( .D(n5484), .CP(wclk), .Q(ram[1243]) );
  DFF ram_reg_1892__2_ ( .D(n5483), .CP(wclk), .Q(ram[1242]) );
  DFF ram_reg_1892__1_ ( .D(n5482), .CP(wclk), .Q(ram[1241]) );
  DFF ram_reg_1892__0_ ( .D(n5481), .CP(wclk), .Q(ram[1240]) );
  DFF ram_reg_1896__7_ ( .D(n5456), .CP(wclk), .Q(ram[1215]) );
  DFF ram_reg_1896__6_ ( .D(n5455), .CP(wclk), .Q(ram[1214]) );
  DFF ram_reg_1896__5_ ( .D(n5454), .CP(wclk), .Q(ram[1213]) );
  DFF ram_reg_1896__4_ ( .D(n5453), .CP(wclk), .Q(ram[1212]) );
  DFF ram_reg_1896__3_ ( .D(n5452), .CP(wclk), .Q(ram[1211]) );
  DFF ram_reg_1896__2_ ( .D(n5451), .CP(wclk), .Q(ram[1210]) );
  DFF ram_reg_1896__1_ ( .D(n5450), .CP(wclk), .Q(ram[1209]) );
  DFF ram_reg_1896__0_ ( .D(n5449), .CP(wclk), .Q(ram[1208]) );
  DFF ram_reg_1900__7_ ( .D(n5424), .CP(wclk), .Q(ram[1183]) );
  DFF ram_reg_1900__6_ ( .D(n5423), .CP(wclk), .Q(ram[1182]) );
  DFF ram_reg_1900__5_ ( .D(n5422), .CP(wclk), .Q(ram[1181]) );
  DFF ram_reg_1900__4_ ( .D(n5421), .CP(wclk), .Q(ram[1180]) );
  DFF ram_reg_1900__3_ ( .D(n5420), .CP(wclk), .Q(ram[1179]) );
  DFF ram_reg_1900__2_ ( .D(n5419), .CP(wclk), .Q(ram[1178]) );
  DFF ram_reg_1900__1_ ( .D(n5418), .CP(wclk), .Q(ram[1177]) );
  DFF ram_reg_1900__0_ ( .D(n5417), .CP(wclk), .Q(ram[1176]) );
  DFF ram_reg_1904__7_ ( .D(n5392), .CP(wclk), .Q(ram[1151]) );
  DFF ram_reg_1904__6_ ( .D(n5391), .CP(wclk), .Q(ram[1150]) );
  DFF ram_reg_1904__5_ ( .D(n5390), .CP(wclk), .Q(ram[1149]) );
  DFF ram_reg_1904__4_ ( .D(n5389), .CP(wclk), .Q(ram[1148]) );
  DFF ram_reg_1904__3_ ( .D(n5388), .CP(wclk), .Q(ram[1147]) );
  DFF ram_reg_1904__2_ ( .D(n5387), .CP(wclk), .Q(ram[1146]) );
  DFF ram_reg_1904__1_ ( .D(n5386), .CP(wclk), .Q(ram[1145]) );
  DFF ram_reg_1904__0_ ( .D(n5385), .CP(wclk), .Q(ram[1144]) );
  DFF ram_reg_1908__7_ ( .D(n5360), .CP(wclk), .Q(ram[1119]) );
  DFF ram_reg_1908__6_ ( .D(n5359), .CP(wclk), .Q(ram[1118]) );
  DFF ram_reg_1908__5_ ( .D(n5358), .CP(wclk), .Q(ram[1117]) );
  DFF ram_reg_1908__4_ ( .D(n5357), .CP(wclk), .Q(ram[1116]) );
  DFF ram_reg_1908__3_ ( .D(n5356), .CP(wclk), .Q(ram[1115]) );
  DFF ram_reg_1908__2_ ( .D(n5355), .CP(wclk), .Q(ram[1114]) );
  DFF ram_reg_1908__1_ ( .D(n5354), .CP(wclk), .Q(ram[1113]) );
  DFF ram_reg_1908__0_ ( .D(n5353), .CP(wclk), .Q(ram[1112]) );
  DFF ram_reg_1912__7_ ( .D(n5328), .CP(wclk), .Q(ram[1087]) );
  DFF ram_reg_1912__6_ ( .D(n5327), .CP(wclk), .Q(ram[1086]) );
  DFF ram_reg_1912__5_ ( .D(n5326), .CP(wclk), .Q(ram[1085]) );
  DFF ram_reg_1912__4_ ( .D(n5325), .CP(wclk), .Q(ram[1084]) );
  DFF ram_reg_1912__3_ ( .D(n5324), .CP(wclk), .Q(ram[1083]) );
  DFF ram_reg_1912__2_ ( .D(n5323), .CP(wclk), .Q(ram[1082]) );
  DFF ram_reg_1912__1_ ( .D(n5322), .CP(wclk), .Q(ram[1081]) );
  DFF ram_reg_1912__0_ ( .D(n5321), .CP(wclk), .Q(ram[1080]) );
  DFF ram_reg_1916__7_ ( .D(n5296), .CP(wclk), .Q(ram[1055]) );
  DFF ram_reg_1916__6_ ( .D(n5295), .CP(wclk), .Q(ram[1054]) );
  DFF ram_reg_1916__5_ ( .D(n5294), .CP(wclk), .Q(ram[1053]) );
  DFF ram_reg_1916__4_ ( .D(n5293), .CP(wclk), .Q(ram[1052]) );
  DFF ram_reg_1916__3_ ( .D(n5292), .CP(wclk), .Q(ram[1051]) );
  DFF ram_reg_1916__2_ ( .D(n5291), .CP(wclk), .Q(ram[1050]) );
  DFF ram_reg_1916__1_ ( .D(n5290), .CP(wclk), .Q(ram[1049]) );
  DFF ram_reg_1916__0_ ( .D(n5289), .CP(wclk), .Q(ram[1048]) );
  DFF ram_reg_1924__7_ ( .D(n5232), .CP(wclk), .Q(ram[991]) );
  DFF ram_reg_1924__6_ ( .D(n5231), .CP(wclk), .Q(ram[990]) );
  DFF ram_reg_1924__5_ ( .D(n5230), .CP(wclk), .Q(ram[989]) );
  DFF ram_reg_1924__4_ ( .D(n5229), .CP(wclk), .Q(ram[988]) );
  DFF ram_reg_1924__3_ ( .D(n5228), .CP(wclk), .Q(ram[987]) );
  DFF ram_reg_1924__2_ ( .D(n5227), .CP(wclk), .Q(ram[986]) );
  DFF ram_reg_1924__1_ ( .D(n5226), .CP(wclk), .Q(ram[985]) );
  DFF ram_reg_1924__0_ ( .D(n5225), .CP(wclk), .Q(ram[984]) );
  DFF ram_reg_1936__7_ ( .D(n5136), .CP(wclk), .Q(ram[895]) );
  DFF ram_reg_1936__6_ ( .D(n5135), .CP(wclk), .Q(ram[894]) );
  DFF ram_reg_1936__5_ ( .D(n5134), .CP(wclk), .Q(ram[893]) );
  DFF ram_reg_1936__4_ ( .D(n5133), .CP(wclk), .Q(ram[892]) );
  DFF ram_reg_1936__3_ ( .D(n5132), .CP(wclk), .Q(ram[891]) );
  DFF ram_reg_1936__2_ ( .D(n5131), .CP(wclk), .Q(ram[890]) );
  DFF ram_reg_1936__1_ ( .D(n5130), .CP(wclk), .Q(ram[889]) );
  DFF ram_reg_1936__0_ ( .D(n5129), .CP(wclk), .Q(ram[888]) );
  DFF ram_reg_1940__7_ ( .D(n5104), .CP(wclk), .Q(ram[863]) );
  DFF ram_reg_1940__6_ ( .D(n5103), .CP(wclk), .Q(ram[862]) );
  DFF ram_reg_1940__5_ ( .D(n5102), .CP(wclk), .Q(ram[861]) );
  DFF ram_reg_1940__4_ ( .D(n5101), .CP(wclk), .Q(ram[860]) );
  DFF ram_reg_1940__3_ ( .D(n5100), .CP(wclk), .Q(ram[859]) );
  DFF ram_reg_1940__2_ ( .D(n5099), .CP(wclk), .Q(ram[858]) );
  DFF ram_reg_1940__1_ ( .D(n5098), .CP(wclk), .Q(ram[857]) );
  DFF ram_reg_1940__0_ ( .D(n5097), .CP(wclk), .Q(ram[856]) );
  DFF ram_reg_1956__7_ ( .D(n4976), .CP(wclk), .Q(ram[735]) );
  DFF ram_reg_1956__6_ ( .D(n4975), .CP(wclk), .Q(ram[734]) );
  DFF ram_reg_1956__5_ ( .D(n4974), .CP(wclk), .Q(ram[733]) );
  DFF ram_reg_1956__4_ ( .D(n4973), .CP(wclk), .Q(ram[732]) );
  DFF ram_reg_1956__3_ ( .D(n4972), .CP(wclk), .Q(ram[731]) );
  DFF ram_reg_1956__2_ ( .D(n4971), .CP(wclk), .Q(ram[730]) );
  DFF ram_reg_1956__1_ ( .D(n4970), .CP(wclk), .Q(ram[729]) );
  DFF ram_reg_1956__0_ ( .D(n4969), .CP(wclk), .Q(ram[728]) );
  DFF ram_reg_1972__7_ ( .D(n4848), .CP(wclk), .Q(ram[607]) );
  DFF ram_reg_1972__6_ ( .D(n4847), .CP(wclk), .Q(ram[606]) );
  DFF ram_reg_1972__5_ ( .D(n4846), .CP(wclk), .Q(ram[605]) );
  DFF ram_reg_1972__4_ ( .D(n4845), .CP(wclk), .Q(ram[604]) );
  DFF ram_reg_1972__3_ ( .D(n4844), .CP(wclk), .Q(ram[603]) );
  DFF ram_reg_1972__2_ ( .D(n4843), .CP(wclk), .Q(ram[602]) );
  DFF ram_reg_1972__1_ ( .D(n4842), .CP(wclk), .Q(ram[601]) );
  DFF ram_reg_1972__0_ ( .D(n4841), .CP(wclk), .Q(ram[600]) );
  DFF ram_reg_1984__7_ ( .D(n4752), .CP(wclk), .Q(ram[511]) );
  DFF ram_reg_1984__6_ ( .D(n4751), .CP(wclk), .Q(ram[510]) );
  DFF ram_reg_1984__5_ ( .D(n4750), .CP(wclk), .Q(ram[509]) );
  DFF ram_reg_1984__4_ ( .D(n4749), .CP(wclk), .Q(ram[508]) );
  DFF ram_reg_1984__3_ ( .D(n4748), .CP(wclk), .Q(ram[507]) );
  DFF ram_reg_1984__2_ ( .D(n4747), .CP(wclk), .Q(ram[506]) );
  DFF ram_reg_1984__1_ ( .D(n4746), .CP(wclk), .Q(ram[505]) );
  DFF ram_reg_1984__0_ ( .D(n4745), .CP(wclk), .Q(ram[504]) );
  DFF ram_reg_1988__7_ ( .D(n4720), .CP(wclk), .Q(ram[479]) );
  DFF ram_reg_1988__6_ ( .D(n4719), .CP(wclk), .Q(ram[478]) );
  DFF ram_reg_1988__5_ ( .D(n4718), .CP(wclk), .Q(ram[477]) );
  DFF ram_reg_1988__4_ ( .D(n4717), .CP(wclk), .Q(ram[476]) );
  DFF ram_reg_1988__3_ ( .D(n4716), .CP(wclk), .Q(ram[475]) );
  DFF ram_reg_1988__2_ ( .D(n4715), .CP(wclk), .Q(ram[474]) );
  DFF ram_reg_1988__1_ ( .D(n4714), .CP(wclk), .Q(ram[473]) );
  DFF ram_reg_1988__0_ ( .D(n4713), .CP(wclk), .Q(ram[472]) );
  DFF ram_reg_2000__7_ ( .D(n4624), .CP(wclk), .Q(ram[383]) );
  DFF ram_reg_2000__6_ ( .D(n4623), .CP(wclk), .Q(ram[382]) );
  DFF ram_reg_2000__5_ ( .D(n4622), .CP(wclk), .Q(ram[381]) );
  DFF ram_reg_2000__4_ ( .D(n4621), .CP(wclk), .Q(ram[380]) );
  DFF ram_reg_2000__3_ ( .D(n4620), .CP(wclk), .Q(ram[379]) );
  DFF ram_reg_2000__2_ ( .D(n4619), .CP(wclk), .Q(ram[378]) );
  DFF ram_reg_2000__1_ ( .D(n4618), .CP(wclk), .Q(ram[377]) );
  DFF ram_reg_2000__0_ ( .D(n4617), .CP(wclk), .Q(ram[376]) );
  DFF ram_reg_2004__7_ ( .D(n4592), .CP(wclk), .Q(ram[351]) );
  DFF ram_reg_2004__6_ ( .D(n4591), .CP(wclk), .Q(ram[350]) );
  DFF ram_reg_2004__5_ ( .D(n4590), .CP(wclk), .Q(ram[349]) );
  DFF ram_reg_2004__4_ ( .D(n4589), .CP(wclk), .Q(ram[348]) );
  DFF ram_reg_2004__3_ ( .D(n4588), .CP(wclk), .Q(ram[347]) );
  DFF ram_reg_2004__2_ ( .D(n4587), .CP(wclk), .Q(ram[346]) );
  DFF ram_reg_2004__1_ ( .D(n4586), .CP(wclk), .Q(ram[345]) );
  DFF ram_reg_2004__0_ ( .D(n4585), .CP(wclk), .Q(ram[344]) );
  DFF ram_reg_2020__7_ ( .D(n4464), .CP(wclk), .Q(ram[223]) );
  DFF ram_reg_2020__6_ ( .D(n4463), .CP(wclk), .Q(ram[222]) );
  DFF ram_reg_2020__5_ ( .D(n4462), .CP(wclk), .Q(ram[221]) );
  DFF ram_reg_2020__4_ ( .D(n4461), .CP(wclk), .Q(ram[220]) );
  DFF ram_reg_2020__3_ ( .D(n4460), .CP(wclk), .Q(ram[219]) );
  DFF ram_reg_2020__2_ ( .D(n4459), .CP(wclk), .Q(ram[218]) );
  DFF ram_reg_2020__1_ ( .D(n4458), .CP(wclk), .Q(ram[217]) );
  DFF ram_reg_2020__0_ ( .D(n4457), .CP(wclk), .Q(ram[216]) );
  DFF ram_reg_2036__7_ ( .D(n4336), .CP(wclk), .Q(ram[95]) );
  DFF ram_reg_2036__6_ ( .D(n4335), .CP(wclk), .Q(ram[94]) );
  DFF ram_reg_2036__5_ ( .D(n4334), .CP(wclk), .Q(ram[93]) );
  DFF ram_reg_2036__4_ ( .D(n4333), .CP(wclk), .Q(ram[92]) );
  DFF ram_reg_2036__3_ ( .D(n4332), .CP(wclk), .Q(ram[91]) );
  DFF ram_reg_2036__2_ ( .D(n4331), .CP(wclk), .Q(ram[90]) );
  DFF ram_reg_2036__1_ ( .D(n4330), .CP(wclk), .Q(ram[89]) );
  DFF ram_reg_2036__0_ ( .D(n4329), .CP(wclk), .Q(ram[88]) );
  DFF ram_reg_2__7_ ( .D(n20608), .CP(wclk), .Q(ram[16367]) );
  DFF ram_reg_2__6_ ( .D(n20607), .CP(wclk), .Q(ram[16366]) );
  DFF ram_reg_2__5_ ( .D(n20606), .CP(wclk), .Q(ram[16365]) );
  DFF ram_reg_2__4_ ( .D(n20605), .CP(wclk), .Q(ram[16364]) );
  DFF ram_reg_2__3_ ( .D(n20604), .CP(wclk), .Q(ram[16363]) );
  DFF ram_reg_2__2_ ( .D(n20603), .CP(wclk), .Q(ram[16362]) );
  DFF ram_reg_2__1_ ( .D(n20602), .CP(wclk), .Q(ram[16361]) );
  DFF ram_reg_2__0_ ( .D(n20601), .CP(wclk), .Q(ram[16360]) );
  DFF ram_reg_6__7_ ( .D(n20576), .CP(wclk), .Q(ram[16335]) );
  DFF ram_reg_6__6_ ( .D(n20575), .CP(wclk), .Q(ram[16334]) );
  DFF ram_reg_6__5_ ( .D(n20574), .CP(wclk), .Q(ram[16333]) );
  DFF ram_reg_6__4_ ( .D(n20573), .CP(wclk), .Q(ram[16332]) );
  DFF ram_reg_6__3_ ( .D(n20572), .CP(wclk), .Q(ram[16331]) );
  DFF ram_reg_6__2_ ( .D(n20571), .CP(wclk), .Q(ram[16330]) );
  DFF ram_reg_6__1_ ( .D(n20570), .CP(wclk), .Q(ram[16329]) );
  DFF ram_reg_6__0_ ( .D(n20569), .CP(wclk), .Q(ram[16328]) );
  DFF ram_reg_10__7_ ( .D(n20544), .CP(wclk), .Q(ram[16303]) );
  DFF ram_reg_10__6_ ( .D(n20543), .CP(wclk), .Q(ram[16302]) );
  DFF ram_reg_10__5_ ( .D(n20542), .CP(wclk), .Q(ram[16301]) );
  DFF ram_reg_10__4_ ( .D(n20541), .CP(wclk), .Q(ram[16300]) );
  DFF ram_reg_10__3_ ( .D(n20540), .CP(wclk), .Q(ram[16299]) );
  DFF ram_reg_10__2_ ( .D(n20539), .CP(wclk), .Q(ram[16298]) );
  DFF ram_reg_10__1_ ( .D(n20538), .CP(wclk), .Q(ram[16297]) );
  DFF ram_reg_10__0_ ( .D(n20537), .CP(wclk), .Q(ram[16296]) );
  DFF ram_reg_14__7_ ( .D(n20512), .CP(wclk), .Q(ram[16271]) );
  DFF ram_reg_14__6_ ( .D(n20511), .CP(wclk), .Q(ram[16270]) );
  DFF ram_reg_14__5_ ( .D(n20510), .CP(wclk), .Q(ram[16269]) );
  DFF ram_reg_14__4_ ( .D(n20509), .CP(wclk), .Q(ram[16268]) );
  DFF ram_reg_14__3_ ( .D(n20508), .CP(wclk), .Q(ram[16267]) );
  DFF ram_reg_14__2_ ( .D(n20507), .CP(wclk), .Q(ram[16266]) );
  DFF ram_reg_14__1_ ( .D(n20506), .CP(wclk), .Q(ram[16265]) );
  DFF ram_reg_14__0_ ( .D(n20505), .CP(wclk), .Q(ram[16264]) );
  DFF ram_reg_18__7_ ( .D(n20480), .CP(wclk), .Q(ram[16239]) );
  DFF ram_reg_18__6_ ( .D(n20479), .CP(wclk), .Q(ram[16238]) );
  DFF ram_reg_18__5_ ( .D(n20478), .CP(wclk), .Q(ram[16237]) );
  DFF ram_reg_18__4_ ( .D(n20477), .CP(wclk), .Q(ram[16236]) );
  DFF ram_reg_18__3_ ( .D(n20476), .CP(wclk), .Q(ram[16235]) );
  DFF ram_reg_18__2_ ( .D(n20475), .CP(wclk), .Q(ram[16234]) );
  DFF ram_reg_18__1_ ( .D(n20474), .CP(wclk), .Q(ram[16233]) );
  DFF ram_reg_18__0_ ( .D(n20473), .CP(wclk), .Q(ram[16232]) );
  DFF ram_reg_22__7_ ( .D(n20448), .CP(wclk), .Q(ram[16207]) );
  DFF ram_reg_22__6_ ( .D(n20447), .CP(wclk), .Q(ram[16206]) );
  DFF ram_reg_22__5_ ( .D(n20446), .CP(wclk), .Q(ram[16205]) );
  DFF ram_reg_22__4_ ( .D(n20445), .CP(wclk), .Q(ram[16204]) );
  DFF ram_reg_22__3_ ( .D(n20444), .CP(wclk), .Q(ram[16203]) );
  DFF ram_reg_22__2_ ( .D(n20443), .CP(wclk), .Q(ram[16202]) );
  DFF ram_reg_22__1_ ( .D(n20442), .CP(wclk), .Q(ram[16201]) );
  DFF ram_reg_22__0_ ( .D(n20441), .CP(wclk), .Q(ram[16200]) );
  DFF ram_reg_26__7_ ( .D(n20416), .CP(wclk), .Q(ram[16175]) );
  DFF ram_reg_26__6_ ( .D(n20415), .CP(wclk), .Q(ram[16174]) );
  DFF ram_reg_26__5_ ( .D(n20414), .CP(wclk), .Q(ram[16173]) );
  DFF ram_reg_26__4_ ( .D(n20413), .CP(wclk), .Q(ram[16172]) );
  DFF ram_reg_26__3_ ( .D(n20412), .CP(wclk), .Q(ram[16171]) );
  DFF ram_reg_26__2_ ( .D(n20411), .CP(wclk), .Q(ram[16170]) );
  DFF ram_reg_26__1_ ( .D(n20410), .CP(wclk), .Q(ram[16169]) );
  DFF ram_reg_26__0_ ( .D(n20409), .CP(wclk), .Q(ram[16168]) );
  DFF ram_reg_30__7_ ( .D(n20384), .CP(wclk), .Q(ram[16143]) );
  DFF ram_reg_30__6_ ( .D(n20383), .CP(wclk), .Q(ram[16142]) );
  DFF ram_reg_30__5_ ( .D(n20382), .CP(wclk), .Q(ram[16141]) );
  DFF ram_reg_30__4_ ( .D(n20381), .CP(wclk), .Q(ram[16140]) );
  DFF ram_reg_30__3_ ( .D(n20380), .CP(wclk), .Q(ram[16139]) );
  DFF ram_reg_30__2_ ( .D(n20379), .CP(wclk), .Q(ram[16138]) );
  DFF ram_reg_30__1_ ( .D(n20378), .CP(wclk), .Q(ram[16137]) );
  DFF ram_reg_30__0_ ( .D(n20377), .CP(wclk), .Q(ram[16136]) );
  DFF ram_reg_34__7_ ( .D(n20352), .CP(wclk), .Q(ram[16111]) );
  DFF ram_reg_34__6_ ( .D(n20351), .CP(wclk), .Q(ram[16110]) );
  DFF ram_reg_34__5_ ( .D(n20350), .CP(wclk), .Q(ram[16109]) );
  DFF ram_reg_34__4_ ( .D(n20349), .CP(wclk), .Q(ram[16108]) );
  DFF ram_reg_34__3_ ( .D(n20348), .CP(wclk), .Q(ram[16107]) );
  DFF ram_reg_34__2_ ( .D(n20347), .CP(wclk), .Q(ram[16106]) );
  DFF ram_reg_34__1_ ( .D(n20346), .CP(wclk), .Q(ram[16105]) );
  DFF ram_reg_34__0_ ( .D(n20345), .CP(wclk), .Q(ram[16104]) );
  DFF ram_reg_38__7_ ( .D(n20320), .CP(wclk), .Q(ram[16079]) );
  DFF ram_reg_38__6_ ( .D(n20319), .CP(wclk), .Q(ram[16078]) );
  DFF ram_reg_38__5_ ( .D(n20318), .CP(wclk), .Q(ram[16077]) );
  DFF ram_reg_38__4_ ( .D(n20317), .CP(wclk), .Q(ram[16076]) );
  DFF ram_reg_38__3_ ( .D(n20316), .CP(wclk), .Q(ram[16075]) );
  DFF ram_reg_38__2_ ( .D(n20315), .CP(wclk), .Q(ram[16074]) );
  DFF ram_reg_38__1_ ( .D(n20314), .CP(wclk), .Q(ram[16073]) );
  DFF ram_reg_38__0_ ( .D(n20313), .CP(wclk), .Q(ram[16072]) );
  DFF ram_reg_42__7_ ( .D(n20288), .CP(wclk), .Q(ram[16047]) );
  DFF ram_reg_42__6_ ( .D(n20287), .CP(wclk), .Q(ram[16046]) );
  DFF ram_reg_42__5_ ( .D(n20286), .CP(wclk), .Q(ram[16045]) );
  DFF ram_reg_42__4_ ( .D(n20285), .CP(wclk), .Q(ram[16044]) );
  DFF ram_reg_42__3_ ( .D(n20284), .CP(wclk), .Q(ram[16043]) );
  DFF ram_reg_42__2_ ( .D(n20283), .CP(wclk), .Q(ram[16042]) );
  DFF ram_reg_42__1_ ( .D(n20282), .CP(wclk), .Q(ram[16041]) );
  DFF ram_reg_42__0_ ( .D(n20281), .CP(wclk), .Q(ram[16040]) );
  DFF ram_reg_46__7_ ( .D(n20256), .CP(wclk), .Q(ram[16015]) );
  DFF ram_reg_46__6_ ( .D(n20255), .CP(wclk), .Q(ram[16014]) );
  DFF ram_reg_46__5_ ( .D(n20254), .CP(wclk), .Q(ram[16013]) );
  DFF ram_reg_46__4_ ( .D(n20253), .CP(wclk), .Q(ram[16012]) );
  DFF ram_reg_46__3_ ( .D(n20252), .CP(wclk), .Q(ram[16011]) );
  DFF ram_reg_46__2_ ( .D(n20251), .CP(wclk), .Q(ram[16010]) );
  DFF ram_reg_46__1_ ( .D(n20250), .CP(wclk), .Q(ram[16009]) );
  DFF ram_reg_46__0_ ( .D(n20249), .CP(wclk), .Q(ram[16008]) );
  DFF ram_reg_50__7_ ( .D(n20224), .CP(wclk), .Q(ram[15983]) );
  DFF ram_reg_50__6_ ( .D(n20223), .CP(wclk), .Q(ram[15982]) );
  DFF ram_reg_50__5_ ( .D(n20222), .CP(wclk), .Q(ram[15981]) );
  DFF ram_reg_50__4_ ( .D(n20221), .CP(wclk), .Q(ram[15980]) );
  DFF ram_reg_50__3_ ( .D(n20220), .CP(wclk), .Q(ram[15979]) );
  DFF ram_reg_50__2_ ( .D(n20219), .CP(wclk), .Q(ram[15978]) );
  DFF ram_reg_50__1_ ( .D(n20218), .CP(wclk), .Q(ram[15977]) );
  DFF ram_reg_50__0_ ( .D(n20217), .CP(wclk), .Q(ram[15976]) );
  DFF ram_reg_54__7_ ( .D(n20192), .CP(wclk), .Q(ram[15951]) );
  DFF ram_reg_54__6_ ( .D(n20191), .CP(wclk), .Q(ram[15950]) );
  DFF ram_reg_54__5_ ( .D(n20190), .CP(wclk), .Q(ram[15949]) );
  DFF ram_reg_54__4_ ( .D(n20189), .CP(wclk), .Q(ram[15948]) );
  DFF ram_reg_54__3_ ( .D(n20188), .CP(wclk), .Q(ram[15947]) );
  DFF ram_reg_54__2_ ( .D(n20187), .CP(wclk), .Q(ram[15946]) );
  DFF ram_reg_54__1_ ( .D(n20186), .CP(wclk), .Q(ram[15945]) );
  DFF ram_reg_54__0_ ( .D(n20185), .CP(wclk), .Q(ram[15944]) );
  DFF ram_reg_58__7_ ( .D(n20160), .CP(wclk), .Q(ram[15919]) );
  DFF ram_reg_58__6_ ( .D(n20159), .CP(wclk), .Q(ram[15918]) );
  DFF ram_reg_58__5_ ( .D(n20158), .CP(wclk), .Q(ram[15917]) );
  DFF ram_reg_58__4_ ( .D(n20157), .CP(wclk), .Q(ram[15916]) );
  DFF ram_reg_58__3_ ( .D(n20156), .CP(wclk), .Q(ram[15915]) );
  DFF ram_reg_58__2_ ( .D(n20155), .CP(wclk), .Q(ram[15914]) );
  DFF ram_reg_58__1_ ( .D(n20154), .CP(wclk), .Q(ram[15913]) );
  DFF ram_reg_58__0_ ( .D(n20153), .CP(wclk), .Q(ram[15912]) );
  DFF ram_reg_62__7_ ( .D(n20128), .CP(wclk), .Q(ram[15887]) );
  DFF ram_reg_62__6_ ( .D(n20127), .CP(wclk), .Q(ram[15886]) );
  DFF ram_reg_62__5_ ( .D(n20126), .CP(wclk), .Q(ram[15885]) );
  DFF ram_reg_62__4_ ( .D(n20125), .CP(wclk), .Q(ram[15884]) );
  DFF ram_reg_62__3_ ( .D(n20124), .CP(wclk), .Q(ram[15883]) );
  DFF ram_reg_62__2_ ( .D(n20123), .CP(wclk), .Q(ram[15882]) );
  DFF ram_reg_62__1_ ( .D(n20122), .CP(wclk), .Q(ram[15881]) );
  DFF ram_reg_62__0_ ( .D(n20121), .CP(wclk), .Q(ram[15880]) );
  DFF ram_reg_66__7_ ( .D(n20096), .CP(wclk), .Q(ram[15855]) );
  DFF ram_reg_66__6_ ( .D(n20095), .CP(wclk), .Q(ram[15854]) );
  DFF ram_reg_66__5_ ( .D(n20094), .CP(wclk), .Q(ram[15853]) );
  DFF ram_reg_66__4_ ( .D(n20093), .CP(wclk), .Q(ram[15852]) );
  DFF ram_reg_66__3_ ( .D(n20092), .CP(wclk), .Q(ram[15851]) );
  DFF ram_reg_66__2_ ( .D(n20091), .CP(wclk), .Q(ram[15850]) );
  DFF ram_reg_66__1_ ( .D(n20090), .CP(wclk), .Q(ram[15849]) );
  DFF ram_reg_66__0_ ( .D(n20089), .CP(wclk), .Q(ram[15848]) );
  DFF ram_reg_70__7_ ( .D(n20064), .CP(wclk), .Q(ram[15823]) );
  DFF ram_reg_70__6_ ( .D(n20063), .CP(wclk), .Q(ram[15822]) );
  DFF ram_reg_70__5_ ( .D(n20062), .CP(wclk), .Q(ram[15821]) );
  DFF ram_reg_70__4_ ( .D(n20061), .CP(wclk), .Q(ram[15820]) );
  DFF ram_reg_70__3_ ( .D(n20060), .CP(wclk), .Q(ram[15819]) );
  DFF ram_reg_70__2_ ( .D(n20059), .CP(wclk), .Q(ram[15818]) );
  DFF ram_reg_70__1_ ( .D(n20058), .CP(wclk), .Q(ram[15817]) );
  DFF ram_reg_70__0_ ( .D(n20057), .CP(wclk), .Q(ram[15816]) );
  DFF ram_reg_74__7_ ( .D(n20032), .CP(wclk), .Q(ram[15791]) );
  DFF ram_reg_74__6_ ( .D(n20031), .CP(wclk), .Q(ram[15790]) );
  DFF ram_reg_74__5_ ( .D(n20030), .CP(wclk), .Q(ram[15789]) );
  DFF ram_reg_74__4_ ( .D(n20029), .CP(wclk), .Q(ram[15788]) );
  DFF ram_reg_74__3_ ( .D(n20028), .CP(wclk), .Q(ram[15787]) );
  DFF ram_reg_74__2_ ( .D(n20027), .CP(wclk), .Q(ram[15786]) );
  DFF ram_reg_74__1_ ( .D(n20026), .CP(wclk), .Q(ram[15785]) );
  DFF ram_reg_74__0_ ( .D(n20025), .CP(wclk), .Q(ram[15784]) );
  DFF ram_reg_78__7_ ( .D(n20000), .CP(wclk), .Q(ram[15759]) );
  DFF ram_reg_78__6_ ( .D(n19999), .CP(wclk), .Q(ram[15758]) );
  DFF ram_reg_78__5_ ( .D(n19998), .CP(wclk), .Q(ram[15757]) );
  DFF ram_reg_78__4_ ( .D(n19997), .CP(wclk), .Q(ram[15756]) );
  DFF ram_reg_78__3_ ( .D(n19996), .CP(wclk), .Q(ram[15755]) );
  DFF ram_reg_78__2_ ( .D(n19995), .CP(wclk), .Q(ram[15754]) );
  DFF ram_reg_78__1_ ( .D(n19994), .CP(wclk), .Q(ram[15753]) );
  DFF ram_reg_78__0_ ( .D(n19993), .CP(wclk), .Q(ram[15752]) );
  DFF ram_reg_82__7_ ( .D(n19968), .CP(wclk), .Q(ram[15727]) );
  DFF ram_reg_82__6_ ( .D(n19967), .CP(wclk), .Q(ram[15726]) );
  DFF ram_reg_82__5_ ( .D(n19966), .CP(wclk), .Q(ram[15725]) );
  DFF ram_reg_82__4_ ( .D(n19965), .CP(wclk), .Q(ram[15724]) );
  DFF ram_reg_82__3_ ( .D(n19964), .CP(wclk), .Q(ram[15723]) );
  DFF ram_reg_82__2_ ( .D(n19963), .CP(wclk), .Q(ram[15722]) );
  DFF ram_reg_82__1_ ( .D(n19962), .CP(wclk), .Q(ram[15721]) );
  DFF ram_reg_82__0_ ( .D(n19961), .CP(wclk), .Q(ram[15720]) );
  DFF ram_reg_86__7_ ( .D(n19936), .CP(wclk), .Q(ram[15695]) );
  DFF ram_reg_86__6_ ( .D(n19935), .CP(wclk), .Q(ram[15694]) );
  DFF ram_reg_86__5_ ( .D(n19934), .CP(wclk), .Q(ram[15693]) );
  DFF ram_reg_86__4_ ( .D(n19933), .CP(wclk), .Q(ram[15692]) );
  DFF ram_reg_86__3_ ( .D(n19932), .CP(wclk), .Q(ram[15691]) );
  DFF ram_reg_86__2_ ( .D(n19931), .CP(wclk), .Q(ram[15690]) );
  DFF ram_reg_86__1_ ( .D(n19930), .CP(wclk), .Q(ram[15689]) );
  DFF ram_reg_86__0_ ( .D(n19929), .CP(wclk), .Q(ram[15688]) );
  DFF ram_reg_90__7_ ( .D(n19904), .CP(wclk), .Q(ram[15663]) );
  DFF ram_reg_90__6_ ( .D(n19903), .CP(wclk), .Q(ram[15662]) );
  DFF ram_reg_90__5_ ( .D(n19902), .CP(wclk), .Q(ram[15661]) );
  DFF ram_reg_90__4_ ( .D(n19901), .CP(wclk), .Q(ram[15660]) );
  DFF ram_reg_90__3_ ( .D(n19900), .CP(wclk), .Q(ram[15659]) );
  DFF ram_reg_90__2_ ( .D(n19899), .CP(wclk), .Q(ram[15658]) );
  DFF ram_reg_90__1_ ( .D(n19898), .CP(wclk), .Q(ram[15657]) );
  DFF ram_reg_90__0_ ( .D(n19897), .CP(wclk), .Q(ram[15656]) );
  DFF ram_reg_94__7_ ( .D(n19872), .CP(wclk), .Q(ram[15631]) );
  DFF ram_reg_94__6_ ( .D(n19871), .CP(wclk), .Q(ram[15630]) );
  DFF ram_reg_94__5_ ( .D(n19870), .CP(wclk), .Q(ram[15629]) );
  DFF ram_reg_94__4_ ( .D(n19869), .CP(wclk), .Q(ram[15628]) );
  DFF ram_reg_94__3_ ( .D(n19868), .CP(wclk), .Q(ram[15627]) );
  DFF ram_reg_94__2_ ( .D(n19867), .CP(wclk), .Q(ram[15626]) );
  DFF ram_reg_94__1_ ( .D(n19866), .CP(wclk), .Q(ram[15625]) );
  DFF ram_reg_94__0_ ( .D(n19865), .CP(wclk), .Q(ram[15624]) );
  DFF ram_reg_98__7_ ( .D(n19840), .CP(wclk), .Q(ram[15599]) );
  DFF ram_reg_98__6_ ( .D(n19839), .CP(wclk), .Q(ram[15598]) );
  DFF ram_reg_98__5_ ( .D(n19838), .CP(wclk), .Q(ram[15597]) );
  DFF ram_reg_98__4_ ( .D(n19837), .CP(wclk), .Q(ram[15596]) );
  DFF ram_reg_98__3_ ( .D(n19836), .CP(wclk), .Q(ram[15595]) );
  DFF ram_reg_98__2_ ( .D(n19835), .CP(wclk), .Q(ram[15594]) );
  DFF ram_reg_98__1_ ( .D(n19834), .CP(wclk), .Q(ram[15593]) );
  DFF ram_reg_98__0_ ( .D(n19833), .CP(wclk), .Q(ram[15592]) );
  DFF ram_reg_102__7_ ( .D(n19808), .CP(wclk), .Q(ram[15567]) );
  DFF ram_reg_102__6_ ( .D(n19807), .CP(wclk), .Q(ram[15566]) );
  DFF ram_reg_102__5_ ( .D(n19806), .CP(wclk), .Q(ram[15565]) );
  DFF ram_reg_102__4_ ( .D(n19805), .CP(wclk), .Q(ram[15564]) );
  DFF ram_reg_102__3_ ( .D(n19804), .CP(wclk), .Q(ram[15563]) );
  DFF ram_reg_102__2_ ( .D(n19803), .CP(wclk), .Q(ram[15562]) );
  DFF ram_reg_102__1_ ( .D(n19802), .CP(wclk), .Q(ram[15561]) );
  DFF ram_reg_102__0_ ( .D(n19801), .CP(wclk), .Q(ram[15560]) );
  DFF ram_reg_106__7_ ( .D(n19776), .CP(wclk), .Q(ram[15535]) );
  DFF ram_reg_106__6_ ( .D(n19775), .CP(wclk), .Q(ram[15534]) );
  DFF ram_reg_106__5_ ( .D(n19774), .CP(wclk), .Q(ram[15533]) );
  DFF ram_reg_106__4_ ( .D(n19773), .CP(wclk), .Q(ram[15532]) );
  DFF ram_reg_106__3_ ( .D(n19772), .CP(wclk), .Q(ram[15531]) );
  DFF ram_reg_106__2_ ( .D(n19771), .CP(wclk), .Q(ram[15530]) );
  DFF ram_reg_106__1_ ( .D(n19770), .CP(wclk), .Q(ram[15529]) );
  DFF ram_reg_106__0_ ( .D(n19769), .CP(wclk), .Q(ram[15528]) );
  DFF ram_reg_110__7_ ( .D(n19744), .CP(wclk), .Q(ram[15503]) );
  DFF ram_reg_110__6_ ( .D(n19743), .CP(wclk), .Q(ram[15502]) );
  DFF ram_reg_110__5_ ( .D(n19742), .CP(wclk), .Q(ram[15501]) );
  DFF ram_reg_110__4_ ( .D(n19741), .CP(wclk), .Q(ram[15500]) );
  DFF ram_reg_110__3_ ( .D(n19740), .CP(wclk), .Q(ram[15499]) );
  DFF ram_reg_110__2_ ( .D(n19739), .CP(wclk), .Q(ram[15498]) );
  DFF ram_reg_110__1_ ( .D(n19738), .CP(wclk), .Q(ram[15497]) );
  DFF ram_reg_110__0_ ( .D(n19737), .CP(wclk), .Q(ram[15496]) );
  DFF ram_reg_114__7_ ( .D(n19712), .CP(wclk), .Q(ram[15471]) );
  DFF ram_reg_114__6_ ( .D(n19711), .CP(wclk), .Q(ram[15470]) );
  DFF ram_reg_114__5_ ( .D(n19710), .CP(wclk), .Q(ram[15469]) );
  DFF ram_reg_114__4_ ( .D(n19709), .CP(wclk), .Q(ram[15468]) );
  DFF ram_reg_114__3_ ( .D(n19708), .CP(wclk), .Q(ram[15467]) );
  DFF ram_reg_114__2_ ( .D(n19707), .CP(wclk), .Q(ram[15466]) );
  DFF ram_reg_114__1_ ( .D(n19706), .CP(wclk), .Q(ram[15465]) );
  DFF ram_reg_114__0_ ( .D(n19705), .CP(wclk), .Q(ram[15464]) );
  DFF ram_reg_118__7_ ( .D(n19680), .CP(wclk), .Q(ram[15439]) );
  DFF ram_reg_118__6_ ( .D(n19679), .CP(wclk), .Q(ram[15438]) );
  DFF ram_reg_118__5_ ( .D(n19678), .CP(wclk), .Q(ram[15437]) );
  DFF ram_reg_118__4_ ( .D(n19677), .CP(wclk), .Q(ram[15436]) );
  DFF ram_reg_118__3_ ( .D(n19676), .CP(wclk), .Q(ram[15435]) );
  DFF ram_reg_118__2_ ( .D(n19675), .CP(wclk), .Q(ram[15434]) );
  DFF ram_reg_118__1_ ( .D(n19674), .CP(wclk), .Q(ram[15433]) );
  DFF ram_reg_118__0_ ( .D(n19673), .CP(wclk), .Q(ram[15432]) );
  DFF ram_reg_122__7_ ( .D(n19648), .CP(wclk), .Q(ram[15407]) );
  DFF ram_reg_122__6_ ( .D(n19647), .CP(wclk), .Q(ram[15406]) );
  DFF ram_reg_122__5_ ( .D(n19646), .CP(wclk), .Q(ram[15405]) );
  DFF ram_reg_122__4_ ( .D(n19645), .CP(wclk), .Q(ram[15404]) );
  DFF ram_reg_122__3_ ( .D(n19644), .CP(wclk), .Q(ram[15403]) );
  DFF ram_reg_122__2_ ( .D(n19643), .CP(wclk), .Q(ram[15402]) );
  DFF ram_reg_122__1_ ( .D(n19642), .CP(wclk), .Q(ram[15401]) );
  DFF ram_reg_122__0_ ( .D(n19641), .CP(wclk), .Q(ram[15400]) );
  DFF ram_reg_126__7_ ( .D(n19616), .CP(wclk), .Q(ram[15375]) );
  DFF ram_reg_126__6_ ( .D(n19615), .CP(wclk), .Q(ram[15374]) );
  DFF ram_reg_126__5_ ( .D(n19614), .CP(wclk), .Q(ram[15373]) );
  DFF ram_reg_126__4_ ( .D(n19613), .CP(wclk), .Q(ram[15372]) );
  DFF ram_reg_126__3_ ( .D(n19612), .CP(wclk), .Q(ram[15371]) );
  DFF ram_reg_126__2_ ( .D(n19611), .CP(wclk), .Q(ram[15370]) );
  DFF ram_reg_126__1_ ( .D(n19610), .CP(wclk), .Q(ram[15369]) );
  DFF ram_reg_126__0_ ( .D(n19609), .CP(wclk), .Q(ram[15368]) );
  DFF ram_reg_130__7_ ( .D(n19584), .CP(wclk), .Q(ram[15343]) );
  DFF ram_reg_130__6_ ( .D(n19583), .CP(wclk), .Q(ram[15342]) );
  DFF ram_reg_130__5_ ( .D(n19582), .CP(wclk), .Q(ram[15341]) );
  DFF ram_reg_130__4_ ( .D(n19581), .CP(wclk), .Q(ram[15340]) );
  DFF ram_reg_130__3_ ( .D(n19580), .CP(wclk), .Q(ram[15339]) );
  DFF ram_reg_130__2_ ( .D(n19579), .CP(wclk), .Q(ram[15338]) );
  DFF ram_reg_130__1_ ( .D(n19578), .CP(wclk), .Q(ram[15337]) );
  DFF ram_reg_130__0_ ( .D(n19577), .CP(wclk), .Q(ram[15336]) );
  DFF ram_reg_134__7_ ( .D(n19552), .CP(wclk), .Q(ram[15311]) );
  DFF ram_reg_134__6_ ( .D(n19551), .CP(wclk), .Q(ram[15310]) );
  DFF ram_reg_134__5_ ( .D(n19550), .CP(wclk), .Q(ram[15309]) );
  DFF ram_reg_134__4_ ( .D(n19549), .CP(wclk), .Q(ram[15308]) );
  DFF ram_reg_134__3_ ( .D(n19548), .CP(wclk), .Q(ram[15307]) );
  DFF ram_reg_134__2_ ( .D(n19547), .CP(wclk), .Q(ram[15306]) );
  DFF ram_reg_134__1_ ( .D(n19546), .CP(wclk), .Q(ram[15305]) );
  DFF ram_reg_134__0_ ( .D(n19545), .CP(wclk), .Q(ram[15304]) );
  DFF ram_reg_142__7_ ( .D(n19488), .CP(wclk), .Q(ram[15247]) );
  DFF ram_reg_142__6_ ( .D(n19487), .CP(wclk), .Q(ram[15246]) );
  DFF ram_reg_142__5_ ( .D(n19486), .CP(wclk), .Q(ram[15245]) );
  DFF ram_reg_142__4_ ( .D(n19485), .CP(wclk), .Q(ram[15244]) );
  DFF ram_reg_142__3_ ( .D(n19484), .CP(wclk), .Q(ram[15243]) );
  DFF ram_reg_142__2_ ( .D(n19483), .CP(wclk), .Q(ram[15242]) );
  DFF ram_reg_142__1_ ( .D(n19482), .CP(wclk), .Q(ram[15241]) );
  DFF ram_reg_142__0_ ( .D(n19481), .CP(wclk), .Q(ram[15240]) );
  DFF ram_reg_146__7_ ( .D(n19456), .CP(wclk), .Q(ram[15215]) );
  DFF ram_reg_146__6_ ( .D(n19455), .CP(wclk), .Q(ram[15214]) );
  DFF ram_reg_146__5_ ( .D(n19454), .CP(wclk), .Q(ram[15213]) );
  DFF ram_reg_146__4_ ( .D(n19453), .CP(wclk), .Q(ram[15212]) );
  DFF ram_reg_146__3_ ( .D(n19452), .CP(wclk), .Q(ram[15211]) );
  DFF ram_reg_146__2_ ( .D(n19451), .CP(wclk), .Q(ram[15210]) );
  DFF ram_reg_146__1_ ( .D(n19450), .CP(wclk), .Q(ram[15209]) );
  DFF ram_reg_146__0_ ( .D(n19449), .CP(wclk), .Q(ram[15208]) );
  DFF ram_reg_150__7_ ( .D(n19424), .CP(wclk), .Q(ram[15183]) );
  DFF ram_reg_150__6_ ( .D(n19423), .CP(wclk), .Q(ram[15182]) );
  DFF ram_reg_150__5_ ( .D(n19422), .CP(wclk), .Q(ram[15181]) );
  DFF ram_reg_150__4_ ( .D(n19421), .CP(wclk), .Q(ram[15180]) );
  DFF ram_reg_150__3_ ( .D(n19420), .CP(wclk), .Q(ram[15179]) );
  DFF ram_reg_150__2_ ( .D(n19419), .CP(wclk), .Q(ram[15178]) );
  DFF ram_reg_150__1_ ( .D(n19418), .CP(wclk), .Q(ram[15177]) );
  DFF ram_reg_150__0_ ( .D(n19417), .CP(wclk), .Q(ram[15176]) );
  DFF ram_reg_154__7_ ( .D(n19392), .CP(wclk), .Q(ram[15151]) );
  DFF ram_reg_154__6_ ( .D(n19391), .CP(wclk), .Q(ram[15150]) );
  DFF ram_reg_154__5_ ( .D(n19390), .CP(wclk), .Q(ram[15149]) );
  DFF ram_reg_154__4_ ( .D(n19389), .CP(wclk), .Q(ram[15148]) );
  DFF ram_reg_154__3_ ( .D(n19388), .CP(wclk), .Q(ram[15147]) );
  DFF ram_reg_154__2_ ( .D(n19387), .CP(wclk), .Q(ram[15146]) );
  DFF ram_reg_154__1_ ( .D(n19386), .CP(wclk), .Q(ram[15145]) );
  DFF ram_reg_154__0_ ( .D(n19385), .CP(wclk), .Q(ram[15144]) );
  DFF ram_reg_158__7_ ( .D(n19360), .CP(wclk), .Q(ram[15119]) );
  DFF ram_reg_158__6_ ( .D(n19359), .CP(wclk), .Q(ram[15118]) );
  DFF ram_reg_158__5_ ( .D(n19358), .CP(wclk), .Q(ram[15117]) );
  DFF ram_reg_158__4_ ( .D(n19357), .CP(wclk), .Q(ram[15116]) );
  DFF ram_reg_158__3_ ( .D(n19356), .CP(wclk), .Q(ram[15115]) );
  DFF ram_reg_158__2_ ( .D(n19355), .CP(wclk), .Q(ram[15114]) );
  DFF ram_reg_158__1_ ( .D(n19354), .CP(wclk), .Q(ram[15113]) );
  DFF ram_reg_158__0_ ( .D(n19353), .CP(wclk), .Q(ram[15112]) );
  DFF ram_reg_162__7_ ( .D(n19328), .CP(wclk), .Q(ram[15087]) );
  DFF ram_reg_162__6_ ( .D(n19327), .CP(wclk), .Q(ram[15086]) );
  DFF ram_reg_162__5_ ( .D(n19326), .CP(wclk), .Q(ram[15085]) );
  DFF ram_reg_162__4_ ( .D(n19325), .CP(wclk), .Q(ram[15084]) );
  DFF ram_reg_162__3_ ( .D(n19324), .CP(wclk), .Q(ram[15083]) );
  DFF ram_reg_162__2_ ( .D(n19323), .CP(wclk), .Q(ram[15082]) );
  DFF ram_reg_162__1_ ( .D(n19322), .CP(wclk), .Q(ram[15081]) );
  DFF ram_reg_162__0_ ( .D(n19321), .CP(wclk), .Q(ram[15080]) );
  DFF ram_reg_166__7_ ( .D(n19296), .CP(wclk), .Q(ram[15055]) );
  DFF ram_reg_166__6_ ( .D(n19295), .CP(wclk), .Q(ram[15054]) );
  DFF ram_reg_166__5_ ( .D(n19294), .CP(wclk), .Q(ram[15053]) );
  DFF ram_reg_166__4_ ( .D(n19293), .CP(wclk), .Q(ram[15052]) );
  DFF ram_reg_166__3_ ( .D(n19292), .CP(wclk), .Q(ram[15051]) );
  DFF ram_reg_166__2_ ( .D(n19291), .CP(wclk), .Q(ram[15050]) );
  DFF ram_reg_166__1_ ( .D(n19290), .CP(wclk), .Q(ram[15049]) );
  DFF ram_reg_166__0_ ( .D(n19289), .CP(wclk), .Q(ram[15048]) );
  DFF ram_reg_178__7_ ( .D(n19200), .CP(wclk), .Q(ram[14959]) );
  DFF ram_reg_178__6_ ( .D(n19199), .CP(wclk), .Q(ram[14958]) );
  DFF ram_reg_178__5_ ( .D(n19198), .CP(wclk), .Q(ram[14957]) );
  DFF ram_reg_178__4_ ( .D(n19197), .CP(wclk), .Q(ram[14956]) );
  DFF ram_reg_178__3_ ( .D(n19196), .CP(wclk), .Q(ram[14955]) );
  DFF ram_reg_178__2_ ( .D(n19195), .CP(wclk), .Q(ram[14954]) );
  DFF ram_reg_178__1_ ( .D(n19194), .CP(wclk), .Q(ram[14953]) );
  DFF ram_reg_178__0_ ( .D(n19193), .CP(wclk), .Q(ram[14952]) );
  DFF ram_reg_182__7_ ( .D(n19168), .CP(wclk), .Q(ram[14927]) );
  DFF ram_reg_182__6_ ( .D(n19167), .CP(wclk), .Q(ram[14926]) );
  DFF ram_reg_182__5_ ( .D(n19166), .CP(wclk), .Q(ram[14925]) );
  DFF ram_reg_182__4_ ( .D(n19165), .CP(wclk), .Q(ram[14924]) );
  DFF ram_reg_182__3_ ( .D(n19164), .CP(wclk), .Q(ram[14923]) );
  DFF ram_reg_182__2_ ( .D(n19163), .CP(wclk), .Q(ram[14922]) );
  DFF ram_reg_182__1_ ( .D(n19162), .CP(wclk), .Q(ram[14921]) );
  DFF ram_reg_182__0_ ( .D(n19161), .CP(wclk), .Q(ram[14920]) );
  DFF ram_reg_194__7_ ( .D(n19072), .CP(wclk), .Q(ram[14831]) );
  DFF ram_reg_194__6_ ( .D(n19071), .CP(wclk), .Q(ram[14830]) );
  DFF ram_reg_194__5_ ( .D(n19070), .CP(wclk), .Q(ram[14829]) );
  DFF ram_reg_194__4_ ( .D(n19069), .CP(wclk), .Q(ram[14828]) );
  DFF ram_reg_194__3_ ( .D(n19068), .CP(wclk), .Q(ram[14827]) );
  DFF ram_reg_194__2_ ( .D(n19067), .CP(wclk), .Q(ram[14826]) );
  DFF ram_reg_194__1_ ( .D(n19066), .CP(wclk), .Q(ram[14825]) );
  DFF ram_reg_194__0_ ( .D(n19065), .CP(wclk), .Q(ram[14824]) );
  DFF ram_reg_198__7_ ( .D(n19040), .CP(wclk), .Q(ram[14799]) );
  DFF ram_reg_198__6_ ( .D(n19039), .CP(wclk), .Q(ram[14798]) );
  DFF ram_reg_198__5_ ( .D(n19038), .CP(wclk), .Q(ram[14797]) );
  DFF ram_reg_198__4_ ( .D(n19037), .CP(wclk), .Q(ram[14796]) );
  DFF ram_reg_198__3_ ( .D(n19036), .CP(wclk), .Q(ram[14795]) );
  DFF ram_reg_198__2_ ( .D(n19035), .CP(wclk), .Q(ram[14794]) );
  DFF ram_reg_198__1_ ( .D(n19034), .CP(wclk), .Q(ram[14793]) );
  DFF ram_reg_198__0_ ( .D(n19033), .CP(wclk), .Q(ram[14792]) );
  DFF ram_reg_202__7_ ( .D(n19008), .CP(wclk), .Q(ram[14767]) );
  DFF ram_reg_202__6_ ( .D(n19007), .CP(wclk), .Q(ram[14766]) );
  DFF ram_reg_202__5_ ( .D(n19006), .CP(wclk), .Q(ram[14765]) );
  DFF ram_reg_202__4_ ( .D(n19005), .CP(wclk), .Q(ram[14764]) );
  DFF ram_reg_202__3_ ( .D(n19004), .CP(wclk), .Q(ram[14763]) );
  DFF ram_reg_202__2_ ( .D(n19003), .CP(wclk), .Q(ram[14762]) );
  DFF ram_reg_202__1_ ( .D(n19002), .CP(wclk), .Q(ram[14761]) );
  DFF ram_reg_202__0_ ( .D(n19001), .CP(wclk), .Q(ram[14760]) );
  DFF ram_reg_206__7_ ( .D(n18976), .CP(wclk), .Q(ram[14735]) );
  DFF ram_reg_206__6_ ( .D(n18975), .CP(wclk), .Q(ram[14734]) );
  DFF ram_reg_206__5_ ( .D(n18974), .CP(wclk), .Q(ram[14733]) );
  DFF ram_reg_206__4_ ( .D(n18973), .CP(wclk), .Q(ram[14732]) );
  DFF ram_reg_206__3_ ( .D(n18972), .CP(wclk), .Q(ram[14731]) );
  DFF ram_reg_206__2_ ( .D(n18971), .CP(wclk), .Q(ram[14730]) );
  DFF ram_reg_206__1_ ( .D(n18970), .CP(wclk), .Q(ram[14729]) );
  DFF ram_reg_206__0_ ( .D(n18969), .CP(wclk), .Q(ram[14728]) );
  DFF ram_reg_210__7_ ( .D(n18944), .CP(wclk), .Q(ram[14703]) );
  DFF ram_reg_210__6_ ( .D(n18943), .CP(wclk), .Q(ram[14702]) );
  DFF ram_reg_210__5_ ( .D(n18942), .CP(wclk), .Q(ram[14701]) );
  DFF ram_reg_210__4_ ( .D(n18941), .CP(wclk), .Q(ram[14700]) );
  DFF ram_reg_210__3_ ( .D(n18940), .CP(wclk), .Q(ram[14699]) );
  DFF ram_reg_210__2_ ( .D(n18939), .CP(wclk), .Q(ram[14698]) );
  DFF ram_reg_210__1_ ( .D(n18938), .CP(wclk), .Q(ram[14697]) );
  DFF ram_reg_210__0_ ( .D(n18937), .CP(wclk), .Q(ram[14696]) );
  DFF ram_reg_214__7_ ( .D(n18912), .CP(wclk), .Q(ram[14671]) );
  DFF ram_reg_214__6_ ( .D(n18911), .CP(wclk), .Q(ram[14670]) );
  DFF ram_reg_214__5_ ( .D(n18910), .CP(wclk), .Q(ram[14669]) );
  DFF ram_reg_214__4_ ( .D(n18909), .CP(wclk), .Q(ram[14668]) );
  DFF ram_reg_214__3_ ( .D(n18908), .CP(wclk), .Q(ram[14667]) );
  DFF ram_reg_214__2_ ( .D(n18907), .CP(wclk), .Q(ram[14666]) );
  DFF ram_reg_214__1_ ( .D(n18906), .CP(wclk), .Q(ram[14665]) );
  DFF ram_reg_214__0_ ( .D(n18905), .CP(wclk), .Q(ram[14664]) );
  DFF ram_reg_218__7_ ( .D(n18880), .CP(wclk), .Q(ram[14639]) );
  DFF ram_reg_218__6_ ( .D(n18879), .CP(wclk), .Q(ram[14638]) );
  DFF ram_reg_218__5_ ( .D(n18878), .CP(wclk), .Q(ram[14637]) );
  DFF ram_reg_218__4_ ( .D(n18877), .CP(wclk), .Q(ram[14636]) );
  DFF ram_reg_218__3_ ( .D(n18876), .CP(wclk), .Q(ram[14635]) );
  DFF ram_reg_218__2_ ( .D(n18875), .CP(wclk), .Q(ram[14634]) );
  DFF ram_reg_218__1_ ( .D(n18874), .CP(wclk), .Q(ram[14633]) );
  DFF ram_reg_218__0_ ( .D(n18873), .CP(wclk), .Q(ram[14632]) );
  DFF ram_reg_222__7_ ( .D(n18848), .CP(wclk), .Q(ram[14607]) );
  DFF ram_reg_222__6_ ( .D(n18847), .CP(wclk), .Q(ram[14606]) );
  DFF ram_reg_222__5_ ( .D(n18846), .CP(wclk), .Q(ram[14605]) );
  DFF ram_reg_222__4_ ( .D(n18845), .CP(wclk), .Q(ram[14604]) );
  DFF ram_reg_222__3_ ( .D(n18844), .CP(wclk), .Q(ram[14603]) );
  DFF ram_reg_222__2_ ( .D(n18843), .CP(wclk), .Q(ram[14602]) );
  DFF ram_reg_222__1_ ( .D(n18842), .CP(wclk), .Q(ram[14601]) );
  DFF ram_reg_222__0_ ( .D(n18841), .CP(wclk), .Q(ram[14600]) );
  DFF ram_reg_226__7_ ( .D(n18816), .CP(wclk), .Q(ram[14575]) );
  DFF ram_reg_226__6_ ( .D(n18815), .CP(wclk), .Q(ram[14574]) );
  DFF ram_reg_226__5_ ( .D(n18814), .CP(wclk), .Q(ram[14573]) );
  DFF ram_reg_226__4_ ( .D(n18813), .CP(wclk), .Q(ram[14572]) );
  DFF ram_reg_226__3_ ( .D(n18812), .CP(wclk), .Q(ram[14571]) );
  DFF ram_reg_226__2_ ( .D(n18811), .CP(wclk), .Q(ram[14570]) );
  DFF ram_reg_226__1_ ( .D(n18810), .CP(wclk), .Q(ram[14569]) );
  DFF ram_reg_226__0_ ( .D(n18809), .CP(wclk), .Q(ram[14568]) );
  DFF ram_reg_230__7_ ( .D(n18784), .CP(wclk), .Q(ram[14543]) );
  DFF ram_reg_230__6_ ( .D(n18783), .CP(wclk), .Q(ram[14542]) );
  DFF ram_reg_230__5_ ( .D(n18782), .CP(wclk), .Q(ram[14541]) );
  DFF ram_reg_230__4_ ( .D(n18781), .CP(wclk), .Q(ram[14540]) );
  DFF ram_reg_230__3_ ( .D(n18780), .CP(wclk), .Q(ram[14539]) );
  DFF ram_reg_230__2_ ( .D(n18779), .CP(wclk), .Q(ram[14538]) );
  DFF ram_reg_230__1_ ( .D(n18778), .CP(wclk), .Q(ram[14537]) );
  DFF ram_reg_230__0_ ( .D(n18777), .CP(wclk), .Q(ram[14536]) );
  DFF ram_reg_238__7_ ( .D(n18720), .CP(wclk), .Q(ram[14479]) );
  DFF ram_reg_238__6_ ( .D(n18719), .CP(wclk), .Q(ram[14478]) );
  DFF ram_reg_238__5_ ( .D(n18718), .CP(wclk), .Q(ram[14477]) );
  DFF ram_reg_238__4_ ( .D(n18717), .CP(wclk), .Q(ram[14476]) );
  DFF ram_reg_238__3_ ( .D(n18716), .CP(wclk), .Q(ram[14475]) );
  DFF ram_reg_238__2_ ( .D(n18715), .CP(wclk), .Q(ram[14474]) );
  DFF ram_reg_238__1_ ( .D(n18714), .CP(wclk), .Q(ram[14473]) );
  DFF ram_reg_238__0_ ( .D(n18713), .CP(wclk), .Q(ram[14472]) );
  DFF ram_reg_242__7_ ( .D(n18688), .CP(wclk), .Q(ram[14447]) );
  DFF ram_reg_242__6_ ( .D(n18687), .CP(wclk), .Q(ram[14446]) );
  DFF ram_reg_242__5_ ( .D(n18686), .CP(wclk), .Q(ram[14445]) );
  DFF ram_reg_242__4_ ( .D(n18685), .CP(wclk), .Q(ram[14444]) );
  DFF ram_reg_242__3_ ( .D(n18684), .CP(wclk), .Q(ram[14443]) );
  DFF ram_reg_242__2_ ( .D(n18683), .CP(wclk), .Q(ram[14442]) );
  DFF ram_reg_242__1_ ( .D(n18682), .CP(wclk), .Q(ram[14441]) );
  DFF ram_reg_242__0_ ( .D(n18681), .CP(wclk), .Q(ram[14440]) );
  DFF ram_reg_246__7_ ( .D(n18656), .CP(wclk), .Q(ram[14415]) );
  DFF ram_reg_246__6_ ( .D(n18655), .CP(wclk), .Q(ram[14414]) );
  DFF ram_reg_246__5_ ( .D(n18654), .CP(wclk), .Q(ram[14413]) );
  DFF ram_reg_246__4_ ( .D(n18653), .CP(wclk), .Q(ram[14412]) );
  DFF ram_reg_246__3_ ( .D(n18652), .CP(wclk), .Q(ram[14411]) );
  DFF ram_reg_246__2_ ( .D(n18651), .CP(wclk), .Q(ram[14410]) );
  DFF ram_reg_246__1_ ( .D(n18650), .CP(wclk), .Q(ram[14409]) );
  DFF ram_reg_246__0_ ( .D(n18649), .CP(wclk), .Q(ram[14408]) );
  DFF ram_reg_258__7_ ( .D(n18560), .CP(wclk), .Q(ram[14319]) );
  DFF ram_reg_258__6_ ( .D(n18559), .CP(wclk), .Q(ram[14318]) );
  DFF ram_reg_258__5_ ( .D(n18558), .CP(wclk), .Q(ram[14317]) );
  DFF ram_reg_258__4_ ( .D(n18557), .CP(wclk), .Q(ram[14316]) );
  DFF ram_reg_258__3_ ( .D(n18556), .CP(wclk), .Q(ram[14315]) );
  DFF ram_reg_258__2_ ( .D(n18555), .CP(wclk), .Q(ram[14314]) );
  DFF ram_reg_258__1_ ( .D(n18554), .CP(wclk), .Q(ram[14313]) );
  DFF ram_reg_258__0_ ( .D(n18553), .CP(wclk), .Q(ram[14312]) );
  DFF ram_reg_262__7_ ( .D(n18528), .CP(wclk), .Q(ram[14287]) );
  DFF ram_reg_262__6_ ( .D(n18527), .CP(wclk), .Q(ram[14286]) );
  DFF ram_reg_262__5_ ( .D(n18526), .CP(wclk), .Q(ram[14285]) );
  DFF ram_reg_262__4_ ( .D(n18525), .CP(wclk), .Q(ram[14284]) );
  DFF ram_reg_262__3_ ( .D(n18524), .CP(wclk), .Q(ram[14283]) );
  DFF ram_reg_262__2_ ( .D(n18523), .CP(wclk), .Q(ram[14282]) );
  DFF ram_reg_262__1_ ( .D(n18522), .CP(wclk), .Q(ram[14281]) );
  DFF ram_reg_262__0_ ( .D(n18521), .CP(wclk), .Q(ram[14280]) );
  DFF ram_reg_266__7_ ( .D(n18496), .CP(wclk), .Q(ram[14255]) );
  DFF ram_reg_266__6_ ( .D(n18495), .CP(wclk), .Q(ram[14254]) );
  DFF ram_reg_266__5_ ( .D(n18494), .CP(wclk), .Q(ram[14253]) );
  DFF ram_reg_266__4_ ( .D(n18493), .CP(wclk), .Q(ram[14252]) );
  DFF ram_reg_266__3_ ( .D(n18492), .CP(wclk), .Q(ram[14251]) );
  DFF ram_reg_266__2_ ( .D(n18491), .CP(wclk), .Q(ram[14250]) );
  DFF ram_reg_266__1_ ( .D(n18490), .CP(wclk), .Q(ram[14249]) );
  DFF ram_reg_266__0_ ( .D(n18489), .CP(wclk), .Q(ram[14248]) );
  DFF ram_reg_270__7_ ( .D(n18464), .CP(wclk), .Q(ram[14223]) );
  DFF ram_reg_270__6_ ( .D(n18463), .CP(wclk), .Q(ram[14222]) );
  DFF ram_reg_270__5_ ( .D(n18462), .CP(wclk), .Q(ram[14221]) );
  DFF ram_reg_270__4_ ( .D(n18461), .CP(wclk), .Q(ram[14220]) );
  DFF ram_reg_270__3_ ( .D(n18460), .CP(wclk), .Q(ram[14219]) );
  DFF ram_reg_270__2_ ( .D(n18459), .CP(wclk), .Q(ram[14218]) );
  DFF ram_reg_270__1_ ( .D(n18458), .CP(wclk), .Q(ram[14217]) );
  DFF ram_reg_270__0_ ( .D(n18457), .CP(wclk), .Q(ram[14216]) );
  DFF ram_reg_274__7_ ( .D(n18432), .CP(wclk), .Q(ram[14191]) );
  DFF ram_reg_274__6_ ( .D(n18431), .CP(wclk), .Q(ram[14190]) );
  DFF ram_reg_274__5_ ( .D(n18430), .CP(wclk), .Q(ram[14189]) );
  DFF ram_reg_274__4_ ( .D(n18429), .CP(wclk), .Q(ram[14188]) );
  DFF ram_reg_274__3_ ( .D(n18428), .CP(wclk), .Q(ram[14187]) );
  DFF ram_reg_274__2_ ( .D(n18427), .CP(wclk), .Q(ram[14186]) );
  DFF ram_reg_274__1_ ( .D(n18426), .CP(wclk), .Q(ram[14185]) );
  DFF ram_reg_274__0_ ( .D(n18425), .CP(wclk), .Q(ram[14184]) );
  DFF ram_reg_278__7_ ( .D(n18400), .CP(wclk), .Q(ram[14159]) );
  DFF ram_reg_278__6_ ( .D(n18399), .CP(wclk), .Q(ram[14158]) );
  DFF ram_reg_278__5_ ( .D(n18398), .CP(wclk), .Q(ram[14157]) );
  DFF ram_reg_278__4_ ( .D(n18397), .CP(wclk), .Q(ram[14156]) );
  DFF ram_reg_278__3_ ( .D(n18396), .CP(wclk), .Q(ram[14155]) );
  DFF ram_reg_278__2_ ( .D(n18395), .CP(wclk), .Q(ram[14154]) );
  DFF ram_reg_278__1_ ( .D(n18394), .CP(wclk), .Q(ram[14153]) );
  DFF ram_reg_278__0_ ( .D(n18393), .CP(wclk), .Q(ram[14152]) );
  DFF ram_reg_282__7_ ( .D(n18368), .CP(wclk), .Q(ram[14127]) );
  DFF ram_reg_282__6_ ( .D(n18367), .CP(wclk), .Q(ram[14126]) );
  DFF ram_reg_282__5_ ( .D(n18366), .CP(wclk), .Q(ram[14125]) );
  DFF ram_reg_282__4_ ( .D(n18365), .CP(wclk), .Q(ram[14124]) );
  DFF ram_reg_282__3_ ( .D(n18364), .CP(wclk), .Q(ram[14123]) );
  DFF ram_reg_282__2_ ( .D(n18363), .CP(wclk), .Q(ram[14122]) );
  DFF ram_reg_282__1_ ( .D(n18362), .CP(wclk), .Q(ram[14121]) );
  DFF ram_reg_282__0_ ( .D(n18361), .CP(wclk), .Q(ram[14120]) );
  DFF ram_reg_286__7_ ( .D(n18336), .CP(wclk), .Q(ram[14095]) );
  DFF ram_reg_286__6_ ( .D(n18335), .CP(wclk), .Q(ram[14094]) );
  DFF ram_reg_286__5_ ( .D(n18334), .CP(wclk), .Q(ram[14093]) );
  DFF ram_reg_286__4_ ( .D(n18333), .CP(wclk), .Q(ram[14092]) );
  DFF ram_reg_286__3_ ( .D(n18332), .CP(wclk), .Q(ram[14091]) );
  DFF ram_reg_286__2_ ( .D(n18331), .CP(wclk), .Q(ram[14090]) );
  DFF ram_reg_286__1_ ( .D(n18330), .CP(wclk), .Q(ram[14089]) );
  DFF ram_reg_286__0_ ( .D(n18329), .CP(wclk), .Q(ram[14088]) );
  DFF ram_reg_290__7_ ( .D(n18304), .CP(wclk), .Q(ram[14063]) );
  DFF ram_reg_290__6_ ( .D(n18303), .CP(wclk), .Q(ram[14062]) );
  DFF ram_reg_290__5_ ( .D(n18302), .CP(wclk), .Q(ram[14061]) );
  DFF ram_reg_290__4_ ( .D(n18301), .CP(wclk), .Q(ram[14060]) );
  DFF ram_reg_290__3_ ( .D(n18300), .CP(wclk), .Q(ram[14059]) );
  DFF ram_reg_290__2_ ( .D(n18299), .CP(wclk), .Q(ram[14058]) );
  DFF ram_reg_290__1_ ( .D(n18298), .CP(wclk), .Q(ram[14057]) );
  DFF ram_reg_290__0_ ( .D(n18297), .CP(wclk), .Q(ram[14056]) );
  DFF ram_reg_294__7_ ( .D(n18272), .CP(wclk), .Q(ram[14031]) );
  DFF ram_reg_294__6_ ( .D(n18271), .CP(wclk), .Q(ram[14030]) );
  DFF ram_reg_294__5_ ( .D(n18270), .CP(wclk), .Q(ram[14029]) );
  DFF ram_reg_294__4_ ( .D(n18269), .CP(wclk), .Q(ram[14028]) );
  DFF ram_reg_294__3_ ( .D(n18268), .CP(wclk), .Q(ram[14027]) );
  DFF ram_reg_294__2_ ( .D(n18267), .CP(wclk), .Q(ram[14026]) );
  DFF ram_reg_294__1_ ( .D(n18266), .CP(wclk), .Q(ram[14025]) );
  DFF ram_reg_294__0_ ( .D(n18265), .CP(wclk), .Q(ram[14024]) );
  DFF ram_reg_298__7_ ( .D(n18240), .CP(wclk), .Q(ram[13999]) );
  DFF ram_reg_298__6_ ( .D(n18239), .CP(wclk), .Q(ram[13998]) );
  DFF ram_reg_298__5_ ( .D(n18238), .CP(wclk), .Q(ram[13997]) );
  DFF ram_reg_298__4_ ( .D(n18237), .CP(wclk), .Q(ram[13996]) );
  DFF ram_reg_298__3_ ( .D(n18236), .CP(wclk), .Q(ram[13995]) );
  DFF ram_reg_298__2_ ( .D(n18235), .CP(wclk), .Q(ram[13994]) );
  DFF ram_reg_298__1_ ( .D(n18234), .CP(wclk), .Q(ram[13993]) );
  DFF ram_reg_298__0_ ( .D(n18233), .CP(wclk), .Q(ram[13992]) );
  DFF ram_reg_302__7_ ( .D(n18208), .CP(wclk), .Q(ram[13967]) );
  DFF ram_reg_302__6_ ( .D(n18207), .CP(wclk), .Q(ram[13966]) );
  DFF ram_reg_302__5_ ( .D(n18206), .CP(wclk), .Q(ram[13965]) );
  DFF ram_reg_302__4_ ( .D(n18205), .CP(wclk), .Q(ram[13964]) );
  DFF ram_reg_302__3_ ( .D(n18204), .CP(wclk), .Q(ram[13963]) );
  DFF ram_reg_302__2_ ( .D(n18203), .CP(wclk), .Q(ram[13962]) );
  DFF ram_reg_302__1_ ( .D(n18202), .CP(wclk), .Q(ram[13961]) );
  DFF ram_reg_302__0_ ( .D(n18201), .CP(wclk), .Q(ram[13960]) );
  DFF ram_reg_306__7_ ( .D(n18176), .CP(wclk), .Q(ram[13935]) );
  DFF ram_reg_306__6_ ( .D(n18175), .CP(wclk), .Q(ram[13934]) );
  DFF ram_reg_306__5_ ( .D(n18174), .CP(wclk), .Q(ram[13933]) );
  DFF ram_reg_306__4_ ( .D(n18173), .CP(wclk), .Q(ram[13932]) );
  DFF ram_reg_306__3_ ( .D(n18172), .CP(wclk), .Q(ram[13931]) );
  DFF ram_reg_306__2_ ( .D(n18171), .CP(wclk), .Q(ram[13930]) );
  DFF ram_reg_306__1_ ( .D(n18170), .CP(wclk), .Q(ram[13929]) );
  DFF ram_reg_306__0_ ( .D(n18169), .CP(wclk), .Q(ram[13928]) );
  DFF ram_reg_310__7_ ( .D(n18144), .CP(wclk), .Q(ram[13903]) );
  DFF ram_reg_310__6_ ( .D(n18143), .CP(wclk), .Q(ram[13902]) );
  DFF ram_reg_310__5_ ( .D(n18142), .CP(wclk), .Q(ram[13901]) );
  DFF ram_reg_310__4_ ( .D(n18141), .CP(wclk), .Q(ram[13900]) );
  DFF ram_reg_310__3_ ( .D(n18140), .CP(wclk), .Q(ram[13899]) );
  DFF ram_reg_310__2_ ( .D(n18139), .CP(wclk), .Q(ram[13898]) );
  DFF ram_reg_310__1_ ( .D(n18138), .CP(wclk), .Q(ram[13897]) );
  DFF ram_reg_310__0_ ( .D(n18137), .CP(wclk), .Q(ram[13896]) );
  DFF ram_reg_318__7_ ( .D(n18080), .CP(wclk), .Q(ram[13839]) );
  DFF ram_reg_318__6_ ( .D(n18079), .CP(wclk), .Q(ram[13838]) );
  DFF ram_reg_318__5_ ( .D(n18078), .CP(wclk), .Q(ram[13837]) );
  DFF ram_reg_318__4_ ( .D(n18077), .CP(wclk), .Q(ram[13836]) );
  DFF ram_reg_318__3_ ( .D(n18076), .CP(wclk), .Q(ram[13835]) );
  DFF ram_reg_318__2_ ( .D(n18075), .CP(wclk), .Q(ram[13834]) );
  DFF ram_reg_318__1_ ( .D(n18074), .CP(wclk), .Q(ram[13833]) );
  DFF ram_reg_318__0_ ( .D(n18073), .CP(wclk), .Q(ram[13832]) );
  DFF ram_reg_322__7_ ( .D(n18048), .CP(wclk), .Q(ram[13807]) );
  DFF ram_reg_322__6_ ( .D(n18047), .CP(wclk), .Q(ram[13806]) );
  DFF ram_reg_322__5_ ( .D(n18046), .CP(wclk), .Q(ram[13805]) );
  DFF ram_reg_322__4_ ( .D(n18045), .CP(wclk), .Q(ram[13804]) );
  DFF ram_reg_322__3_ ( .D(n18044), .CP(wclk), .Q(ram[13803]) );
  DFF ram_reg_322__2_ ( .D(n18043), .CP(wclk), .Q(ram[13802]) );
  DFF ram_reg_322__1_ ( .D(n18042), .CP(wclk), .Q(ram[13801]) );
  DFF ram_reg_322__0_ ( .D(n18041), .CP(wclk), .Q(ram[13800]) );
  DFF ram_reg_326__7_ ( .D(n18016), .CP(wclk), .Q(ram[13775]) );
  DFF ram_reg_326__6_ ( .D(n18015), .CP(wclk), .Q(ram[13774]) );
  DFF ram_reg_326__5_ ( .D(n18014), .CP(wclk), .Q(ram[13773]) );
  DFF ram_reg_326__4_ ( .D(n18013), .CP(wclk), .Q(ram[13772]) );
  DFF ram_reg_326__3_ ( .D(n18012), .CP(wclk), .Q(ram[13771]) );
  DFF ram_reg_326__2_ ( .D(n18011), .CP(wclk), .Q(ram[13770]) );
  DFF ram_reg_326__1_ ( .D(n18010), .CP(wclk), .Q(ram[13769]) );
  DFF ram_reg_326__0_ ( .D(n18009), .CP(wclk), .Q(ram[13768]) );
  DFF ram_reg_330__7_ ( .D(n17984), .CP(wclk), .Q(ram[13743]) );
  DFF ram_reg_330__6_ ( .D(n17983), .CP(wclk), .Q(ram[13742]) );
  DFF ram_reg_330__5_ ( .D(n17982), .CP(wclk), .Q(ram[13741]) );
  DFF ram_reg_330__4_ ( .D(n17981), .CP(wclk), .Q(ram[13740]) );
  DFF ram_reg_330__3_ ( .D(n17980), .CP(wclk), .Q(ram[13739]) );
  DFF ram_reg_330__2_ ( .D(n17979), .CP(wclk), .Q(ram[13738]) );
  DFF ram_reg_330__1_ ( .D(n17978), .CP(wclk), .Q(ram[13737]) );
  DFF ram_reg_330__0_ ( .D(n17977), .CP(wclk), .Q(ram[13736]) );
  DFF ram_reg_334__7_ ( .D(n17952), .CP(wclk), .Q(ram[13711]) );
  DFF ram_reg_334__6_ ( .D(n17951), .CP(wclk), .Q(ram[13710]) );
  DFF ram_reg_334__5_ ( .D(n17950), .CP(wclk), .Q(ram[13709]) );
  DFF ram_reg_334__4_ ( .D(n17949), .CP(wclk), .Q(ram[13708]) );
  DFF ram_reg_334__3_ ( .D(n17948), .CP(wclk), .Q(ram[13707]) );
  DFF ram_reg_334__2_ ( .D(n17947), .CP(wclk), .Q(ram[13706]) );
  DFF ram_reg_334__1_ ( .D(n17946), .CP(wclk), .Q(ram[13705]) );
  DFF ram_reg_334__0_ ( .D(n17945), .CP(wclk), .Q(ram[13704]) );
  DFF ram_reg_338__7_ ( .D(n17920), .CP(wclk), .Q(ram[13679]) );
  DFF ram_reg_338__6_ ( .D(n17919), .CP(wclk), .Q(ram[13678]) );
  DFF ram_reg_338__5_ ( .D(n17918), .CP(wclk), .Q(ram[13677]) );
  DFF ram_reg_338__4_ ( .D(n17917), .CP(wclk), .Q(ram[13676]) );
  DFF ram_reg_338__3_ ( .D(n17916), .CP(wclk), .Q(ram[13675]) );
  DFF ram_reg_338__2_ ( .D(n17915), .CP(wclk), .Q(ram[13674]) );
  DFF ram_reg_338__1_ ( .D(n17914), .CP(wclk), .Q(ram[13673]) );
  DFF ram_reg_338__0_ ( .D(n17913), .CP(wclk), .Q(ram[13672]) );
  DFF ram_reg_342__7_ ( .D(n17888), .CP(wclk), .Q(ram[13647]) );
  DFF ram_reg_342__6_ ( .D(n17887), .CP(wclk), .Q(ram[13646]) );
  DFF ram_reg_342__5_ ( .D(n17886), .CP(wclk), .Q(ram[13645]) );
  DFF ram_reg_342__4_ ( .D(n17885), .CP(wclk), .Q(ram[13644]) );
  DFF ram_reg_342__3_ ( .D(n17884), .CP(wclk), .Q(ram[13643]) );
  DFF ram_reg_342__2_ ( .D(n17883), .CP(wclk), .Q(ram[13642]) );
  DFF ram_reg_342__1_ ( .D(n17882), .CP(wclk), .Q(ram[13641]) );
  DFF ram_reg_342__0_ ( .D(n17881), .CP(wclk), .Q(ram[13640]) );
  DFF ram_reg_346__7_ ( .D(n17856), .CP(wclk), .Q(ram[13615]) );
  DFF ram_reg_346__6_ ( .D(n17855), .CP(wclk), .Q(ram[13614]) );
  DFF ram_reg_346__5_ ( .D(n17854), .CP(wclk), .Q(ram[13613]) );
  DFF ram_reg_346__4_ ( .D(n17853), .CP(wclk), .Q(ram[13612]) );
  DFF ram_reg_346__3_ ( .D(n17852), .CP(wclk), .Q(ram[13611]) );
  DFF ram_reg_346__2_ ( .D(n17851), .CP(wclk), .Q(ram[13610]) );
  DFF ram_reg_346__1_ ( .D(n17850), .CP(wclk), .Q(ram[13609]) );
  DFF ram_reg_346__0_ ( .D(n17849), .CP(wclk), .Q(ram[13608]) );
  DFF ram_reg_350__7_ ( .D(n17824), .CP(wclk), .Q(ram[13583]) );
  DFF ram_reg_350__6_ ( .D(n17823), .CP(wclk), .Q(ram[13582]) );
  DFF ram_reg_350__5_ ( .D(n17822), .CP(wclk), .Q(ram[13581]) );
  DFF ram_reg_350__4_ ( .D(n17821), .CP(wclk), .Q(ram[13580]) );
  DFF ram_reg_350__3_ ( .D(n17820), .CP(wclk), .Q(ram[13579]) );
  DFF ram_reg_350__2_ ( .D(n17819), .CP(wclk), .Q(ram[13578]) );
  DFF ram_reg_350__1_ ( .D(n17818), .CP(wclk), .Q(ram[13577]) );
  DFF ram_reg_350__0_ ( .D(n17817), .CP(wclk), .Q(ram[13576]) );
  DFF ram_reg_354__7_ ( .D(n17792), .CP(wclk), .Q(ram[13551]) );
  DFF ram_reg_354__6_ ( .D(n17791), .CP(wclk), .Q(ram[13550]) );
  DFF ram_reg_354__5_ ( .D(n17790), .CP(wclk), .Q(ram[13549]) );
  DFF ram_reg_354__4_ ( .D(n17789), .CP(wclk), .Q(ram[13548]) );
  DFF ram_reg_354__3_ ( .D(n17788), .CP(wclk), .Q(ram[13547]) );
  DFF ram_reg_354__2_ ( .D(n17787), .CP(wclk), .Q(ram[13546]) );
  DFF ram_reg_354__1_ ( .D(n17786), .CP(wclk), .Q(ram[13545]) );
  DFF ram_reg_354__0_ ( .D(n17785), .CP(wclk), .Q(ram[13544]) );
  DFF ram_reg_358__7_ ( .D(n17760), .CP(wclk), .Q(ram[13519]) );
  DFF ram_reg_358__6_ ( .D(n17759), .CP(wclk), .Q(ram[13518]) );
  DFF ram_reg_358__5_ ( .D(n17758), .CP(wclk), .Q(ram[13517]) );
  DFF ram_reg_358__4_ ( .D(n17757), .CP(wclk), .Q(ram[13516]) );
  DFF ram_reg_358__3_ ( .D(n17756), .CP(wclk), .Q(ram[13515]) );
  DFF ram_reg_358__2_ ( .D(n17755), .CP(wclk), .Q(ram[13514]) );
  DFF ram_reg_358__1_ ( .D(n17754), .CP(wclk), .Q(ram[13513]) );
  DFF ram_reg_358__0_ ( .D(n17753), .CP(wclk), .Q(ram[13512]) );
  DFF ram_reg_362__7_ ( .D(n17728), .CP(wclk), .Q(ram[13487]) );
  DFF ram_reg_362__6_ ( .D(n17727), .CP(wclk), .Q(ram[13486]) );
  DFF ram_reg_362__5_ ( .D(n17726), .CP(wclk), .Q(ram[13485]) );
  DFF ram_reg_362__4_ ( .D(n17725), .CP(wclk), .Q(ram[13484]) );
  DFF ram_reg_362__3_ ( .D(n17724), .CP(wclk), .Q(ram[13483]) );
  DFF ram_reg_362__2_ ( .D(n17723), .CP(wclk), .Q(ram[13482]) );
  DFF ram_reg_362__1_ ( .D(n17722), .CP(wclk), .Q(ram[13481]) );
  DFF ram_reg_362__0_ ( .D(n17721), .CP(wclk), .Q(ram[13480]) );
  DFF ram_reg_366__7_ ( .D(n17696), .CP(wclk), .Q(ram[13455]) );
  DFF ram_reg_366__6_ ( .D(n17695), .CP(wclk), .Q(ram[13454]) );
  DFF ram_reg_366__5_ ( .D(n17694), .CP(wclk), .Q(ram[13453]) );
  DFF ram_reg_366__4_ ( .D(n17693), .CP(wclk), .Q(ram[13452]) );
  DFF ram_reg_366__3_ ( .D(n17692), .CP(wclk), .Q(ram[13451]) );
  DFF ram_reg_366__2_ ( .D(n17691), .CP(wclk), .Q(ram[13450]) );
  DFF ram_reg_366__1_ ( .D(n17690), .CP(wclk), .Q(ram[13449]) );
  DFF ram_reg_366__0_ ( .D(n17689), .CP(wclk), .Q(ram[13448]) );
  DFF ram_reg_370__7_ ( .D(n17664), .CP(wclk), .Q(ram[13423]) );
  DFF ram_reg_370__6_ ( .D(n17663), .CP(wclk), .Q(ram[13422]) );
  DFF ram_reg_370__5_ ( .D(n17662), .CP(wclk), .Q(ram[13421]) );
  DFF ram_reg_370__4_ ( .D(n17661), .CP(wclk), .Q(ram[13420]) );
  DFF ram_reg_370__3_ ( .D(n17660), .CP(wclk), .Q(ram[13419]) );
  DFF ram_reg_370__2_ ( .D(n17659), .CP(wclk), .Q(ram[13418]) );
  DFF ram_reg_370__1_ ( .D(n17658), .CP(wclk), .Q(ram[13417]) );
  DFF ram_reg_370__0_ ( .D(n17657), .CP(wclk), .Q(ram[13416]) );
  DFF ram_reg_374__7_ ( .D(n17632), .CP(wclk), .Q(ram[13391]) );
  DFF ram_reg_374__6_ ( .D(n17631), .CP(wclk), .Q(ram[13390]) );
  DFF ram_reg_374__5_ ( .D(n17630), .CP(wclk), .Q(ram[13389]) );
  DFF ram_reg_374__4_ ( .D(n17629), .CP(wclk), .Q(ram[13388]) );
  DFF ram_reg_374__3_ ( .D(n17628), .CP(wclk), .Q(ram[13387]) );
  DFF ram_reg_374__2_ ( .D(n17627), .CP(wclk), .Q(ram[13386]) );
  DFF ram_reg_374__1_ ( .D(n17626), .CP(wclk), .Q(ram[13385]) );
  DFF ram_reg_374__0_ ( .D(n17625), .CP(wclk), .Q(ram[13384]) );
  DFF ram_reg_378__7_ ( .D(n17600), .CP(wclk), .Q(ram[13359]) );
  DFF ram_reg_378__6_ ( .D(n17599), .CP(wclk), .Q(ram[13358]) );
  DFF ram_reg_378__5_ ( .D(n17598), .CP(wclk), .Q(ram[13357]) );
  DFF ram_reg_378__4_ ( .D(n17597), .CP(wclk), .Q(ram[13356]) );
  DFF ram_reg_378__3_ ( .D(n17596), .CP(wclk), .Q(ram[13355]) );
  DFF ram_reg_378__2_ ( .D(n17595), .CP(wclk), .Q(ram[13354]) );
  DFF ram_reg_378__1_ ( .D(n17594), .CP(wclk), .Q(ram[13353]) );
  DFF ram_reg_378__0_ ( .D(n17593), .CP(wclk), .Q(ram[13352]) );
  DFF ram_reg_382__7_ ( .D(n17568), .CP(wclk), .Q(ram[13327]) );
  DFF ram_reg_382__6_ ( .D(n17567), .CP(wclk), .Q(ram[13326]) );
  DFF ram_reg_382__5_ ( .D(n17566), .CP(wclk), .Q(ram[13325]) );
  DFF ram_reg_382__4_ ( .D(n17565), .CP(wclk), .Q(ram[13324]) );
  DFF ram_reg_382__3_ ( .D(n17564), .CP(wclk), .Q(ram[13323]) );
  DFF ram_reg_382__2_ ( .D(n17563), .CP(wclk), .Q(ram[13322]) );
  DFF ram_reg_382__1_ ( .D(n17562), .CP(wclk), .Q(ram[13321]) );
  DFF ram_reg_382__0_ ( .D(n17561), .CP(wclk), .Q(ram[13320]) );
  DFF ram_reg_386__7_ ( .D(n17536), .CP(wclk), .Q(ram[13295]) );
  DFF ram_reg_386__6_ ( .D(n17535), .CP(wclk), .Q(ram[13294]) );
  DFF ram_reg_386__5_ ( .D(n17534), .CP(wclk), .Q(ram[13293]) );
  DFF ram_reg_386__4_ ( .D(n17533), .CP(wclk), .Q(ram[13292]) );
  DFF ram_reg_386__3_ ( .D(n17532), .CP(wclk), .Q(ram[13291]) );
  DFF ram_reg_386__2_ ( .D(n17531), .CP(wclk), .Q(ram[13290]) );
  DFF ram_reg_386__1_ ( .D(n17530), .CP(wclk), .Q(ram[13289]) );
  DFF ram_reg_386__0_ ( .D(n17529), .CP(wclk), .Q(ram[13288]) );
  DFF ram_reg_390__7_ ( .D(n17504), .CP(wclk), .Q(ram[13263]) );
  DFF ram_reg_390__6_ ( .D(n17503), .CP(wclk), .Q(ram[13262]) );
  DFF ram_reg_390__5_ ( .D(n17502), .CP(wclk), .Q(ram[13261]) );
  DFF ram_reg_390__4_ ( .D(n17501), .CP(wclk), .Q(ram[13260]) );
  DFF ram_reg_390__3_ ( .D(n17500), .CP(wclk), .Q(ram[13259]) );
  DFF ram_reg_390__2_ ( .D(n17499), .CP(wclk), .Q(ram[13258]) );
  DFF ram_reg_390__1_ ( .D(n17498), .CP(wclk), .Q(ram[13257]) );
  DFF ram_reg_390__0_ ( .D(n17497), .CP(wclk), .Q(ram[13256]) );
  DFF ram_reg_402__7_ ( .D(n17408), .CP(wclk), .Q(ram[13167]) );
  DFF ram_reg_402__6_ ( .D(n17407), .CP(wclk), .Q(ram[13166]) );
  DFF ram_reg_402__5_ ( .D(n17406), .CP(wclk), .Q(ram[13165]) );
  DFF ram_reg_402__4_ ( .D(n17405), .CP(wclk), .Q(ram[13164]) );
  DFF ram_reg_402__3_ ( .D(n17404), .CP(wclk), .Q(ram[13163]) );
  DFF ram_reg_402__2_ ( .D(n17403), .CP(wclk), .Q(ram[13162]) );
  DFF ram_reg_402__1_ ( .D(n17402), .CP(wclk), .Q(ram[13161]) );
  DFF ram_reg_402__0_ ( .D(n17401), .CP(wclk), .Q(ram[13160]) );
  DFF ram_reg_406__7_ ( .D(n17376), .CP(wclk), .Q(ram[13135]) );
  DFF ram_reg_406__6_ ( .D(n17375), .CP(wclk), .Q(ram[13134]) );
  DFF ram_reg_406__5_ ( .D(n17374), .CP(wclk), .Q(ram[13133]) );
  DFF ram_reg_406__4_ ( .D(n17373), .CP(wclk), .Q(ram[13132]) );
  DFF ram_reg_406__3_ ( .D(n17372), .CP(wclk), .Q(ram[13131]) );
  DFF ram_reg_406__2_ ( .D(n17371), .CP(wclk), .Q(ram[13130]) );
  DFF ram_reg_406__1_ ( .D(n17370), .CP(wclk), .Q(ram[13129]) );
  DFF ram_reg_406__0_ ( .D(n17369), .CP(wclk), .Q(ram[13128]) );
  DFF ram_reg_410__7_ ( .D(n17344), .CP(wclk), .Q(ram[13103]) );
  DFF ram_reg_410__6_ ( .D(n17343), .CP(wclk), .Q(ram[13102]) );
  DFF ram_reg_410__5_ ( .D(n17342), .CP(wclk), .Q(ram[13101]) );
  DFF ram_reg_410__4_ ( .D(n17341), .CP(wclk), .Q(ram[13100]) );
  DFF ram_reg_410__3_ ( .D(n17340), .CP(wclk), .Q(ram[13099]) );
  DFF ram_reg_410__2_ ( .D(n17339), .CP(wclk), .Q(ram[13098]) );
  DFF ram_reg_410__1_ ( .D(n17338), .CP(wclk), .Q(ram[13097]) );
  DFF ram_reg_410__0_ ( .D(n17337), .CP(wclk), .Q(ram[13096]) );
  DFF ram_reg_414__7_ ( .D(n17312), .CP(wclk), .Q(ram[13071]) );
  DFF ram_reg_414__6_ ( .D(n17311), .CP(wclk), .Q(ram[13070]) );
  DFF ram_reg_414__5_ ( .D(n17310), .CP(wclk), .Q(ram[13069]) );
  DFF ram_reg_414__4_ ( .D(n17309), .CP(wclk), .Q(ram[13068]) );
  DFF ram_reg_414__3_ ( .D(n17308), .CP(wclk), .Q(ram[13067]) );
  DFF ram_reg_414__2_ ( .D(n17307), .CP(wclk), .Q(ram[13066]) );
  DFF ram_reg_414__1_ ( .D(n17306), .CP(wclk), .Q(ram[13065]) );
  DFF ram_reg_414__0_ ( .D(n17305), .CP(wclk), .Q(ram[13064]) );
  DFF ram_reg_418__7_ ( .D(n17280), .CP(wclk), .Q(ram[13039]) );
  DFF ram_reg_418__6_ ( .D(n17279), .CP(wclk), .Q(ram[13038]) );
  DFF ram_reg_418__5_ ( .D(n17278), .CP(wclk), .Q(ram[13037]) );
  DFF ram_reg_418__4_ ( .D(n17277), .CP(wclk), .Q(ram[13036]) );
  DFF ram_reg_418__3_ ( .D(n17276), .CP(wclk), .Q(ram[13035]) );
  DFF ram_reg_418__2_ ( .D(n17275), .CP(wclk), .Q(ram[13034]) );
  DFF ram_reg_418__1_ ( .D(n17274), .CP(wclk), .Q(ram[13033]) );
  DFF ram_reg_418__0_ ( .D(n17273), .CP(wclk), .Q(ram[13032]) );
  DFF ram_reg_422__7_ ( .D(n17248), .CP(wclk), .Q(ram[13007]) );
  DFF ram_reg_422__6_ ( .D(n17247), .CP(wclk), .Q(ram[13006]) );
  DFF ram_reg_422__5_ ( .D(n17246), .CP(wclk), .Q(ram[13005]) );
  DFF ram_reg_422__4_ ( .D(n17245), .CP(wclk), .Q(ram[13004]) );
  DFF ram_reg_422__3_ ( .D(n17244), .CP(wclk), .Q(ram[13003]) );
  DFF ram_reg_422__2_ ( .D(n17243), .CP(wclk), .Q(ram[13002]) );
  DFF ram_reg_422__1_ ( .D(n17242), .CP(wclk), .Q(ram[13001]) );
  DFF ram_reg_422__0_ ( .D(n17241), .CP(wclk), .Q(ram[13000]) );
  DFF ram_reg_438__7_ ( .D(n17120), .CP(wclk), .Q(ram[12879]) );
  DFF ram_reg_438__6_ ( .D(n17119), .CP(wclk), .Q(ram[12878]) );
  DFF ram_reg_438__5_ ( .D(n17118), .CP(wclk), .Q(ram[12877]) );
  DFF ram_reg_438__4_ ( .D(n17117), .CP(wclk), .Q(ram[12876]) );
  DFF ram_reg_438__3_ ( .D(n17116), .CP(wclk), .Q(ram[12875]) );
  DFF ram_reg_438__2_ ( .D(n17115), .CP(wclk), .Q(ram[12874]) );
  DFF ram_reg_438__1_ ( .D(n17114), .CP(wclk), .Q(ram[12873]) );
  DFF ram_reg_438__0_ ( .D(n17113), .CP(wclk), .Q(ram[12872]) );
  DFF ram_reg_450__7_ ( .D(n17024), .CP(wclk), .Q(ram[12783]) );
  DFF ram_reg_450__6_ ( .D(n17023), .CP(wclk), .Q(ram[12782]) );
  DFF ram_reg_450__5_ ( .D(n17022), .CP(wclk), .Q(ram[12781]) );
  DFF ram_reg_450__4_ ( .D(n17021), .CP(wclk), .Q(ram[12780]) );
  DFF ram_reg_450__3_ ( .D(n17020), .CP(wclk), .Q(ram[12779]) );
  DFF ram_reg_450__2_ ( .D(n17019), .CP(wclk), .Q(ram[12778]) );
  DFF ram_reg_450__1_ ( .D(n17018), .CP(wclk), .Q(ram[12777]) );
  DFF ram_reg_450__0_ ( .D(n17017), .CP(wclk), .Q(ram[12776]) );
  DFF ram_reg_454__7_ ( .D(n16992), .CP(wclk), .Q(ram[12751]) );
  DFF ram_reg_454__6_ ( .D(n16991), .CP(wclk), .Q(ram[12750]) );
  DFF ram_reg_454__5_ ( .D(n16990), .CP(wclk), .Q(ram[12749]) );
  DFF ram_reg_454__4_ ( .D(n16989), .CP(wclk), .Q(ram[12748]) );
  DFF ram_reg_454__3_ ( .D(n16988), .CP(wclk), .Q(ram[12747]) );
  DFF ram_reg_454__2_ ( .D(n16987), .CP(wclk), .Q(ram[12746]) );
  DFF ram_reg_454__1_ ( .D(n16986), .CP(wclk), .Q(ram[12745]) );
  DFF ram_reg_454__0_ ( .D(n16985), .CP(wclk), .Q(ram[12744]) );
  DFF ram_reg_462__7_ ( .D(n16928), .CP(wclk), .Q(ram[12687]) );
  DFF ram_reg_462__6_ ( .D(n16927), .CP(wclk), .Q(ram[12686]) );
  DFF ram_reg_462__5_ ( .D(n16926), .CP(wclk), .Q(ram[12685]) );
  DFF ram_reg_462__4_ ( .D(n16925), .CP(wclk), .Q(ram[12684]) );
  DFF ram_reg_462__3_ ( .D(n16924), .CP(wclk), .Q(ram[12683]) );
  DFF ram_reg_462__2_ ( .D(n16923), .CP(wclk), .Q(ram[12682]) );
  DFF ram_reg_462__1_ ( .D(n16922), .CP(wclk), .Q(ram[12681]) );
  DFF ram_reg_462__0_ ( .D(n16921), .CP(wclk), .Q(ram[12680]) );
  DFF ram_reg_466__7_ ( .D(n16896), .CP(wclk), .Q(ram[12655]) );
  DFF ram_reg_466__6_ ( .D(n16895), .CP(wclk), .Q(ram[12654]) );
  DFF ram_reg_466__5_ ( .D(n16894), .CP(wclk), .Q(ram[12653]) );
  DFF ram_reg_466__4_ ( .D(n16893), .CP(wclk), .Q(ram[12652]) );
  DFF ram_reg_466__3_ ( .D(n16892), .CP(wclk), .Q(ram[12651]) );
  DFF ram_reg_466__2_ ( .D(n16891), .CP(wclk), .Q(ram[12650]) );
  DFF ram_reg_466__1_ ( .D(n16890), .CP(wclk), .Q(ram[12649]) );
  DFF ram_reg_466__0_ ( .D(n16889), .CP(wclk), .Q(ram[12648]) );
  DFF ram_reg_470__7_ ( .D(n16864), .CP(wclk), .Q(ram[12623]) );
  DFF ram_reg_470__6_ ( .D(n16863), .CP(wclk), .Q(ram[12622]) );
  DFF ram_reg_470__5_ ( .D(n16862), .CP(wclk), .Q(ram[12621]) );
  DFF ram_reg_470__4_ ( .D(n16861), .CP(wclk), .Q(ram[12620]) );
  DFF ram_reg_470__3_ ( .D(n16860), .CP(wclk), .Q(ram[12619]) );
  DFF ram_reg_470__2_ ( .D(n16859), .CP(wclk), .Q(ram[12618]) );
  DFF ram_reg_470__1_ ( .D(n16858), .CP(wclk), .Q(ram[12617]) );
  DFF ram_reg_470__0_ ( .D(n16857), .CP(wclk), .Q(ram[12616]) );
  DFF ram_reg_474__7_ ( .D(n16832), .CP(wclk), .Q(ram[12591]) );
  DFF ram_reg_474__6_ ( .D(n16831), .CP(wclk), .Q(ram[12590]) );
  DFF ram_reg_474__5_ ( .D(n16830), .CP(wclk), .Q(ram[12589]) );
  DFF ram_reg_474__4_ ( .D(n16829), .CP(wclk), .Q(ram[12588]) );
  DFF ram_reg_474__3_ ( .D(n16828), .CP(wclk), .Q(ram[12587]) );
  DFF ram_reg_474__2_ ( .D(n16827), .CP(wclk), .Q(ram[12586]) );
  DFF ram_reg_474__1_ ( .D(n16826), .CP(wclk), .Q(ram[12585]) );
  DFF ram_reg_474__0_ ( .D(n16825), .CP(wclk), .Q(ram[12584]) );
  DFF ram_reg_478__7_ ( .D(n16800), .CP(wclk), .Q(ram[12559]) );
  DFF ram_reg_478__6_ ( .D(n16799), .CP(wclk), .Q(ram[12558]) );
  DFF ram_reg_478__5_ ( .D(n16798), .CP(wclk), .Q(ram[12557]) );
  DFF ram_reg_478__4_ ( .D(n16797), .CP(wclk), .Q(ram[12556]) );
  DFF ram_reg_478__3_ ( .D(n16796), .CP(wclk), .Q(ram[12555]) );
  DFF ram_reg_478__2_ ( .D(n16795), .CP(wclk), .Q(ram[12554]) );
  DFF ram_reg_478__1_ ( .D(n16794), .CP(wclk), .Q(ram[12553]) );
  DFF ram_reg_478__0_ ( .D(n16793), .CP(wclk), .Q(ram[12552]) );
  DFF ram_reg_482__7_ ( .D(n16768), .CP(wclk), .Q(ram[12527]) );
  DFF ram_reg_482__6_ ( .D(n16767), .CP(wclk), .Q(ram[12526]) );
  DFF ram_reg_482__5_ ( .D(n16766), .CP(wclk), .Q(ram[12525]) );
  DFF ram_reg_482__4_ ( .D(n16765), .CP(wclk), .Q(ram[12524]) );
  DFF ram_reg_482__3_ ( .D(n16764), .CP(wclk), .Q(ram[12523]) );
  DFF ram_reg_482__2_ ( .D(n16763), .CP(wclk), .Q(ram[12522]) );
  DFF ram_reg_482__1_ ( .D(n16762), .CP(wclk), .Q(ram[12521]) );
  DFF ram_reg_482__0_ ( .D(n16761), .CP(wclk), .Q(ram[12520]) );
  DFF ram_reg_486__7_ ( .D(n16736), .CP(wclk), .Q(ram[12495]) );
  DFF ram_reg_486__6_ ( .D(n16735), .CP(wclk), .Q(ram[12494]) );
  DFF ram_reg_486__5_ ( .D(n16734), .CP(wclk), .Q(ram[12493]) );
  DFF ram_reg_486__4_ ( .D(n16733), .CP(wclk), .Q(ram[12492]) );
  DFF ram_reg_486__3_ ( .D(n16732), .CP(wclk), .Q(ram[12491]) );
  DFF ram_reg_486__2_ ( .D(n16731), .CP(wclk), .Q(ram[12490]) );
  DFF ram_reg_486__1_ ( .D(n16730), .CP(wclk), .Q(ram[12489]) );
  DFF ram_reg_486__0_ ( .D(n16729), .CP(wclk), .Q(ram[12488]) );
  DFF ram_reg_498__7_ ( .D(n16640), .CP(wclk), .Q(ram[12399]) );
  DFF ram_reg_498__6_ ( .D(n16639), .CP(wclk), .Q(ram[12398]) );
  DFF ram_reg_498__5_ ( .D(n16638), .CP(wclk), .Q(ram[12397]) );
  DFF ram_reg_498__4_ ( .D(n16637), .CP(wclk), .Q(ram[12396]) );
  DFF ram_reg_498__3_ ( .D(n16636), .CP(wclk), .Q(ram[12395]) );
  DFF ram_reg_498__2_ ( .D(n16635), .CP(wclk), .Q(ram[12394]) );
  DFF ram_reg_498__1_ ( .D(n16634), .CP(wclk), .Q(ram[12393]) );
  DFF ram_reg_498__0_ ( .D(n16633), .CP(wclk), .Q(ram[12392]) );
  DFF ram_reg_502__7_ ( .D(n16608), .CP(wclk), .Q(ram[12367]) );
  DFF ram_reg_502__6_ ( .D(n16607), .CP(wclk), .Q(ram[12366]) );
  DFF ram_reg_502__5_ ( .D(n16606), .CP(wclk), .Q(ram[12365]) );
  DFF ram_reg_502__4_ ( .D(n16605), .CP(wclk), .Q(ram[12364]) );
  DFF ram_reg_502__3_ ( .D(n16604), .CP(wclk), .Q(ram[12363]) );
  DFF ram_reg_502__2_ ( .D(n16603), .CP(wclk), .Q(ram[12362]) );
  DFF ram_reg_502__1_ ( .D(n16602), .CP(wclk), .Q(ram[12361]) );
  DFF ram_reg_502__0_ ( .D(n16601), .CP(wclk), .Q(ram[12360]) );
  DFF ram_reg_514__7_ ( .D(n16512), .CP(wclk), .Q(ram[12271]) );
  DFF ram_reg_514__6_ ( .D(n16511), .CP(wclk), .Q(ram[12270]) );
  DFF ram_reg_514__5_ ( .D(n16510), .CP(wclk), .Q(ram[12269]) );
  DFF ram_reg_514__4_ ( .D(n16509), .CP(wclk), .Q(ram[12268]) );
  DFF ram_reg_514__3_ ( .D(n16508), .CP(wclk), .Q(ram[12267]) );
  DFF ram_reg_514__2_ ( .D(n16507), .CP(wclk), .Q(ram[12266]) );
  DFF ram_reg_514__1_ ( .D(n16506), .CP(wclk), .Q(ram[12265]) );
  DFF ram_reg_514__0_ ( .D(n16505), .CP(wclk), .Q(ram[12264]) );
  DFF ram_reg_518__7_ ( .D(n16480), .CP(wclk), .Q(ram[12239]) );
  DFF ram_reg_518__6_ ( .D(n16479), .CP(wclk), .Q(ram[12238]) );
  DFF ram_reg_518__5_ ( .D(n16478), .CP(wclk), .Q(ram[12237]) );
  DFF ram_reg_518__4_ ( .D(n16477), .CP(wclk), .Q(ram[12236]) );
  DFF ram_reg_518__3_ ( .D(n16476), .CP(wclk), .Q(ram[12235]) );
  DFF ram_reg_518__2_ ( .D(n16475), .CP(wclk), .Q(ram[12234]) );
  DFF ram_reg_518__1_ ( .D(n16474), .CP(wclk), .Q(ram[12233]) );
  DFF ram_reg_518__0_ ( .D(n16473), .CP(wclk), .Q(ram[12232]) );
  DFF ram_reg_526__7_ ( .D(n16416), .CP(wclk), .Q(ram[12175]) );
  DFF ram_reg_526__6_ ( .D(n16415), .CP(wclk), .Q(ram[12174]) );
  DFF ram_reg_526__5_ ( .D(n16414), .CP(wclk), .Q(ram[12173]) );
  DFF ram_reg_526__4_ ( .D(n16413), .CP(wclk), .Q(ram[12172]) );
  DFF ram_reg_526__3_ ( .D(n16412), .CP(wclk), .Q(ram[12171]) );
  DFF ram_reg_526__2_ ( .D(n16411), .CP(wclk), .Q(ram[12170]) );
  DFF ram_reg_526__1_ ( .D(n16410), .CP(wclk), .Q(ram[12169]) );
  DFF ram_reg_526__0_ ( .D(n16409), .CP(wclk), .Q(ram[12168]) );
  DFF ram_reg_530__7_ ( .D(n16384), .CP(wclk), .Q(ram[12143]) );
  DFF ram_reg_530__6_ ( .D(n16383), .CP(wclk), .Q(ram[12142]) );
  DFF ram_reg_530__5_ ( .D(n16382), .CP(wclk), .Q(ram[12141]) );
  DFF ram_reg_530__4_ ( .D(n16381), .CP(wclk), .Q(ram[12140]) );
  DFF ram_reg_530__3_ ( .D(n16380), .CP(wclk), .Q(ram[12139]) );
  DFF ram_reg_530__2_ ( .D(n16379), .CP(wclk), .Q(ram[12138]) );
  DFF ram_reg_530__1_ ( .D(n16378), .CP(wclk), .Q(ram[12137]) );
  DFF ram_reg_530__0_ ( .D(n16377), .CP(wclk), .Q(ram[12136]) );
  DFF ram_reg_534__7_ ( .D(n16352), .CP(wclk), .Q(ram[12111]) );
  DFF ram_reg_534__6_ ( .D(n16351), .CP(wclk), .Q(ram[12110]) );
  DFF ram_reg_534__5_ ( .D(n16350), .CP(wclk), .Q(ram[12109]) );
  DFF ram_reg_534__4_ ( .D(n16349), .CP(wclk), .Q(ram[12108]) );
  DFF ram_reg_534__3_ ( .D(n16348), .CP(wclk), .Q(ram[12107]) );
  DFF ram_reg_534__2_ ( .D(n16347), .CP(wclk), .Q(ram[12106]) );
  DFF ram_reg_534__1_ ( .D(n16346), .CP(wclk), .Q(ram[12105]) );
  DFF ram_reg_534__0_ ( .D(n16345), .CP(wclk), .Q(ram[12104]) );
  DFF ram_reg_538__7_ ( .D(n16320), .CP(wclk), .Q(ram[12079]) );
  DFF ram_reg_538__6_ ( .D(n16319), .CP(wclk), .Q(ram[12078]) );
  DFF ram_reg_538__5_ ( .D(n16318), .CP(wclk), .Q(ram[12077]) );
  DFF ram_reg_538__4_ ( .D(n16317), .CP(wclk), .Q(ram[12076]) );
  DFF ram_reg_538__3_ ( .D(n16316), .CP(wclk), .Q(ram[12075]) );
  DFF ram_reg_538__2_ ( .D(n16315), .CP(wclk), .Q(ram[12074]) );
  DFF ram_reg_538__1_ ( .D(n16314), .CP(wclk), .Q(ram[12073]) );
  DFF ram_reg_538__0_ ( .D(n16313), .CP(wclk), .Q(ram[12072]) );
  DFF ram_reg_542__7_ ( .D(n16288), .CP(wclk), .Q(ram[12047]) );
  DFF ram_reg_542__6_ ( .D(n16287), .CP(wclk), .Q(ram[12046]) );
  DFF ram_reg_542__5_ ( .D(n16286), .CP(wclk), .Q(ram[12045]) );
  DFF ram_reg_542__4_ ( .D(n16285), .CP(wclk), .Q(ram[12044]) );
  DFF ram_reg_542__3_ ( .D(n16284), .CP(wclk), .Q(ram[12043]) );
  DFF ram_reg_542__2_ ( .D(n16283), .CP(wclk), .Q(ram[12042]) );
  DFF ram_reg_542__1_ ( .D(n16282), .CP(wclk), .Q(ram[12041]) );
  DFF ram_reg_542__0_ ( .D(n16281), .CP(wclk), .Q(ram[12040]) );
  DFF ram_reg_546__7_ ( .D(n16256), .CP(wclk), .Q(ram[12015]) );
  DFF ram_reg_546__6_ ( .D(n16255), .CP(wclk), .Q(ram[12014]) );
  DFF ram_reg_546__5_ ( .D(n16254), .CP(wclk), .Q(ram[12013]) );
  DFF ram_reg_546__4_ ( .D(n16253), .CP(wclk), .Q(ram[12012]) );
  DFF ram_reg_546__3_ ( .D(n16252), .CP(wclk), .Q(ram[12011]) );
  DFF ram_reg_546__2_ ( .D(n16251), .CP(wclk), .Q(ram[12010]) );
  DFF ram_reg_546__1_ ( .D(n16250), .CP(wclk), .Q(ram[12009]) );
  DFF ram_reg_546__0_ ( .D(n16249), .CP(wclk), .Q(ram[12008]) );
  DFF ram_reg_550__7_ ( .D(n16224), .CP(wclk), .Q(ram[11983]) );
  DFF ram_reg_550__6_ ( .D(n16223), .CP(wclk), .Q(ram[11982]) );
  DFF ram_reg_550__5_ ( .D(n16222), .CP(wclk), .Q(ram[11981]) );
  DFF ram_reg_550__4_ ( .D(n16221), .CP(wclk), .Q(ram[11980]) );
  DFF ram_reg_550__3_ ( .D(n16220), .CP(wclk), .Q(ram[11979]) );
  DFF ram_reg_550__2_ ( .D(n16219), .CP(wclk), .Q(ram[11978]) );
  DFF ram_reg_550__1_ ( .D(n16218), .CP(wclk), .Q(ram[11977]) );
  DFF ram_reg_550__0_ ( .D(n16217), .CP(wclk), .Q(ram[11976]) );
  DFF ram_reg_562__7_ ( .D(n16128), .CP(wclk), .Q(ram[11887]) );
  DFF ram_reg_562__6_ ( .D(n16127), .CP(wclk), .Q(ram[11886]) );
  DFF ram_reg_562__5_ ( .D(n16126), .CP(wclk), .Q(ram[11885]) );
  DFF ram_reg_562__4_ ( .D(n16125), .CP(wclk), .Q(ram[11884]) );
  DFF ram_reg_562__3_ ( .D(n16124), .CP(wclk), .Q(ram[11883]) );
  DFF ram_reg_562__2_ ( .D(n16123), .CP(wclk), .Q(ram[11882]) );
  DFF ram_reg_562__1_ ( .D(n16122), .CP(wclk), .Q(ram[11881]) );
  DFF ram_reg_562__0_ ( .D(n16121), .CP(wclk), .Q(ram[11880]) );
  DFF ram_reg_566__7_ ( .D(n16096), .CP(wclk), .Q(ram[11855]) );
  DFF ram_reg_566__6_ ( .D(n16095), .CP(wclk), .Q(ram[11854]) );
  DFF ram_reg_566__5_ ( .D(n16094), .CP(wclk), .Q(ram[11853]) );
  DFF ram_reg_566__4_ ( .D(n16093), .CP(wclk), .Q(ram[11852]) );
  DFF ram_reg_566__3_ ( .D(n16092), .CP(wclk), .Q(ram[11851]) );
  DFF ram_reg_566__2_ ( .D(n16091), .CP(wclk), .Q(ram[11850]) );
  DFF ram_reg_566__1_ ( .D(n16090), .CP(wclk), .Q(ram[11849]) );
  DFF ram_reg_566__0_ ( .D(n16089), .CP(wclk), .Q(ram[11848]) );
  DFF ram_reg_578__7_ ( .D(n16000), .CP(wclk), .Q(ram[11759]) );
  DFF ram_reg_578__6_ ( .D(n15999), .CP(wclk), .Q(ram[11758]) );
  DFF ram_reg_578__5_ ( .D(n15998), .CP(wclk), .Q(ram[11757]) );
  DFF ram_reg_578__4_ ( .D(n15997), .CP(wclk), .Q(ram[11756]) );
  DFF ram_reg_578__3_ ( .D(n15996), .CP(wclk), .Q(ram[11755]) );
  DFF ram_reg_578__2_ ( .D(n15995), .CP(wclk), .Q(ram[11754]) );
  DFF ram_reg_578__1_ ( .D(n15994), .CP(wclk), .Q(ram[11753]) );
  DFF ram_reg_578__0_ ( .D(n15993), .CP(wclk), .Q(ram[11752]) );
  DFF ram_reg_582__7_ ( .D(n15968), .CP(wclk), .Q(ram[11727]) );
  DFF ram_reg_582__6_ ( .D(n15967), .CP(wclk), .Q(ram[11726]) );
  DFF ram_reg_582__5_ ( .D(n15966), .CP(wclk), .Q(ram[11725]) );
  DFF ram_reg_582__4_ ( .D(n15965), .CP(wclk), .Q(ram[11724]) );
  DFF ram_reg_582__3_ ( .D(n15964), .CP(wclk), .Q(ram[11723]) );
  DFF ram_reg_582__2_ ( .D(n15963), .CP(wclk), .Q(ram[11722]) );
  DFF ram_reg_582__1_ ( .D(n15962), .CP(wclk), .Q(ram[11721]) );
  DFF ram_reg_582__0_ ( .D(n15961), .CP(wclk), .Q(ram[11720]) );
  DFF ram_reg_586__7_ ( .D(n15936), .CP(wclk), .Q(ram[11695]) );
  DFF ram_reg_586__6_ ( .D(n15935), .CP(wclk), .Q(ram[11694]) );
  DFF ram_reg_586__5_ ( .D(n15934), .CP(wclk), .Q(ram[11693]) );
  DFF ram_reg_586__4_ ( .D(n15933), .CP(wclk), .Q(ram[11692]) );
  DFF ram_reg_586__3_ ( .D(n15932), .CP(wclk), .Q(ram[11691]) );
  DFF ram_reg_586__2_ ( .D(n15931), .CP(wclk), .Q(ram[11690]) );
  DFF ram_reg_586__1_ ( .D(n15930), .CP(wclk), .Q(ram[11689]) );
  DFF ram_reg_586__0_ ( .D(n15929), .CP(wclk), .Q(ram[11688]) );
  DFF ram_reg_590__7_ ( .D(n15904), .CP(wclk), .Q(ram[11663]) );
  DFF ram_reg_590__6_ ( .D(n15903), .CP(wclk), .Q(ram[11662]) );
  DFF ram_reg_590__5_ ( .D(n15902), .CP(wclk), .Q(ram[11661]) );
  DFF ram_reg_590__4_ ( .D(n15901), .CP(wclk), .Q(ram[11660]) );
  DFF ram_reg_590__3_ ( .D(n15900), .CP(wclk), .Q(ram[11659]) );
  DFF ram_reg_590__2_ ( .D(n15899), .CP(wclk), .Q(ram[11658]) );
  DFF ram_reg_590__1_ ( .D(n15898), .CP(wclk), .Q(ram[11657]) );
  DFF ram_reg_590__0_ ( .D(n15897), .CP(wclk), .Q(ram[11656]) );
  DFF ram_reg_594__7_ ( .D(n15872), .CP(wclk), .Q(ram[11631]) );
  DFF ram_reg_594__6_ ( .D(n15871), .CP(wclk), .Q(ram[11630]) );
  DFF ram_reg_594__5_ ( .D(n15870), .CP(wclk), .Q(ram[11629]) );
  DFF ram_reg_594__4_ ( .D(n15869), .CP(wclk), .Q(ram[11628]) );
  DFF ram_reg_594__3_ ( .D(n15868), .CP(wclk), .Q(ram[11627]) );
  DFF ram_reg_594__2_ ( .D(n15867), .CP(wclk), .Q(ram[11626]) );
  DFF ram_reg_594__1_ ( .D(n15866), .CP(wclk), .Q(ram[11625]) );
  DFF ram_reg_594__0_ ( .D(n15865), .CP(wclk), .Q(ram[11624]) );
  DFF ram_reg_598__7_ ( .D(n15840), .CP(wclk), .Q(ram[11599]) );
  DFF ram_reg_598__6_ ( .D(n15839), .CP(wclk), .Q(ram[11598]) );
  DFF ram_reg_598__5_ ( .D(n15838), .CP(wclk), .Q(ram[11597]) );
  DFF ram_reg_598__4_ ( .D(n15837), .CP(wclk), .Q(ram[11596]) );
  DFF ram_reg_598__3_ ( .D(n15836), .CP(wclk), .Q(ram[11595]) );
  DFF ram_reg_598__2_ ( .D(n15835), .CP(wclk), .Q(ram[11594]) );
  DFF ram_reg_598__1_ ( .D(n15834), .CP(wclk), .Q(ram[11593]) );
  DFF ram_reg_598__0_ ( .D(n15833), .CP(wclk), .Q(ram[11592]) );
  DFF ram_reg_602__7_ ( .D(n15808), .CP(wclk), .Q(ram[11567]) );
  DFF ram_reg_602__6_ ( .D(n15807), .CP(wclk), .Q(ram[11566]) );
  DFF ram_reg_602__5_ ( .D(n15806), .CP(wclk), .Q(ram[11565]) );
  DFF ram_reg_602__4_ ( .D(n15805), .CP(wclk), .Q(ram[11564]) );
  DFF ram_reg_602__3_ ( .D(n15804), .CP(wclk), .Q(ram[11563]) );
  DFF ram_reg_602__2_ ( .D(n15803), .CP(wclk), .Q(ram[11562]) );
  DFF ram_reg_602__1_ ( .D(n15802), .CP(wclk), .Q(ram[11561]) );
  DFF ram_reg_602__0_ ( .D(n15801), .CP(wclk), .Q(ram[11560]) );
  DFF ram_reg_606__7_ ( .D(n15776), .CP(wclk), .Q(ram[11535]) );
  DFF ram_reg_606__6_ ( .D(n15775), .CP(wclk), .Q(ram[11534]) );
  DFF ram_reg_606__5_ ( .D(n15774), .CP(wclk), .Q(ram[11533]) );
  DFF ram_reg_606__4_ ( .D(n15773), .CP(wclk), .Q(ram[11532]) );
  DFF ram_reg_606__3_ ( .D(n15772), .CP(wclk), .Q(ram[11531]) );
  DFF ram_reg_606__2_ ( .D(n15771), .CP(wclk), .Q(ram[11530]) );
  DFF ram_reg_606__1_ ( .D(n15770), .CP(wclk), .Q(ram[11529]) );
  DFF ram_reg_606__0_ ( .D(n15769), .CP(wclk), .Q(ram[11528]) );
  DFF ram_reg_610__7_ ( .D(n15744), .CP(wclk), .Q(ram[11503]) );
  DFF ram_reg_610__6_ ( .D(n15743), .CP(wclk), .Q(ram[11502]) );
  DFF ram_reg_610__5_ ( .D(n15742), .CP(wclk), .Q(ram[11501]) );
  DFF ram_reg_610__4_ ( .D(n15741), .CP(wclk), .Q(ram[11500]) );
  DFF ram_reg_610__3_ ( .D(n15740), .CP(wclk), .Q(ram[11499]) );
  DFF ram_reg_610__2_ ( .D(n15739), .CP(wclk), .Q(ram[11498]) );
  DFF ram_reg_610__1_ ( .D(n15738), .CP(wclk), .Q(ram[11497]) );
  DFF ram_reg_610__0_ ( .D(n15737), .CP(wclk), .Q(ram[11496]) );
  DFF ram_reg_614__7_ ( .D(n15712), .CP(wclk), .Q(ram[11471]) );
  DFF ram_reg_614__6_ ( .D(n15711), .CP(wclk), .Q(ram[11470]) );
  DFF ram_reg_614__5_ ( .D(n15710), .CP(wclk), .Q(ram[11469]) );
  DFF ram_reg_614__4_ ( .D(n15709), .CP(wclk), .Q(ram[11468]) );
  DFF ram_reg_614__3_ ( .D(n15708), .CP(wclk), .Q(ram[11467]) );
  DFF ram_reg_614__2_ ( .D(n15707), .CP(wclk), .Q(ram[11466]) );
  DFF ram_reg_614__1_ ( .D(n15706), .CP(wclk), .Q(ram[11465]) );
  DFF ram_reg_614__0_ ( .D(n15705), .CP(wclk), .Q(ram[11464]) );
  DFF ram_reg_618__7_ ( .D(n15680), .CP(wclk), .Q(ram[11439]) );
  DFF ram_reg_618__6_ ( .D(n15679), .CP(wclk), .Q(ram[11438]) );
  DFF ram_reg_618__5_ ( .D(n15678), .CP(wclk), .Q(ram[11437]) );
  DFF ram_reg_618__4_ ( .D(n15677), .CP(wclk), .Q(ram[11436]) );
  DFF ram_reg_618__3_ ( .D(n15676), .CP(wclk), .Q(ram[11435]) );
  DFF ram_reg_618__2_ ( .D(n15675), .CP(wclk), .Q(ram[11434]) );
  DFF ram_reg_618__1_ ( .D(n15674), .CP(wclk), .Q(ram[11433]) );
  DFF ram_reg_618__0_ ( .D(n15673), .CP(wclk), .Q(ram[11432]) );
  DFF ram_reg_622__7_ ( .D(n15648), .CP(wclk), .Q(ram[11407]) );
  DFF ram_reg_622__6_ ( .D(n15647), .CP(wclk), .Q(ram[11406]) );
  DFF ram_reg_622__5_ ( .D(n15646), .CP(wclk), .Q(ram[11405]) );
  DFF ram_reg_622__4_ ( .D(n15645), .CP(wclk), .Q(ram[11404]) );
  DFF ram_reg_622__3_ ( .D(n15644), .CP(wclk), .Q(ram[11403]) );
  DFF ram_reg_622__2_ ( .D(n15643), .CP(wclk), .Q(ram[11402]) );
  DFF ram_reg_622__1_ ( .D(n15642), .CP(wclk), .Q(ram[11401]) );
  DFF ram_reg_622__0_ ( .D(n15641), .CP(wclk), .Q(ram[11400]) );
  DFF ram_reg_626__7_ ( .D(n15616), .CP(wclk), .Q(ram[11375]) );
  DFF ram_reg_626__6_ ( .D(n15615), .CP(wclk), .Q(ram[11374]) );
  DFF ram_reg_626__5_ ( .D(n15614), .CP(wclk), .Q(ram[11373]) );
  DFF ram_reg_626__4_ ( .D(n15613), .CP(wclk), .Q(ram[11372]) );
  DFF ram_reg_626__3_ ( .D(n15612), .CP(wclk), .Q(ram[11371]) );
  DFF ram_reg_626__2_ ( .D(n15611), .CP(wclk), .Q(ram[11370]) );
  DFF ram_reg_626__1_ ( .D(n15610), .CP(wclk), .Q(ram[11369]) );
  DFF ram_reg_626__0_ ( .D(n15609), .CP(wclk), .Q(ram[11368]) );
  DFF ram_reg_630__7_ ( .D(n15584), .CP(wclk), .Q(ram[11343]) );
  DFF ram_reg_630__6_ ( .D(n15583), .CP(wclk), .Q(ram[11342]) );
  DFF ram_reg_630__5_ ( .D(n15582), .CP(wclk), .Q(ram[11341]) );
  DFF ram_reg_630__4_ ( .D(n15581), .CP(wclk), .Q(ram[11340]) );
  DFF ram_reg_630__3_ ( .D(n15580), .CP(wclk), .Q(ram[11339]) );
  DFF ram_reg_630__2_ ( .D(n15579), .CP(wclk), .Q(ram[11338]) );
  DFF ram_reg_630__1_ ( .D(n15578), .CP(wclk), .Q(ram[11337]) );
  DFF ram_reg_630__0_ ( .D(n15577), .CP(wclk), .Q(ram[11336]) );
  DFF ram_reg_634__7_ ( .D(n15552), .CP(wclk), .Q(ram[11311]) );
  DFF ram_reg_634__6_ ( .D(n15551), .CP(wclk), .Q(ram[11310]) );
  DFF ram_reg_634__5_ ( .D(n15550), .CP(wclk), .Q(ram[11309]) );
  DFF ram_reg_634__4_ ( .D(n15549), .CP(wclk), .Q(ram[11308]) );
  DFF ram_reg_634__3_ ( .D(n15548), .CP(wclk), .Q(ram[11307]) );
  DFF ram_reg_634__2_ ( .D(n15547), .CP(wclk), .Q(ram[11306]) );
  DFF ram_reg_634__1_ ( .D(n15546), .CP(wclk), .Q(ram[11305]) );
  DFF ram_reg_634__0_ ( .D(n15545), .CP(wclk), .Q(ram[11304]) );
  DFF ram_reg_638__7_ ( .D(n15520), .CP(wclk), .Q(ram[11279]) );
  DFF ram_reg_638__6_ ( .D(n15519), .CP(wclk), .Q(ram[11278]) );
  DFF ram_reg_638__5_ ( .D(n15518), .CP(wclk), .Q(ram[11277]) );
  DFF ram_reg_638__4_ ( .D(n15517), .CP(wclk), .Q(ram[11276]) );
  DFF ram_reg_638__3_ ( .D(n15516), .CP(wclk), .Q(ram[11275]) );
  DFF ram_reg_638__2_ ( .D(n15515), .CP(wclk), .Q(ram[11274]) );
  DFF ram_reg_638__1_ ( .D(n15514), .CP(wclk), .Q(ram[11273]) );
  DFF ram_reg_638__0_ ( .D(n15513), .CP(wclk), .Q(ram[11272]) );
  DFF ram_reg_646__7_ ( .D(n15456), .CP(wclk), .Q(ram[11215]) );
  DFF ram_reg_646__6_ ( .D(n15455), .CP(wclk), .Q(ram[11214]) );
  DFF ram_reg_646__5_ ( .D(n15454), .CP(wclk), .Q(ram[11213]) );
  DFF ram_reg_646__4_ ( .D(n15453), .CP(wclk), .Q(ram[11212]) );
  DFF ram_reg_646__3_ ( .D(n15452), .CP(wclk), .Q(ram[11211]) );
  DFF ram_reg_646__2_ ( .D(n15451), .CP(wclk), .Q(ram[11210]) );
  DFF ram_reg_646__1_ ( .D(n15450), .CP(wclk), .Q(ram[11209]) );
  DFF ram_reg_646__0_ ( .D(n15449), .CP(wclk), .Q(ram[11208]) );
  DFF ram_reg_658__7_ ( .D(n15360), .CP(wclk), .Q(ram[11119]) );
  DFF ram_reg_658__6_ ( .D(n15359), .CP(wclk), .Q(ram[11118]) );
  DFF ram_reg_658__5_ ( .D(n15358), .CP(wclk), .Q(ram[11117]) );
  DFF ram_reg_658__4_ ( .D(n15357), .CP(wclk), .Q(ram[11116]) );
  DFF ram_reg_658__3_ ( .D(n15356), .CP(wclk), .Q(ram[11115]) );
  DFF ram_reg_658__2_ ( .D(n15355), .CP(wclk), .Q(ram[11114]) );
  DFF ram_reg_658__1_ ( .D(n15354), .CP(wclk), .Q(ram[11113]) );
  DFF ram_reg_658__0_ ( .D(n15353), .CP(wclk), .Q(ram[11112]) );
  DFF ram_reg_662__7_ ( .D(n15328), .CP(wclk), .Q(ram[11087]) );
  DFF ram_reg_662__6_ ( .D(n15327), .CP(wclk), .Q(ram[11086]) );
  DFF ram_reg_662__5_ ( .D(n15326), .CP(wclk), .Q(ram[11085]) );
  DFF ram_reg_662__4_ ( .D(n15325), .CP(wclk), .Q(ram[11084]) );
  DFF ram_reg_662__3_ ( .D(n15324), .CP(wclk), .Q(ram[11083]) );
  DFF ram_reg_662__2_ ( .D(n15323), .CP(wclk), .Q(ram[11082]) );
  DFF ram_reg_662__1_ ( .D(n15322), .CP(wclk), .Q(ram[11081]) );
  DFF ram_reg_662__0_ ( .D(n15321), .CP(wclk), .Q(ram[11080]) );
  DFF ram_reg_678__7_ ( .D(n15200), .CP(wclk), .Q(ram[10959]) );
  DFF ram_reg_678__6_ ( .D(n15199), .CP(wclk), .Q(ram[10958]) );
  DFF ram_reg_678__5_ ( .D(n15198), .CP(wclk), .Q(ram[10957]) );
  DFF ram_reg_678__4_ ( .D(n15197), .CP(wclk), .Q(ram[10956]) );
  DFF ram_reg_678__3_ ( .D(n15196), .CP(wclk), .Q(ram[10955]) );
  DFF ram_reg_678__2_ ( .D(n15195), .CP(wclk), .Q(ram[10954]) );
  DFF ram_reg_678__1_ ( .D(n15194), .CP(wclk), .Q(ram[10953]) );
  DFF ram_reg_678__0_ ( .D(n15193), .CP(wclk), .Q(ram[10952]) );
  DFF ram_reg_694__7_ ( .D(n15072), .CP(wclk), .Q(ram[10831]) );
  DFF ram_reg_694__6_ ( .D(n15071), .CP(wclk), .Q(ram[10830]) );
  DFF ram_reg_694__5_ ( .D(n15070), .CP(wclk), .Q(ram[10829]) );
  DFF ram_reg_694__4_ ( .D(n15069), .CP(wclk), .Q(ram[10828]) );
  DFF ram_reg_694__3_ ( .D(n15068), .CP(wclk), .Q(ram[10827]) );
  DFF ram_reg_694__2_ ( .D(n15067), .CP(wclk), .Q(ram[10826]) );
  DFF ram_reg_694__1_ ( .D(n15066), .CP(wclk), .Q(ram[10825]) );
  DFF ram_reg_694__0_ ( .D(n15065), .CP(wclk), .Q(ram[10824]) );
  DFF ram_reg_706__7_ ( .D(n14976), .CP(wclk), .Q(ram[10735]) );
  DFF ram_reg_706__6_ ( .D(n14975), .CP(wclk), .Q(ram[10734]) );
  DFF ram_reg_706__5_ ( .D(n14974), .CP(wclk), .Q(ram[10733]) );
  DFF ram_reg_706__4_ ( .D(n14973), .CP(wclk), .Q(ram[10732]) );
  DFF ram_reg_706__3_ ( .D(n14972), .CP(wclk), .Q(ram[10731]) );
  DFF ram_reg_706__2_ ( .D(n14971), .CP(wclk), .Q(ram[10730]) );
  DFF ram_reg_706__1_ ( .D(n14970), .CP(wclk), .Q(ram[10729]) );
  DFF ram_reg_706__0_ ( .D(n14969), .CP(wclk), .Q(ram[10728]) );
  DFF ram_reg_710__7_ ( .D(n14944), .CP(wclk), .Q(ram[10703]) );
  DFF ram_reg_710__6_ ( .D(n14943), .CP(wclk), .Q(ram[10702]) );
  DFF ram_reg_710__5_ ( .D(n14942), .CP(wclk), .Q(ram[10701]) );
  DFF ram_reg_710__4_ ( .D(n14941), .CP(wclk), .Q(ram[10700]) );
  DFF ram_reg_710__3_ ( .D(n14940), .CP(wclk), .Q(ram[10699]) );
  DFF ram_reg_710__2_ ( .D(n14939), .CP(wclk), .Q(ram[10698]) );
  DFF ram_reg_710__1_ ( .D(n14938), .CP(wclk), .Q(ram[10697]) );
  DFF ram_reg_710__0_ ( .D(n14937), .CP(wclk), .Q(ram[10696]) );
  DFF ram_reg_722__7_ ( .D(n14848), .CP(wclk), .Q(ram[10607]) );
  DFF ram_reg_722__6_ ( .D(n14847), .CP(wclk), .Q(ram[10606]) );
  DFF ram_reg_722__5_ ( .D(n14846), .CP(wclk), .Q(ram[10605]) );
  DFF ram_reg_722__4_ ( .D(n14845), .CP(wclk), .Q(ram[10604]) );
  DFF ram_reg_722__3_ ( .D(n14844), .CP(wclk), .Q(ram[10603]) );
  DFF ram_reg_722__2_ ( .D(n14843), .CP(wclk), .Q(ram[10602]) );
  DFF ram_reg_722__1_ ( .D(n14842), .CP(wclk), .Q(ram[10601]) );
  DFF ram_reg_722__0_ ( .D(n14841), .CP(wclk), .Q(ram[10600]) );
  DFF ram_reg_726__7_ ( .D(n14816), .CP(wclk), .Q(ram[10575]) );
  DFF ram_reg_726__6_ ( .D(n14815), .CP(wclk), .Q(ram[10574]) );
  DFF ram_reg_726__5_ ( .D(n14814), .CP(wclk), .Q(ram[10573]) );
  DFF ram_reg_726__4_ ( .D(n14813), .CP(wclk), .Q(ram[10572]) );
  DFF ram_reg_726__3_ ( .D(n14812), .CP(wclk), .Q(ram[10571]) );
  DFF ram_reg_726__2_ ( .D(n14811), .CP(wclk), .Q(ram[10570]) );
  DFF ram_reg_726__1_ ( .D(n14810), .CP(wclk), .Q(ram[10569]) );
  DFF ram_reg_726__0_ ( .D(n14809), .CP(wclk), .Q(ram[10568]) );
  DFF ram_reg_734__7_ ( .D(n14752), .CP(wclk), .Q(ram[10511]) );
  DFF ram_reg_734__6_ ( .D(n14751), .CP(wclk), .Q(ram[10510]) );
  DFF ram_reg_734__5_ ( .D(n14750), .CP(wclk), .Q(ram[10509]) );
  DFF ram_reg_734__4_ ( .D(n14749), .CP(wclk), .Q(ram[10508]) );
  DFF ram_reg_734__3_ ( .D(n14748), .CP(wclk), .Q(ram[10507]) );
  DFF ram_reg_734__2_ ( .D(n14747), .CP(wclk), .Q(ram[10506]) );
  DFF ram_reg_734__1_ ( .D(n14746), .CP(wclk), .Q(ram[10505]) );
  DFF ram_reg_734__0_ ( .D(n14745), .CP(wclk), .Q(ram[10504]) );
  DFF ram_reg_742__7_ ( .D(n14688), .CP(wclk), .Q(ram[10447]) );
  DFF ram_reg_742__6_ ( .D(n14687), .CP(wclk), .Q(ram[10446]) );
  DFF ram_reg_742__5_ ( .D(n14686), .CP(wclk), .Q(ram[10445]) );
  DFF ram_reg_742__4_ ( .D(n14685), .CP(wclk), .Q(ram[10444]) );
  DFF ram_reg_742__3_ ( .D(n14684), .CP(wclk), .Q(ram[10443]) );
  DFF ram_reg_742__2_ ( .D(n14683), .CP(wclk), .Q(ram[10442]) );
  DFF ram_reg_742__1_ ( .D(n14682), .CP(wclk), .Q(ram[10441]) );
  DFF ram_reg_742__0_ ( .D(n14681), .CP(wclk), .Q(ram[10440]) );
  DFF ram_reg_758__7_ ( .D(n14560), .CP(wclk), .Q(ram[10319]) );
  DFF ram_reg_758__6_ ( .D(n14559), .CP(wclk), .Q(ram[10318]) );
  DFF ram_reg_758__5_ ( .D(n14558), .CP(wclk), .Q(ram[10317]) );
  DFF ram_reg_758__4_ ( .D(n14557), .CP(wclk), .Q(ram[10316]) );
  DFF ram_reg_758__3_ ( .D(n14556), .CP(wclk), .Q(ram[10315]) );
  DFF ram_reg_758__2_ ( .D(n14555), .CP(wclk), .Q(ram[10314]) );
  DFF ram_reg_758__1_ ( .D(n14554), .CP(wclk), .Q(ram[10313]) );
  DFF ram_reg_758__0_ ( .D(n14553), .CP(wclk), .Q(ram[10312]) );
  DFF ram_reg_770__7_ ( .D(n14464), .CP(wclk), .Q(ram[10223]) );
  DFF ram_reg_770__6_ ( .D(n14463), .CP(wclk), .Q(ram[10222]) );
  DFF ram_reg_770__5_ ( .D(n14462), .CP(wclk), .Q(ram[10221]) );
  DFF ram_reg_770__4_ ( .D(n14461), .CP(wclk), .Q(ram[10220]) );
  DFF ram_reg_770__3_ ( .D(n14460), .CP(wclk), .Q(ram[10219]) );
  DFF ram_reg_770__2_ ( .D(n14459), .CP(wclk), .Q(ram[10218]) );
  DFF ram_reg_770__1_ ( .D(n14458), .CP(wclk), .Q(ram[10217]) );
  DFF ram_reg_770__0_ ( .D(n14457), .CP(wclk), .Q(ram[10216]) );
  DFF ram_reg_774__7_ ( .D(n14432), .CP(wclk), .Q(ram[10191]) );
  DFF ram_reg_774__6_ ( .D(n14431), .CP(wclk), .Q(ram[10190]) );
  DFF ram_reg_774__5_ ( .D(n14430), .CP(wclk), .Q(ram[10189]) );
  DFF ram_reg_774__4_ ( .D(n14429), .CP(wclk), .Q(ram[10188]) );
  DFF ram_reg_774__3_ ( .D(n14428), .CP(wclk), .Q(ram[10187]) );
  DFF ram_reg_774__2_ ( .D(n14427), .CP(wclk), .Q(ram[10186]) );
  DFF ram_reg_774__1_ ( .D(n14426), .CP(wclk), .Q(ram[10185]) );
  DFF ram_reg_774__0_ ( .D(n14425), .CP(wclk), .Q(ram[10184]) );
  DFF ram_reg_782__7_ ( .D(n14368), .CP(wclk), .Q(ram[10127]) );
  DFF ram_reg_782__6_ ( .D(n14367), .CP(wclk), .Q(ram[10126]) );
  DFF ram_reg_782__5_ ( .D(n14366), .CP(wclk), .Q(ram[10125]) );
  DFF ram_reg_782__4_ ( .D(n14365), .CP(wclk), .Q(ram[10124]) );
  DFF ram_reg_782__3_ ( .D(n14364), .CP(wclk), .Q(ram[10123]) );
  DFF ram_reg_782__2_ ( .D(n14363), .CP(wclk), .Q(ram[10122]) );
  DFF ram_reg_782__1_ ( .D(n14362), .CP(wclk), .Q(ram[10121]) );
  DFF ram_reg_782__0_ ( .D(n14361), .CP(wclk), .Q(ram[10120]) );
  DFF ram_reg_786__7_ ( .D(n14336), .CP(wclk), .Q(ram[10095]) );
  DFF ram_reg_786__6_ ( .D(n14335), .CP(wclk), .Q(ram[10094]) );
  DFF ram_reg_786__5_ ( .D(n14334), .CP(wclk), .Q(ram[10093]) );
  DFF ram_reg_786__4_ ( .D(n14333), .CP(wclk), .Q(ram[10092]) );
  DFF ram_reg_786__3_ ( .D(n14332), .CP(wclk), .Q(ram[10091]) );
  DFF ram_reg_786__2_ ( .D(n14331), .CP(wclk), .Q(ram[10090]) );
  DFF ram_reg_786__1_ ( .D(n14330), .CP(wclk), .Q(ram[10089]) );
  DFF ram_reg_786__0_ ( .D(n14329), .CP(wclk), .Q(ram[10088]) );
  DFF ram_reg_790__7_ ( .D(n14304), .CP(wclk), .Q(ram[10063]) );
  DFF ram_reg_790__6_ ( .D(n14303), .CP(wclk), .Q(ram[10062]) );
  DFF ram_reg_790__5_ ( .D(n14302), .CP(wclk), .Q(ram[10061]) );
  DFF ram_reg_790__4_ ( .D(n14301), .CP(wclk), .Q(ram[10060]) );
  DFF ram_reg_790__3_ ( .D(n14300), .CP(wclk), .Q(ram[10059]) );
  DFF ram_reg_790__2_ ( .D(n14299), .CP(wclk), .Q(ram[10058]) );
  DFF ram_reg_790__1_ ( .D(n14298), .CP(wclk), .Q(ram[10057]) );
  DFF ram_reg_790__0_ ( .D(n14297), .CP(wclk), .Q(ram[10056]) );
  DFF ram_reg_794__7_ ( .D(n14272), .CP(wclk), .Q(ram[10031]) );
  DFF ram_reg_794__6_ ( .D(n14271), .CP(wclk), .Q(ram[10030]) );
  DFF ram_reg_794__5_ ( .D(n14270), .CP(wclk), .Q(ram[10029]) );
  DFF ram_reg_794__4_ ( .D(n14269), .CP(wclk), .Q(ram[10028]) );
  DFF ram_reg_794__3_ ( .D(n14268), .CP(wclk), .Q(ram[10027]) );
  DFF ram_reg_794__2_ ( .D(n14267), .CP(wclk), .Q(ram[10026]) );
  DFF ram_reg_794__1_ ( .D(n14266), .CP(wclk), .Q(ram[10025]) );
  DFF ram_reg_794__0_ ( .D(n14265), .CP(wclk), .Q(ram[10024]) );
  DFF ram_reg_798__7_ ( .D(n14240), .CP(wclk), .Q(ram[9999]) );
  DFF ram_reg_798__6_ ( .D(n14239), .CP(wclk), .Q(ram[9998]) );
  DFF ram_reg_798__5_ ( .D(n14238), .CP(wclk), .Q(ram[9997]) );
  DFF ram_reg_798__4_ ( .D(n14237), .CP(wclk), .Q(ram[9996]) );
  DFF ram_reg_798__3_ ( .D(n14236), .CP(wclk), .Q(ram[9995]) );
  DFF ram_reg_798__2_ ( .D(n14235), .CP(wclk), .Q(ram[9994]) );
  DFF ram_reg_798__1_ ( .D(n14234), .CP(wclk), .Q(ram[9993]) );
  DFF ram_reg_798__0_ ( .D(n14233), .CP(wclk), .Q(ram[9992]) );
  DFF ram_reg_802__7_ ( .D(n14208), .CP(wclk), .Q(ram[9967]) );
  DFF ram_reg_802__6_ ( .D(n14207), .CP(wclk), .Q(ram[9966]) );
  DFF ram_reg_802__5_ ( .D(n14206), .CP(wclk), .Q(ram[9965]) );
  DFF ram_reg_802__4_ ( .D(n14205), .CP(wclk), .Q(ram[9964]) );
  DFF ram_reg_802__3_ ( .D(n14204), .CP(wclk), .Q(ram[9963]) );
  DFF ram_reg_802__2_ ( .D(n14203), .CP(wclk), .Q(ram[9962]) );
  DFF ram_reg_802__1_ ( .D(n14202), .CP(wclk), .Q(ram[9961]) );
  DFF ram_reg_802__0_ ( .D(n14201), .CP(wclk), .Q(ram[9960]) );
  DFF ram_reg_806__7_ ( .D(n14176), .CP(wclk), .Q(ram[9935]) );
  DFF ram_reg_806__6_ ( .D(n14175), .CP(wclk), .Q(ram[9934]) );
  DFF ram_reg_806__5_ ( .D(n14174), .CP(wclk), .Q(ram[9933]) );
  DFF ram_reg_806__4_ ( .D(n14173), .CP(wclk), .Q(ram[9932]) );
  DFF ram_reg_806__3_ ( .D(n14172), .CP(wclk), .Q(ram[9931]) );
  DFF ram_reg_806__2_ ( .D(n14171), .CP(wclk), .Q(ram[9930]) );
  DFF ram_reg_806__1_ ( .D(n14170), .CP(wclk), .Q(ram[9929]) );
  DFF ram_reg_806__0_ ( .D(n14169), .CP(wclk), .Q(ram[9928]) );
  DFF ram_reg_818__7_ ( .D(n14080), .CP(wclk), .Q(ram[9839]) );
  DFF ram_reg_818__6_ ( .D(n14079), .CP(wclk), .Q(ram[9838]) );
  DFF ram_reg_818__5_ ( .D(n14078), .CP(wclk), .Q(ram[9837]) );
  DFF ram_reg_818__4_ ( .D(n14077), .CP(wclk), .Q(ram[9836]) );
  DFF ram_reg_818__3_ ( .D(n14076), .CP(wclk), .Q(ram[9835]) );
  DFF ram_reg_818__2_ ( .D(n14075), .CP(wclk), .Q(ram[9834]) );
  DFF ram_reg_818__1_ ( .D(n14074), .CP(wclk), .Q(ram[9833]) );
  DFF ram_reg_818__0_ ( .D(n14073), .CP(wclk), .Q(ram[9832]) );
  DFF ram_reg_822__7_ ( .D(n14048), .CP(wclk), .Q(ram[9807]) );
  DFF ram_reg_822__6_ ( .D(n14047), .CP(wclk), .Q(ram[9806]) );
  DFF ram_reg_822__5_ ( .D(n14046), .CP(wclk), .Q(ram[9805]) );
  DFF ram_reg_822__4_ ( .D(n14045), .CP(wclk), .Q(ram[9804]) );
  DFF ram_reg_822__3_ ( .D(n14044), .CP(wclk), .Q(ram[9803]) );
  DFF ram_reg_822__2_ ( .D(n14043), .CP(wclk), .Q(ram[9802]) );
  DFF ram_reg_822__1_ ( .D(n14042), .CP(wclk), .Q(ram[9801]) );
  DFF ram_reg_822__0_ ( .D(n14041), .CP(wclk), .Q(ram[9800]) );
  DFF ram_reg_834__7_ ( .D(n13952), .CP(wclk), .Q(ram[9711]) );
  DFF ram_reg_834__6_ ( .D(n13951), .CP(wclk), .Q(ram[9710]) );
  DFF ram_reg_834__5_ ( .D(n13950), .CP(wclk), .Q(ram[9709]) );
  DFF ram_reg_834__4_ ( .D(n13949), .CP(wclk), .Q(ram[9708]) );
  DFF ram_reg_834__3_ ( .D(n13948), .CP(wclk), .Q(ram[9707]) );
  DFF ram_reg_834__2_ ( .D(n13947), .CP(wclk), .Q(ram[9706]) );
  DFF ram_reg_834__1_ ( .D(n13946), .CP(wclk), .Q(ram[9705]) );
  DFF ram_reg_834__0_ ( .D(n13945), .CP(wclk), .Q(ram[9704]) );
  DFF ram_reg_838__7_ ( .D(n13920), .CP(wclk), .Q(ram[9679]) );
  DFF ram_reg_838__6_ ( .D(n13919), .CP(wclk), .Q(ram[9678]) );
  DFF ram_reg_838__5_ ( .D(n13918), .CP(wclk), .Q(ram[9677]) );
  DFF ram_reg_838__4_ ( .D(n13917), .CP(wclk), .Q(ram[9676]) );
  DFF ram_reg_838__3_ ( .D(n13916), .CP(wclk), .Q(ram[9675]) );
  DFF ram_reg_838__2_ ( .D(n13915), .CP(wclk), .Q(ram[9674]) );
  DFF ram_reg_838__1_ ( .D(n13914), .CP(wclk), .Q(ram[9673]) );
  DFF ram_reg_838__0_ ( .D(n13913), .CP(wclk), .Q(ram[9672]) );
  DFF ram_reg_842__7_ ( .D(n13888), .CP(wclk), .Q(ram[9647]) );
  DFF ram_reg_842__6_ ( .D(n13887), .CP(wclk), .Q(ram[9646]) );
  DFF ram_reg_842__5_ ( .D(n13886), .CP(wclk), .Q(ram[9645]) );
  DFF ram_reg_842__4_ ( .D(n13885), .CP(wclk), .Q(ram[9644]) );
  DFF ram_reg_842__3_ ( .D(n13884), .CP(wclk), .Q(ram[9643]) );
  DFF ram_reg_842__2_ ( .D(n13883), .CP(wclk), .Q(ram[9642]) );
  DFF ram_reg_842__1_ ( .D(n13882), .CP(wclk), .Q(ram[9641]) );
  DFF ram_reg_842__0_ ( .D(n13881), .CP(wclk), .Q(ram[9640]) );
  DFF ram_reg_846__7_ ( .D(n13856), .CP(wclk), .Q(ram[9615]) );
  DFF ram_reg_846__6_ ( .D(n13855), .CP(wclk), .Q(ram[9614]) );
  DFF ram_reg_846__5_ ( .D(n13854), .CP(wclk), .Q(ram[9613]) );
  DFF ram_reg_846__4_ ( .D(n13853), .CP(wclk), .Q(ram[9612]) );
  DFF ram_reg_846__3_ ( .D(n13852), .CP(wclk), .Q(ram[9611]) );
  DFF ram_reg_846__2_ ( .D(n13851), .CP(wclk), .Q(ram[9610]) );
  DFF ram_reg_846__1_ ( .D(n13850), .CP(wclk), .Q(ram[9609]) );
  DFF ram_reg_846__0_ ( .D(n13849), .CP(wclk), .Q(ram[9608]) );
  DFF ram_reg_850__7_ ( .D(n13824), .CP(wclk), .Q(ram[9583]) );
  DFF ram_reg_850__6_ ( .D(n13823), .CP(wclk), .Q(ram[9582]) );
  DFF ram_reg_850__5_ ( .D(n13822), .CP(wclk), .Q(ram[9581]) );
  DFF ram_reg_850__4_ ( .D(n13821), .CP(wclk), .Q(ram[9580]) );
  DFF ram_reg_850__3_ ( .D(n13820), .CP(wclk), .Q(ram[9579]) );
  DFF ram_reg_850__2_ ( .D(n13819), .CP(wclk), .Q(ram[9578]) );
  DFF ram_reg_850__1_ ( .D(n13818), .CP(wclk), .Q(ram[9577]) );
  DFF ram_reg_850__0_ ( .D(n13817), .CP(wclk), .Q(ram[9576]) );
  DFF ram_reg_854__7_ ( .D(n13792), .CP(wclk), .Q(ram[9551]) );
  DFF ram_reg_854__6_ ( .D(n13791), .CP(wclk), .Q(ram[9550]) );
  DFF ram_reg_854__5_ ( .D(n13790), .CP(wclk), .Q(ram[9549]) );
  DFF ram_reg_854__4_ ( .D(n13789), .CP(wclk), .Q(ram[9548]) );
  DFF ram_reg_854__3_ ( .D(n13788), .CP(wclk), .Q(ram[9547]) );
  DFF ram_reg_854__2_ ( .D(n13787), .CP(wclk), .Q(ram[9546]) );
  DFF ram_reg_854__1_ ( .D(n13786), .CP(wclk), .Q(ram[9545]) );
  DFF ram_reg_854__0_ ( .D(n13785), .CP(wclk), .Q(ram[9544]) );
  DFF ram_reg_858__7_ ( .D(n13760), .CP(wclk), .Q(ram[9519]) );
  DFF ram_reg_858__6_ ( .D(n13759), .CP(wclk), .Q(ram[9518]) );
  DFF ram_reg_858__5_ ( .D(n13758), .CP(wclk), .Q(ram[9517]) );
  DFF ram_reg_858__4_ ( .D(n13757), .CP(wclk), .Q(ram[9516]) );
  DFF ram_reg_858__3_ ( .D(n13756), .CP(wclk), .Q(ram[9515]) );
  DFF ram_reg_858__2_ ( .D(n13755), .CP(wclk), .Q(ram[9514]) );
  DFF ram_reg_858__1_ ( .D(n13754), .CP(wclk), .Q(ram[9513]) );
  DFF ram_reg_858__0_ ( .D(n13753), .CP(wclk), .Q(ram[9512]) );
  DFF ram_reg_862__7_ ( .D(n13728), .CP(wclk), .Q(ram[9487]) );
  DFF ram_reg_862__6_ ( .D(n13727), .CP(wclk), .Q(ram[9486]) );
  DFF ram_reg_862__5_ ( .D(n13726), .CP(wclk), .Q(ram[9485]) );
  DFF ram_reg_862__4_ ( .D(n13725), .CP(wclk), .Q(ram[9484]) );
  DFF ram_reg_862__3_ ( .D(n13724), .CP(wclk), .Q(ram[9483]) );
  DFF ram_reg_862__2_ ( .D(n13723), .CP(wclk), .Q(ram[9482]) );
  DFF ram_reg_862__1_ ( .D(n13722), .CP(wclk), .Q(ram[9481]) );
  DFF ram_reg_862__0_ ( .D(n13721), .CP(wclk), .Q(ram[9480]) );
  DFF ram_reg_866__7_ ( .D(n13696), .CP(wclk), .Q(ram[9455]) );
  DFF ram_reg_866__6_ ( .D(n13695), .CP(wclk), .Q(ram[9454]) );
  DFF ram_reg_866__5_ ( .D(n13694), .CP(wclk), .Q(ram[9453]) );
  DFF ram_reg_866__4_ ( .D(n13693), .CP(wclk), .Q(ram[9452]) );
  DFF ram_reg_866__3_ ( .D(n13692), .CP(wclk), .Q(ram[9451]) );
  DFF ram_reg_866__2_ ( .D(n13691), .CP(wclk), .Q(ram[9450]) );
  DFF ram_reg_866__1_ ( .D(n13690), .CP(wclk), .Q(ram[9449]) );
  DFF ram_reg_866__0_ ( .D(n13689), .CP(wclk), .Q(ram[9448]) );
  DFF ram_reg_870__7_ ( .D(n13664), .CP(wclk), .Q(ram[9423]) );
  DFF ram_reg_870__6_ ( .D(n13663), .CP(wclk), .Q(ram[9422]) );
  DFF ram_reg_870__5_ ( .D(n13662), .CP(wclk), .Q(ram[9421]) );
  DFF ram_reg_870__4_ ( .D(n13661), .CP(wclk), .Q(ram[9420]) );
  DFF ram_reg_870__3_ ( .D(n13660), .CP(wclk), .Q(ram[9419]) );
  DFF ram_reg_870__2_ ( .D(n13659), .CP(wclk), .Q(ram[9418]) );
  DFF ram_reg_870__1_ ( .D(n13658), .CP(wclk), .Q(ram[9417]) );
  DFF ram_reg_870__0_ ( .D(n13657), .CP(wclk), .Q(ram[9416]) );
  DFF ram_reg_874__7_ ( .D(n13632), .CP(wclk), .Q(ram[9391]) );
  DFF ram_reg_874__6_ ( .D(n13631), .CP(wclk), .Q(ram[9390]) );
  DFF ram_reg_874__5_ ( .D(n13630), .CP(wclk), .Q(ram[9389]) );
  DFF ram_reg_874__4_ ( .D(n13629), .CP(wclk), .Q(ram[9388]) );
  DFF ram_reg_874__3_ ( .D(n13628), .CP(wclk), .Q(ram[9387]) );
  DFF ram_reg_874__2_ ( .D(n13627), .CP(wclk), .Q(ram[9386]) );
  DFF ram_reg_874__1_ ( .D(n13626), .CP(wclk), .Q(ram[9385]) );
  DFF ram_reg_874__0_ ( .D(n13625), .CP(wclk), .Q(ram[9384]) );
  DFF ram_reg_878__7_ ( .D(n13600), .CP(wclk), .Q(ram[9359]) );
  DFF ram_reg_878__6_ ( .D(n13599), .CP(wclk), .Q(ram[9358]) );
  DFF ram_reg_878__5_ ( .D(n13598), .CP(wclk), .Q(ram[9357]) );
  DFF ram_reg_878__4_ ( .D(n13597), .CP(wclk), .Q(ram[9356]) );
  DFF ram_reg_878__3_ ( .D(n13596), .CP(wclk), .Q(ram[9355]) );
  DFF ram_reg_878__2_ ( .D(n13595), .CP(wclk), .Q(ram[9354]) );
  DFF ram_reg_878__1_ ( .D(n13594), .CP(wclk), .Q(ram[9353]) );
  DFF ram_reg_878__0_ ( .D(n13593), .CP(wclk), .Q(ram[9352]) );
  DFF ram_reg_882__7_ ( .D(n13568), .CP(wclk), .Q(ram[9327]) );
  DFF ram_reg_882__6_ ( .D(n13567), .CP(wclk), .Q(ram[9326]) );
  DFF ram_reg_882__5_ ( .D(n13566), .CP(wclk), .Q(ram[9325]) );
  DFF ram_reg_882__4_ ( .D(n13565), .CP(wclk), .Q(ram[9324]) );
  DFF ram_reg_882__3_ ( .D(n13564), .CP(wclk), .Q(ram[9323]) );
  DFF ram_reg_882__2_ ( .D(n13563), .CP(wclk), .Q(ram[9322]) );
  DFF ram_reg_882__1_ ( .D(n13562), .CP(wclk), .Q(ram[9321]) );
  DFF ram_reg_882__0_ ( .D(n13561), .CP(wclk), .Q(ram[9320]) );
  DFF ram_reg_886__7_ ( .D(n13536), .CP(wclk), .Q(ram[9295]) );
  DFF ram_reg_886__6_ ( .D(n13535), .CP(wclk), .Q(ram[9294]) );
  DFF ram_reg_886__5_ ( .D(n13534), .CP(wclk), .Q(ram[9293]) );
  DFF ram_reg_886__4_ ( .D(n13533), .CP(wclk), .Q(ram[9292]) );
  DFF ram_reg_886__3_ ( .D(n13532), .CP(wclk), .Q(ram[9291]) );
  DFF ram_reg_886__2_ ( .D(n13531), .CP(wclk), .Q(ram[9290]) );
  DFF ram_reg_886__1_ ( .D(n13530), .CP(wclk), .Q(ram[9289]) );
  DFF ram_reg_886__0_ ( .D(n13529), .CP(wclk), .Q(ram[9288]) );
  DFF ram_reg_890__7_ ( .D(n13504), .CP(wclk), .Q(ram[9263]) );
  DFF ram_reg_890__6_ ( .D(n13503), .CP(wclk), .Q(ram[9262]) );
  DFF ram_reg_890__5_ ( .D(n13502), .CP(wclk), .Q(ram[9261]) );
  DFF ram_reg_890__4_ ( .D(n13501), .CP(wclk), .Q(ram[9260]) );
  DFF ram_reg_890__3_ ( .D(n13500), .CP(wclk), .Q(ram[9259]) );
  DFF ram_reg_890__2_ ( .D(n13499), .CP(wclk), .Q(ram[9258]) );
  DFF ram_reg_890__1_ ( .D(n13498), .CP(wclk), .Q(ram[9257]) );
  DFF ram_reg_890__0_ ( .D(n13497), .CP(wclk), .Q(ram[9256]) );
  DFF ram_reg_894__7_ ( .D(n13472), .CP(wclk), .Q(ram[9231]) );
  DFF ram_reg_894__6_ ( .D(n13471), .CP(wclk), .Q(ram[9230]) );
  DFF ram_reg_894__5_ ( .D(n13470), .CP(wclk), .Q(ram[9229]) );
  DFF ram_reg_894__4_ ( .D(n13469), .CP(wclk), .Q(ram[9228]) );
  DFF ram_reg_894__3_ ( .D(n13468), .CP(wclk), .Q(ram[9227]) );
  DFF ram_reg_894__2_ ( .D(n13467), .CP(wclk), .Q(ram[9226]) );
  DFF ram_reg_894__1_ ( .D(n13466), .CP(wclk), .Q(ram[9225]) );
  DFF ram_reg_894__0_ ( .D(n13465), .CP(wclk), .Q(ram[9224]) );
  DFF ram_reg_902__7_ ( .D(n13408), .CP(wclk), .Q(ram[9167]) );
  DFF ram_reg_902__6_ ( .D(n13407), .CP(wclk), .Q(ram[9166]) );
  DFF ram_reg_902__5_ ( .D(n13406), .CP(wclk), .Q(ram[9165]) );
  DFF ram_reg_902__4_ ( .D(n13405), .CP(wclk), .Q(ram[9164]) );
  DFF ram_reg_902__3_ ( .D(n13404), .CP(wclk), .Q(ram[9163]) );
  DFF ram_reg_902__2_ ( .D(n13403), .CP(wclk), .Q(ram[9162]) );
  DFF ram_reg_902__1_ ( .D(n13402), .CP(wclk), .Q(ram[9161]) );
  DFF ram_reg_902__0_ ( .D(n13401), .CP(wclk), .Q(ram[9160]) );
  DFF ram_reg_914__7_ ( .D(n13312), .CP(wclk), .Q(ram[9071]) );
  DFF ram_reg_914__6_ ( .D(n13311), .CP(wclk), .Q(ram[9070]) );
  DFF ram_reg_914__5_ ( .D(n13310), .CP(wclk), .Q(ram[9069]) );
  DFF ram_reg_914__4_ ( .D(n13309), .CP(wclk), .Q(ram[9068]) );
  DFF ram_reg_914__3_ ( .D(n13308), .CP(wclk), .Q(ram[9067]) );
  DFF ram_reg_914__2_ ( .D(n13307), .CP(wclk), .Q(ram[9066]) );
  DFF ram_reg_914__1_ ( .D(n13306), .CP(wclk), .Q(ram[9065]) );
  DFF ram_reg_914__0_ ( .D(n13305), .CP(wclk), .Q(ram[9064]) );
  DFF ram_reg_918__7_ ( .D(n13280), .CP(wclk), .Q(ram[9039]) );
  DFF ram_reg_918__6_ ( .D(n13279), .CP(wclk), .Q(ram[9038]) );
  DFF ram_reg_918__5_ ( .D(n13278), .CP(wclk), .Q(ram[9037]) );
  DFF ram_reg_918__4_ ( .D(n13277), .CP(wclk), .Q(ram[9036]) );
  DFF ram_reg_918__3_ ( .D(n13276), .CP(wclk), .Q(ram[9035]) );
  DFF ram_reg_918__2_ ( .D(n13275), .CP(wclk), .Q(ram[9034]) );
  DFF ram_reg_918__1_ ( .D(n13274), .CP(wclk), .Q(ram[9033]) );
  DFF ram_reg_918__0_ ( .D(n13273), .CP(wclk), .Q(ram[9032]) );
  DFF ram_reg_934__7_ ( .D(n13152), .CP(wclk), .Q(ram[8911]) );
  DFF ram_reg_934__6_ ( .D(n13151), .CP(wclk), .Q(ram[8910]) );
  DFF ram_reg_934__5_ ( .D(n13150), .CP(wclk), .Q(ram[8909]) );
  DFF ram_reg_934__4_ ( .D(n13149), .CP(wclk), .Q(ram[8908]) );
  DFF ram_reg_934__3_ ( .D(n13148), .CP(wclk), .Q(ram[8907]) );
  DFF ram_reg_934__2_ ( .D(n13147), .CP(wclk), .Q(ram[8906]) );
  DFF ram_reg_934__1_ ( .D(n13146), .CP(wclk), .Q(ram[8905]) );
  DFF ram_reg_934__0_ ( .D(n13145), .CP(wclk), .Q(ram[8904]) );
  DFF ram_reg_950__7_ ( .D(n13024), .CP(wclk), .Q(ram[8783]) );
  DFF ram_reg_950__6_ ( .D(n13023), .CP(wclk), .Q(ram[8782]) );
  DFF ram_reg_950__5_ ( .D(n13022), .CP(wclk), .Q(ram[8781]) );
  DFF ram_reg_950__4_ ( .D(n13021), .CP(wclk), .Q(ram[8780]) );
  DFF ram_reg_950__3_ ( .D(n13020), .CP(wclk), .Q(ram[8779]) );
  DFF ram_reg_950__2_ ( .D(n13019), .CP(wclk), .Q(ram[8778]) );
  DFF ram_reg_950__1_ ( .D(n13018), .CP(wclk), .Q(ram[8777]) );
  DFF ram_reg_950__0_ ( .D(n13017), .CP(wclk), .Q(ram[8776]) );
  DFF ram_reg_962__7_ ( .D(n12928), .CP(wclk), .Q(ram[8687]) );
  DFF ram_reg_962__6_ ( .D(n12927), .CP(wclk), .Q(ram[8686]) );
  DFF ram_reg_962__5_ ( .D(n12926), .CP(wclk), .Q(ram[8685]) );
  DFF ram_reg_962__4_ ( .D(n12925), .CP(wclk), .Q(ram[8684]) );
  DFF ram_reg_962__3_ ( .D(n12924), .CP(wclk), .Q(ram[8683]) );
  DFF ram_reg_962__2_ ( .D(n12923), .CP(wclk), .Q(ram[8682]) );
  DFF ram_reg_962__1_ ( .D(n12922), .CP(wclk), .Q(ram[8681]) );
  DFF ram_reg_962__0_ ( .D(n12921), .CP(wclk), .Q(ram[8680]) );
  DFF ram_reg_966__7_ ( .D(n12896), .CP(wclk), .Q(ram[8655]) );
  DFF ram_reg_966__6_ ( .D(n12895), .CP(wclk), .Q(ram[8654]) );
  DFF ram_reg_966__5_ ( .D(n12894), .CP(wclk), .Q(ram[8653]) );
  DFF ram_reg_966__4_ ( .D(n12893), .CP(wclk), .Q(ram[8652]) );
  DFF ram_reg_966__3_ ( .D(n12892), .CP(wclk), .Q(ram[8651]) );
  DFF ram_reg_966__2_ ( .D(n12891), .CP(wclk), .Q(ram[8650]) );
  DFF ram_reg_966__1_ ( .D(n12890), .CP(wclk), .Q(ram[8649]) );
  DFF ram_reg_966__0_ ( .D(n12889), .CP(wclk), .Q(ram[8648]) );
  DFF ram_reg_978__7_ ( .D(n12800), .CP(wclk), .Q(ram[8559]) );
  DFF ram_reg_978__6_ ( .D(n12799), .CP(wclk), .Q(ram[8558]) );
  DFF ram_reg_978__5_ ( .D(n12798), .CP(wclk), .Q(ram[8557]) );
  DFF ram_reg_978__4_ ( .D(n12797), .CP(wclk), .Q(ram[8556]) );
  DFF ram_reg_978__3_ ( .D(n12796), .CP(wclk), .Q(ram[8555]) );
  DFF ram_reg_978__2_ ( .D(n12795), .CP(wclk), .Q(ram[8554]) );
  DFF ram_reg_978__1_ ( .D(n12794), .CP(wclk), .Q(ram[8553]) );
  DFF ram_reg_978__0_ ( .D(n12793), .CP(wclk), .Q(ram[8552]) );
  DFF ram_reg_982__7_ ( .D(n12768), .CP(wclk), .Q(ram[8527]) );
  DFF ram_reg_982__6_ ( .D(n12767), .CP(wclk), .Q(ram[8526]) );
  DFF ram_reg_982__5_ ( .D(n12766), .CP(wclk), .Q(ram[8525]) );
  DFF ram_reg_982__4_ ( .D(n12765), .CP(wclk), .Q(ram[8524]) );
  DFF ram_reg_982__3_ ( .D(n12764), .CP(wclk), .Q(ram[8523]) );
  DFF ram_reg_982__2_ ( .D(n12763), .CP(wclk), .Q(ram[8522]) );
  DFF ram_reg_982__1_ ( .D(n12762), .CP(wclk), .Q(ram[8521]) );
  DFF ram_reg_982__0_ ( .D(n12761), .CP(wclk), .Q(ram[8520]) );
  DFF ram_reg_998__7_ ( .D(n12640), .CP(wclk), .Q(ram[8399]) );
  DFF ram_reg_998__6_ ( .D(n12639), .CP(wclk), .Q(ram[8398]) );
  DFF ram_reg_998__5_ ( .D(n12638), .CP(wclk), .Q(ram[8397]) );
  DFF ram_reg_998__4_ ( .D(n12637), .CP(wclk), .Q(ram[8396]) );
  DFF ram_reg_998__3_ ( .D(n12636), .CP(wclk), .Q(ram[8395]) );
  DFF ram_reg_998__2_ ( .D(n12635), .CP(wclk), .Q(ram[8394]) );
  DFF ram_reg_998__1_ ( .D(n12634), .CP(wclk), .Q(ram[8393]) );
  DFF ram_reg_998__0_ ( .D(n12633), .CP(wclk), .Q(ram[8392]) );
  DFF ram_reg_1014__7_ ( .D(n12512), .CP(wclk), .Q(ram[8271]) );
  DFF ram_reg_1014__6_ ( .D(n12511), .CP(wclk), .Q(ram[8270]) );
  DFF ram_reg_1014__5_ ( .D(n12510), .CP(wclk), .Q(ram[8269]) );
  DFF ram_reg_1014__4_ ( .D(n12509), .CP(wclk), .Q(ram[8268]) );
  DFF ram_reg_1014__3_ ( .D(n12508), .CP(wclk), .Q(ram[8267]) );
  DFF ram_reg_1014__2_ ( .D(n12507), .CP(wclk), .Q(ram[8266]) );
  DFF ram_reg_1014__1_ ( .D(n12506), .CP(wclk), .Q(ram[8265]) );
  DFF ram_reg_1014__0_ ( .D(n12505), .CP(wclk), .Q(ram[8264]) );
  DFF ram_reg_1026__7_ ( .D(n12416), .CP(wclk), .Q(ram[8175]) );
  DFF ram_reg_1026__6_ ( .D(n12415), .CP(wclk), .Q(ram[8174]) );
  DFF ram_reg_1026__5_ ( .D(n12414), .CP(wclk), .Q(ram[8173]) );
  DFF ram_reg_1026__4_ ( .D(n12413), .CP(wclk), .Q(ram[8172]) );
  DFF ram_reg_1026__3_ ( .D(n12412), .CP(wclk), .Q(ram[8171]) );
  DFF ram_reg_1026__2_ ( .D(n12411), .CP(wclk), .Q(ram[8170]) );
  DFF ram_reg_1026__1_ ( .D(n12410), .CP(wclk), .Q(ram[8169]) );
  DFF ram_reg_1026__0_ ( .D(n12409), .CP(wclk), .Q(ram[8168]) );
  DFF ram_reg_1030__7_ ( .D(n12384), .CP(wclk), .Q(ram[8143]) );
  DFF ram_reg_1030__6_ ( .D(n12383), .CP(wclk), .Q(ram[8142]) );
  DFF ram_reg_1030__5_ ( .D(n12382), .CP(wclk), .Q(ram[8141]) );
  DFF ram_reg_1030__4_ ( .D(n12381), .CP(wclk), .Q(ram[8140]) );
  DFF ram_reg_1030__3_ ( .D(n12380), .CP(wclk), .Q(ram[8139]) );
  DFF ram_reg_1030__2_ ( .D(n12379), .CP(wclk), .Q(ram[8138]) );
  DFF ram_reg_1030__1_ ( .D(n12378), .CP(wclk), .Q(ram[8137]) );
  DFF ram_reg_1030__0_ ( .D(n12377), .CP(wclk), .Q(ram[8136]) );
  DFF ram_reg_1034__7_ ( .D(n12352), .CP(wclk), .Q(ram[8111]) );
  DFF ram_reg_1034__6_ ( .D(n12351), .CP(wclk), .Q(ram[8110]) );
  DFF ram_reg_1034__5_ ( .D(n12350), .CP(wclk), .Q(ram[8109]) );
  DFF ram_reg_1034__4_ ( .D(n12349), .CP(wclk), .Q(ram[8108]) );
  DFF ram_reg_1034__3_ ( .D(n12348), .CP(wclk), .Q(ram[8107]) );
  DFF ram_reg_1034__2_ ( .D(n12347), .CP(wclk), .Q(ram[8106]) );
  DFF ram_reg_1034__1_ ( .D(n12346), .CP(wclk), .Q(ram[8105]) );
  DFF ram_reg_1034__0_ ( .D(n12345), .CP(wclk), .Q(ram[8104]) );
  DFF ram_reg_1038__7_ ( .D(n12320), .CP(wclk), .Q(ram[8079]) );
  DFF ram_reg_1038__6_ ( .D(n12319), .CP(wclk), .Q(ram[8078]) );
  DFF ram_reg_1038__5_ ( .D(n12318), .CP(wclk), .Q(ram[8077]) );
  DFF ram_reg_1038__4_ ( .D(n12317), .CP(wclk), .Q(ram[8076]) );
  DFF ram_reg_1038__3_ ( .D(n12316), .CP(wclk), .Q(ram[8075]) );
  DFF ram_reg_1038__2_ ( .D(n12315), .CP(wclk), .Q(ram[8074]) );
  DFF ram_reg_1038__1_ ( .D(n12314), .CP(wclk), .Q(ram[8073]) );
  DFF ram_reg_1038__0_ ( .D(n12313), .CP(wclk), .Q(ram[8072]) );
  DFF ram_reg_1042__7_ ( .D(n12288), .CP(wclk), .Q(ram[8047]) );
  DFF ram_reg_1042__6_ ( .D(n12287), .CP(wclk), .Q(ram[8046]) );
  DFF ram_reg_1042__5_ ( .D(n12286), .CP(wclk), .Q(ram[8045]) );
  DFF ram_reg_1042__4_ ( .D(n12285), .CP(wclk), .Q(ram[8044]) );
  DFF ram_reg_1042__3_ ( .D(n12284), .CP(wclk), .Q(ram[8043]) );
  DFF ram_reg_1042__2_ ( .D(n12283), .CP(wclk), .Q(ram[8042]) );
  DFF ram_reg_1042__1_ ( .D(n12282), .CP(wclk), .Q(ram[8041]) );
  DFF ram_reg_1042__0_ ( .D(n12281), .CP(wclk), .Q(ram[8040]) );
  DFF ram_reg_1046__7_ ( .D(n12256), .CP(wclk), .Q(ram[8015]) );
  DFF ram_reg_1046__6_ ( .D(n12255), .CP(wclk), .Q(ram[8014]) );
  DFF ram_reg_1046__5_ ( .D(n12254), .CP(wclk), .Q(ram[8013]) );
  DFF ram_reg_1046__4_ ( .D(n12253), .CP(wclk), .Q(ram[8012]) );
  DFF ram_reg_1046__3_ ( .D(n12252), .CP(wclk), .Q(ram[8011]) );
  DFF ram_reg_1046__2_ ( .D(n12251), .CP(wclk), .Q(ram[8010]) );
  DFF ram_reg_1046__1_ ( .D(n12250), .CP(wclk), .Q(ram[8009]) );
  DFF ram_reg_1046__0_ ( .D(n12249), .CP(wclk), .Q(ram[8008]) );
  DFF ram_reg_1050__7_ ( .D(n12224), .CP(wclk), .Q(ram[7983]) );
  DFF ram_reg_1050__6_ ( .D(n12223), .CP(wclk), .Q(ram[7982]) );
  DFF ram_reg_1050__5_ ( .D(n12222), .CP(wclk), .Q(ram[7981]) );
  DFF ram_reg_1050__4_ ( .D(n12221), .CP(wclk), .Q(ram[7980]) );
  DFF ram_reg_1050__3_ ( .D(n12220), .CP(wclk), .Q(ram[7979]) );
  DFF ram_reg_1050__2_ ( .D(n12219), .CP(wclk), .Q(ram[7978]) );
  DFF ram_reg_1050__1_ ( .D(n12218), .CP(wclk), .Q(ram[7977]) );
  DFF ram_reg_1050__0_ ( .D(n12217), .CP(wclk), .Q(ram[7976]) );
  DFF ram_reg_1054__7_ ( .D(n12192), .CP(wclk), .Q(ram[7951]) );
  DFF ram_reg_1054__6_ ( .D(n12191), .CP(wclk), .Q(ram[7950]) );
  DFF ram_reg_1054__5_ ( .D(n12190), .CP(wclk), .Q(ram[7949]) );
  DFF ram_reg_1054__4_ ( .D(n12189), .CP(wclk), .Q(ram[7948]) );
  DFF ram_reg_1054__3_ ( .D(n12188), .CP(wclk), .Q(ram[7947]) );
  DFF ram_reg_1054__2_ ( .D(n12187), .CP(wclk), .Q(ram[7946]) );
  DFF ram_reg_1054__1_ ( .D(n12186), .CP(wclk), .Q(ram[7945]) );
  DFF ram_reg_1054__0_ ( .D(n12185), .CP(wclk), .Q(ram[7944]) );
  DFF ram_reg_1058__7_ ( .D(n12160), .CP(wclk), .Q(ram[7919]) );
  DFF ram_reg_1058__6_ ( .D(n12159), .CP(wclk), .Q(ram[7918]) );
  DFF ram_reg_1058__5_ ( .D(n12158), .CP(wclk), .Q(ram[7917]) );
  DFF ram_reg_1058__4_ ( .D(n12157), .CP(wclk), .Q(ram[7916]) );
  DFF ram_reg_1058__3_ ( .D(n12156), .CP(wclk), .Q(ram[7915]) );
  DFF ram_reg_1058__2_ ( .D(n12155), .CP(wclk), .Q(ram[7914]) );
  DFF ram_reg_1058__1_ ( .D(n12154), .CP(wclk), .Q(ram[7913]) );
  DFF ram_reg_1058__0_ ( .D(n12153), .CP(wclk), .Q(ram[7912]) );
  DFF ram_reg_1062__7_ ( .D(n12128), .CP(wclk), .Q(ram[7887]) );
  DFF ram_reg_1062__6_ ( .D(n12127), .CP(wclk), .Q(ram[7886]) );
  DFF ram_reg_1062__5_ ( .D(n12126), .CP(wclk), .Q(ram[7885]) );
  DFF ram_reg_1062__4_ ( .D(n12125), .CP(wclk), .Q(ram[7884]) );
  DFF ram_reg_1062__3_ ( .D(n12124), .CP(wclk), .Q(ram[7883]) );
  DFF ram_reg_1062__2_ ( .D(n12123), .CP(wclk), .Q(ram[7882]) );
  DFF ram_reg_1062__1_ ( .D(n12122), .CP(wclk), .Q(ram[7881]) );
  DFF ram_reg_1062__0_ ( .D(n12121), .CP(wclk), .Q(ram[7880]) );
  DFF ram_reg_1070__7_ ( .D(n12064), .CP(wclk), .Q(ram[7823]) );
  DFF ram_reg_1070__6_ ( .D(n12063), .CP(wclk), .Q(ram[7822]) );
  DFF ram_reg_1070__5_ ( .D(n12062), .CP(wclk), .Q(ram[7821]) );
  DFF ram_reg_1070__4_ ( .D(n12061), .CP(wclk), .Q(ram[7820]) );
  DFF ram_reg_1070__3_ ( .D(n12060), .CP(wclk), .Q(ram[7819]) );
  DFF ram_reg_1070__2_ ( .D(n12059), .CP(wclk), .Q(ram[7818]) );
  DFF ram_reg_1070__1_ ( .D(n12058), .CP(wclk), .Q(ram[7817]) );
  DFF ram_reg_1070__0_ ( .D(n12057), .CP(wclk), .Q(ram[7816]) );
  DFF ram_reg_1074__7_ ( .D(n12032), .CP(wclk), .Q(ram[7791]) );
  DFF ram_reg_1074__6_ ( .D(n12031), .CP(wclk), .Q(ram[7790]) );
  DFF ram_reg_1074__5_ ( .D(n12030), .CP(wclk), .Q(ram[7789]) );
  DFF ram_reg_1074__4_ ( .D(n12029), .CP(wclk), .Q(ram[7788]) );
  DFF ram_reg_1074__3_ ( .D(n12028), .CP(wclk), .Q(ram[7787]) );
  DFF ram_reg_1074__2_ ( .D(n12027), .CP(wclk), .Q(ram[7786]) );
  DFF ram_reg_1074__1_ ( .D(n12026), .CP(wclk), .Q(ram[7785]) );
  DFF ram_reg_1074__0_ ( .D(n12025), .CP(wclk), .Q(ram[7784]) );
  DFF ram_reg_1078__7_ ( .D(n12000), .CP(wclk), .Q(ram[7759]) );
  DFF ram_reg_1078__6_ ( .D(n11999), .CP(wclk), .Q(ram[7758]) );
  DFF ram_reg_1078__5_ ( .D(n11998), .CP(wclk), .Q(ram[7757]) );
  DFF ram_reg_1078__4_ ( .D(n11997), .CP(wclk), .Q(ram[7756]) );
  DFF ram_reg_1078__3_ ( .D(n11996), .CP(wclk), .Q(ram[7755]) );
  DFF ram_reg_1078__2_ ( .D(n11995), .CP(wclk), .Q(ram[7754]) );
  DFF ram_reg_1078__1_ ( .D(n11994), .CP(wclk), .Q(ram[7753]) );
  DFF ram_reg_1078__0_ ( .D(n11993), .CP(wclk), .Q(ram[7752]) );
  DFF ram_reg_1086__7_ ( .D(n11936), .CP(wclk), .Q(ram[7695]) );
  DFF ram_reg_1086__6_ ( .D(n11935), .CP(wclk), .Q(ram[7694]) );
  DFF ram_reg_1086__5_ ( .D(n11934), .CP(wclk), .Q(ram[7693]) );
  DFF ram_reg_1086__4_ ( .D(n11933), .CP(wclk), .Q(ram[7692]) );
  DFF ram_reg_1086__3_ ( .D(n11932), .CP(wclk), .Q(ram[7691]) );
  DFF ram_reg_1086__2_ ( .D(n11931), .CP(wclk), .Q(ram[7690]) );
  DFF ram_reg_1086__1_ ( .D(n11930), .CP(wclk), .Q(ram[7689]) );
  DFF ram_reg_1086__0_ ( .D(n11929), .CP(wclk), .Q(ram[7688]) );
  DFF ram_reg_1090__7_ ( .D(n11904), .CP(wclk), .Q(ram[7663]) );
  DFF ram_reg_1090__6_ ( .D(n11903), .CP(wclk), .Q(ram[7662]) );
  DFF ram_reg_1090__5_ ( .D(n11902), .CP(wclk), .Q(ram[7661]) );
  DFF ram_reg_1090__4_ ( .D(n11901), .CP(wclk), .Q(ram[7660]) );
  DFF ram_reg_1090__3_ ( .D(n11900), .CP(wclk), .Q(ram[7659]) );
  DFF ram_reg_1090__2_ ( .D(n11899), .CP(wclk), .Q(ram[7658]) );
  DFF ram_reg_1090__1_ ( .D(n11898), .CP(wclk), .Q(ram[7657]) );
  DFF ram_reg_1090__0_ ( .D(n11897), .CP(wclk), .Q(ram[7656]) );
  DFF ram_reg_1094__7_ ( .D(n11872), .CP(wclk), .Q(ram[7631]) );
  DFF ram_reg_1094__6_ ( .D(n11871), .CP(wclk), .Q(ram[7630]) );
  DFF ram_reg_1094__5_ ( .D(n11870), .CP(wclk), .Q(ram[7629]) );
  DFF ram_reg_1094__4_ ( .D(n11869), .CP(wclk), .Q(ram[7628]) );
  DFF ram_reg_1094__3_ ( .D(n11868), .CP(wclk), .Q(ram[7627]) );
  DFF ram_reg_1094__2_ ( .D(n11867), .CP(wclk), .Q(ram[7626]) );
  DFF ram_reg_1094__1_ ( .D(n11866), .CP(wclk), .Q(ram[7625]) );
  DFF ram_reg_1094__0_ ( .D(n11865), .CP(wclk), .Q(ram[7624]) );
  DFF ram_reg_1098__7_ ( .D(n11840), .CP(wclk), .Q(ram[7599]) );
  DFF ram_reg_1098__6_ ( .D(n11839), .CP(wclk), .Q(ram[7598]) );
  DFF ram_reg_1098__5_ ( .D(n11838), .CP(wclk), .Q(ram[7597]) );
  DFF ram_reg_1098__4_ ( .D(n11837), .CP(wclk), .Q(ram[7596]) );
  DFF ram_reg_1098__3_ ( .D(n11836), .CP(wclk), .Q(ram[7595]) );
  DFF ram_reg_1098__2_ ( .D(n11835), .CP(wclk), .Q(ram[7594]) );
  DFF ram_reg_1098__1_ ( .D(n11834), .CP(wclk), .Q(ram[7593]) );
  DFF ram_reg_1098__0_ ( .D(n11833), .CP(wclk), .Q(ram[7592]) );
  DFF ram_reg_1102__7_ ( .D(n11808), .CP(wclk), .Q(ram[7567]) );
  DFF ram_reg_1102__6_ ( .D(n11807), .CP(wclk), .Q(ram[7566]) );
  DFF ram_reg_1102__5_ ( .D(n11806), .CP(wclk), .Q(ram[7565]) );
  DFF ram_reg_1102__4_ ( .D(n11805), .CP(wclk), .Q(ram[7564]) );
  DFF ram_reg_1102__3_ ( .D(n11804), .CP(wclk), .Q(ram[7563]) );
  DFF ram_reg_1102__2_ ( .D(n11803), .CP(wclk), .Q(ram[7562]) );
  DFF ram_reg_1102__1_ ( .D(n11802), .CP(wclk), .Q(ram[7561]) );
  DFF ram_reg_1102__0_ ( .D(n11801), .CP(wclk), .Q(ram[7560]) );
  DFF ram_reg_1106__7_ ( .D(n11776), .CP(wclk), .Q(ram[7535]) );
  DFF ram_reg_1106__6_ ( .D(n11775), .CP(wclk), .Q(ram[7534]) );
  DFF ram_reg_1106__5_ ( .D(n11774), .CP(wclk), .Q(ram[7533]) );
  DFF ram_reg_1106__4_ ( .D(n11773), .CP(wclk), .Q(ram[7532]) );
  DFF ram_reg_1106__3_ ( .D(n11772), .CP(wclk), .Q(ram[7531]) );
  DFF ram_reg_1106__2_ ( .D(n11771), .CP(wclk), .Q(ram[7530]) );
  DFF ram_reg_1106__1_ ( .D(n11770), .CP(wclk), .Q(ram[7529]) );
  DFF ram_reg_1106__0_ ( .D(n11769), .CP(wclk), .Q(ram[7528]) );
  DFF ram_reg_1110__7_ ( .D(n11744), .CP(wclk), .Q(ram[7503]) );
  DFF ram_reg_1110__6_ ( .D(n11743), .CP(wclk), .Q(ram[7502]) );
  DFF ram_reg_1110__5_ ( .D(n11742), .CP(wclk), .Q(ram[7501]) );
  DFF ram_reg_1110__4_ ( .D(n11741), .CP(wclk), .Q(ram[7500]) );
  DFF ram_reg_1110__3_ ( .D(n11740), .CP(wclk), .Q(ram[7499]) );
  DFF ram_reg_1110__2_ ( .D(n11739), .CP(wclk), .Q(ram[7498]) );
  DFF ram_reg_1110__1_ ( .D(n11738), .CP(wclk), .Q(ram[7497]) );
  DFF ram_reg_1110__0_ ( .D(n11737), .CP(wclk), .Q(ram[7496]) );
  DFF ram_reg_1114__7_ ( .D(n11712), .CP(wclk), .Q(ram[7471]) );
  DFF ram_reg_1114__6_ ( .D(n11711), .CP(wclk), .Q(ram[7470]) );
  DFF ram_reg_1114__5_ ( .D(n11710), .CP(wclk), .Q(ram[7469]) );
  DFF ram_reg_1114__4_ ( .D(n11709), .CP(wclk), .Q(ram[7468]) );
  DFF ram_reg_1114__3_ ( .D(n11708), .CP(wclk), .Q(ram[7467]) );
  DFF ram_reg_1114__2_ ( .D(n11707), .CP(wclk), .Q(ram[7466]) );
  DFF ram_reg_1114__1_ ( .D(n11706), .CP(wclk), .Q(ram[7465]) );
  DFF ram_reg_1114__0_ ( .D(n11705), .CP(wclk), .Q(ram[7464]) );
  DFF ram_reg_1118__7_ ( .D(n11680), .CP(wclk), .Q(ram[7439]) );
  DFF ram_reg_1118__6_ ( .D(n11679), .CP(wclk), .Q(ram[7438]) );
  DFF ram_reg_1118__5_ ( .D(n11678), .CP(wclk), .Q(ram[7437]) );
  DFF ram_reg_1118__4_ ( .D(n11677), .CP(wclk), .Q(ram[7436]) );
  DFF ram_reg_1118__3_ ( .D(n11676), .CP(wclk), .Q(ram[7435]) );
  DFF ram_reg_1118__2_ ( .D(n11675), .CP(wclk), .Q(ram[7434]) );
  DFF ram_reg_1118__1_ ( .D(n11674), .CP(wclk), .Q(ram[7433]) );
  DFF ram_reg_1118__0_ ( .D(n11673), .CP(wclk), .Q(ram[7432]) );
  DFF ram_reg_1122__7_ ( .D(n11648), .CP(wclk), .Q(ram[7407]) );
  DFF ram_reg_1122__6_ ( .D(n11647), .CP(wclk), .Q(ram[7406]) );
  DFF ram_reg_1122__5_ ( .D(n11646), .CP(wclk), .Q(ram[7405]) );
  DFF ram_reg_1122__4_ ( .D(n11645), .CP(wclk), .Q(ram[7404]) );
  DFF ram_reg_1122__3_ ( .D(n11644), .CP(wclk), .Q(ram[7403]) );
  DFF ram_reg_1122__2_ ( .D(n11643), .CP(wclk), .Q(ram[7402]) );
  DFF ram_reg_1122__1_ ( .D(n11642), .CP(wclk), .Q(ram[7401]) );
  DFF ram_reg_1122__0_ ( .D(n11641), .CP(wclk), .Q(ram[7400]) );
  DFF ram_reg_1126__7_ ( .D(n11616), .CP(wclk), .Q(ram[7375]) );
  DFF ram_reg_1126__6_ ( .D(n11615), .CP(wclk), .Q(ram[7374]) );
  DFF ram_reg_1126__5_ ( .D(n11614), .CP(wclk), .Q(ram[7373]) );
  DFF ram_reg_1126__4_ ( .D(n11613), .CP(wclk), .Q(ram[7372]) );
  DFF ram_reg_1126__3_ ( .D(n11612), .CP(wclk), .Q(ram[7371]) );
  DFF ram_reg_1126__2_ ( .D(n11611), .CP(wclk), .Q(ram[7370]) );
  DFF ram_reg_1126__1_ ( .D(n11610), .CP(wclk), .Q(ram[7369]) );
  DFF ram_reg_1126__0_ ( .D(n11609), .CP(wclk), .Q(ram[7368]) );
  DFF ram_reg_1130__7_ ( .D(n11584), .CP(wclk), .Q(ram[7343]) );
  DFF ram_reg_1130__6_ ( .D(n11583), .CP(wclk), .Q(ram[7342]) );
  DFF ram_reg_1130__5_ ( .D(n11582), .CP(wclk), .Q(ram[7341]) );
  DFF ram_reg_1130__4_ ( .D(n11581), .CP(wclk), .Q(ram[7340]) );
  DFF ram_reg_1130__3_ ( .D(n11580), .CP(wclk), .Q(ram[7339]) );
  DFF ram_reg_1130__2_ ( .D(n11579), .CP(wclk), .Q(ram[7338]) );
  DFF ram_reg_1130__1_ ( .D(n11578), .CP(wclk), .Q(ram[7337]) );
  DFF ram_reg_1130__0_ ( .D(n11577), .CP(wclk), .Q(ram[7336]) );
  DFF ram_reg_1134__7_ ( .D(n11552), .CP(wclk), .Q(ram[7311]) );
  DFF ram_reg_1134__6_ ( .D(n11551), .CP(wclk), .Q(ram[7310]) );
  DFF ram_reg_1134__5_ ( .D(n11550), .CP(wclk), .Q(ram[7309]) );
  DFF ram_reg_1134__4_ ( .D(n11549), .CP(wclk), .Q(ram[7308]) );
  DFF ram_reg_1134__3_ ( .D(n11548), .CP(wclk), .Q(ram[7307]) );
  DFF ram_reg_1134__2_ ( .D(n11547), .CP(wclk), .Q(ram[7306]) );
  DFF ram_reg_1134__1_ ( .D(n11546), .CP(wclk), .Q(ram[7305]) );
  DFF ram_reg_1134__0_ ( .D(n11545), .CP(wclk), .Q(ram[7304]) );
  DFF ram_reg_1138__7_ ( .D(n11520), .CP(wclk), .Q(ram[7279]) );
  DFF ram_reg_1138__6_ ( .D(n11519), .CP(wclk), .Q(ram[7278]) );
  DFF ram_reg_1138__5_ ( .D(n11518), .CP(wclk), .Q(ram[7277]) );
  DFF ram_reg_1138__4_ ( .D(n11517), .CP(wclk), .Q(ram[7276]) );
  DFF ram_reg_1138__3_ ( .D(n11516), .CP(wclk), .Q(ram[7275]) );
  DFF ram_reg_1138__2_ ( .D(n11515), .CP(wclk), .Q(ram[7274]) );
  DFF ram_reg_1138__1_ ( .D(n11514), .CP(wclk), .Q(ram[7273]) );
  DFF ram_reg_1138__0_ ( .D(n11513), .CP(wclk), .Q(ram[7272]) );
  DFF ram_reg_1142__7_ ( .D(n11488), .CP(wclk), .Q(ram[7247]) );
  DFF ram_reg_1142__6_ ( .D(n11487), .CP(wclk), .Q(ram[7246]) );
  DFF ram_reg_1142__5_ ( .D(n11486), .CP(wclk), .Q(ram[7245]) );
  DFF ram_reg_1142__4_ ( .D(n11485), .CP(wclk), .Q(ram[7244]) );
  DFF ram_reg_1142__3_ ( .D(n11484), .CP(wclk), .Q(ram[7243]) );
  DFF ram_reg_1142__2_ ( .D(n11483), .CP(wclk), .Q(ram[7242]) );
  DFF ram_reg_1142__1_ ( .D(n11482), .CP(wclk), .Q(ram[7241]) );
  DFF ram_reg_1142__0_ ( .D(n11481), .CP(wclk), .Q(ram[7240]) );
  DFF ram_reg_1146__7_ ( .D(n11456), .CP(wclk), .Q(ram[7215]) );
  DFF ram_reg_1146__6_ ( .D(n11455), .CP(wclk), .Q(ram[7214]) );
  DFF ram_reg_1146__5_ ( .D(n11454), .CP(wclk), .Q(ram[7213]) );
  DFF ram_reg_1146__4_ ( .D(n11453), .CP(wclk), .Q(ram[7212]) );
  DFF ram_reg_1146__3_ ( .D(n11452), .CP(wclk), .Q(ram[7211]) );
  DFF ram_reg_1146__2_ ( .D(n11451), .CP(wclk), .Q(ram[7210]) );
  DFF ram_reg_1146__1_ ( .D(n11450), .CP(wclk), .Q(ram[7209]) );
  DFF ram_reg_1146__0_ ( .D(n11449), .CP(wclk), .Q(ram[7208]) );
  DFF ram_reg_1150__7_ ( .D(n11424), .CP(wclk), .Q(ram[7183]) );
  DFF ram_reg_1150__6_ ( .D(n11423), .CP(wclk), .Q(ram[7182]) );
  DFF ram_reg_1150__5_ ( .D(n11422), .CP(wclk), .Q(ram[7181]) );
  DFF ram_reg_1150__4_ ( .D(n11421), .CP(wclk), .Q(ram[7180]) );
  DFF ram_reg_1150__3_ ( .D(n11420), .CP(wclk), .Q(ram[7179]) );
  DFF ram_reg_1150__2_ ( .D(n11419), .CP(wclk), .Q(ram[7178]) );
  DFF ram_reg_1150__1_ ( .D(n11418), .CP(wclk), .Q(ram[7177]) );
  DFF ram_reg_1150__0_ ( .D(n11417), .CP(wclk), .Q(ram[7176]) );
  DFF ram_reg_1154__7_ ( .D(n11392), .CP(wclk), .Q(ram[7151]) );
  DFF ram_reg_1154__6_ ( .D(n11391), .CP(wclk), .Q(ram[7150]) );
  DFF ram_reg_1154__5_ ( .D(n11390), .CP(wclk), .Q(ram[7149]) );
  DFF ram_reg_1154__4_ ( .D(n11389), .CP(wclk), .Q(ram[7148]) );
  DFF ram_reg_1154__3_ ( .D(n11388), .CP(wclk), .Q(ram[7147]) );
  DFF ram_reg_1154__2_ ( .D(n11387), .CP(wclk), .Q(ram[7146]) );
  DFF ram_reg_1154__1_ ( .D(n11386), .CP(wclk), .Q(ram[7145]) );
  DFF ram_reg_1154__0_ ( .D(n11385), .CP(wclk), .Q(ram[7144]) );
  DFF ram_reg_1158__7_ ( .D(n11360), .CP(wclk), .Q(ram[7119]) );
  DFF ram_reg_1158__6_ ( .D(n11359), .CP(wclk), .Q(ram[7118]) );
  DFF ram_reg_1158__5_ ( .D(n11358), .CP(wclk), .Q(ram[7117]) );
  DFF ram_reg_1158__4_ ( .D(n11357), .CP(wclk), .Q(ram[7116]) );
  DFF ram_reg_1158__3_ ( .D(n11356), .CP(wclk), .Q(ram[7115]) );
  DFF ram_reg_1158__2_ ( .D(n11355), .CP(wclk), .Q(ram[7114]) );
  DFF ram_reg_1158__1_ ( .D(n11354), .CP(wclk), .Q(ram[7113]) );
  DFF ram_reg_1158__0_ ( .D(n11353), .CP(wclk), .Q(ram[7112]) );
  DFF ram_reg_1170__7_ ( .D(n11264), .CP(wclk), .Q(ram[7023]) );
  DFF ram_reg_1170__6_ ( .D(n11263), .CP(wclk), .Q(ram[7022]) );
  DFF ram_reg_1170__5_ ( .D(n11262), .CP(wclk), .Q(ram[7021]) );
  DFF ram_reg_1170__4_ ( .D(n11261), .CP(wclk), .Q(ram[7020]) );
  DFF ram_reg_1170__3_ ( .D(n11260), .CP(wclk), .Q(ram[7019]) );
  DFF ram_reg_1170__2_ ( .D(n11259), .CP(wclk), .Q(ram[7018]) );
  DFF ram_reg_1170__1_ ( .D(n11258), .CP(wclk), .Q(ram[7017]) );
  DFF ram_reg_1170__0_ ( .D(n11257), .CP(wclk), .Q(ram[7016]) );
  DFF ram_reg_1174__7_ ( .D(n11232), .CP(wclk), .Q(ram[6991]) );
  DFF ram_reg_1174__6_ ( .D(n11231), .CP(wclk), .Q(ram[6990]) );
  DFF ram_reg_1174__5_ ( .D(n11230), .CP(wclk), .Q(ram[6989]) );
  DFF ram_reg_1174__4_ ( .D(n11229), .CP(wclk), .Q(ram[6988]) );
  DFF ram_reg_1174__3_ ( .D(n11228), .CP(wclk), .Q(ram[6987]) );
  DFF ram_reg_1174__2_ ( .D(n11227), .CP(wclk), .Q(ram[6986]) );
  DFF ram_reg_1174__1_ ( .D(n11226), .CP(wclk), .Q(ram[6985]) );
  DFF ram_reg_1174__0_ ( .D(n11225), .CP(wclk), .Q(ram[6984]) );
  DFF ram_reg_1190__7_ ( .D(n11104), .CP(wclk), .Q(ram[6863]) );
  DFF ram_reg_1190__6_ ( .D(n11103), .CP(wclk), .Q(ram[6862]) );
  DFF ram_reg_1190__5_ ( .D(n11102), .CP(wclk), .Q(ram[6861]) );
  DFF ram_reg_1190__4_ ( .D(n11101), .CP(wclk), .Q(ram[6860]) );
  DFF ram_reg_1190__3_ ( .D(n11100), .CP(wclk), .Q(ram[6859]) );
  DFF ram_reg_1190__2_ ( .D(n11099), .CP(wclk), .Q(ram[6858]) );
  DFF ram_reg_1190__1_ ( .D(n11098), .CP(wclk), .Q(ram[6857]) );
  DFF ram_reg_1190__0_ ( .D(n11097), .CP(wclk), .Q(ram[6856]) );
  DFF ram_reg_1206__7_ ( .D(n10976), .CP(wclk), .Q(ram[6735]) );
  DFF ram_reg_1206__6_ ( .D(n10975), .CP(wclk), .Q(ram[6734]) );
  DFF ram_reg_1206__5_ ( .D(n10974), .CP(wclk), .Q(ram[6733]) );
  DFF ram_reg_1206__4_ ( .D(n10973), .CP(wclk), .Q(ram[6732]) );
  DFF ram_reg_1206__3_ ( .D(n10972), .CP(wclk), .Q(ram[6731]) );
  DFF ram_reg_1206__2_ ( .D(n10971), .CP(wclk), .Q(ram[6730]) );
  DFF ram_reg_1206__1_ ( .D(n10970), .CP(wclk), .Q(ram[6729]) );
  DFF ram_reg_1206__0_ ( .D(n10969), .CP(wclk), .Q(ram[6728]) );
  DFF ram_reg_1218__7_ ( .D(n10880), .CP(wclk), .Q(ram[6639]) );
  DFF ram_reg_1218__6_ ( .D(n10879), .CP(wclk), .Q(ram[6638]) );
  DFF ram_reg_1218__5_ ( .D(n10878), .CP(wclk), .Q(ram[6637]) );
  DFF ram_reg_1218__4_ ( .D(n10877), .CP(wclk), .Q(ram[6636]) );
  DFF ram_reg_1218__3_ ( .D(n10876), .CP(wclk), .Q(ram[6635]) );
  DFF ram_reg_1218__2_ ( .D(n10875), .CP(wclk), .Q(ram[6634]) );
  DFF ram_reg_1218__1_ ( .D(n10874), .CP(wclk), .Q(ram[6633]) );
  DFF ram_reg_1218__0_ ( .D(n10873), .CP(wclk), .Q(ram[6632]) );
  DFF ram_reg_1222__7_ ( .D(n10848), .CP(wclk), .Q(ram[6607]) );
  DFF ram_reg_1222__6_ ( .D(n10847), .CP(wclk), .Q(ram[6606]) );
  DFF ram_reg_1222__5_ ( .D(n10846), .CP(wclk), .Q(ram[6605]) );
  DFF ram_reg_1222__4_ ( .D(n10845), .CP(wclk), .Q(ram[6604]) );
  DFF ram_reg_1222__3_ ( .D(n10844), .CP(wclk), .Q(ram[6603]) );
  DFF ram_reg_1222__2_ ( .D(n10843), .CP(wclk), .Q(ram[6602]) );
  DFF ram_reg_1222__1_ ( .D(n10842), .CP(wclk), .Q(ram[6601]) );
  DFF ram_reg_1222__0_ ( .D(n10841), .CP(wclk), .Q(ram[6600]) );
  DFF ram_reg_1230__7_ ( .D(n10784), .CP(wclk), .Q(ram[6543]) );
  DFF ram_reg_1230__6_ ( .D(n10783), .CP(wclk), .Q(ram[6542]) );
  DFF ram_reg_1230__5_ ( .D(n10782), .CP(wclk), .Q(ram[6541]) );
  DFF ram_reg_1230__4_ ( .D(n10781), .CP(wclk), .Q(ram[6540]) );
  DFF ram_reg_1230__3_ ( .D(n10780), .CP(wclk), .Q(ram[6539]) );
  DFF ram_reg_1230__2_ ( .D(n10779), .CP(wclk), .Q(ram[6538]) );
  DFF ram_reg_1230__1_ ( .D(n10778), .CP(wclk), .Q(ram[6537]) );
  DFF ram_reg_1230__0_ ( .D(n10777), .CP(wclk), .Q(ram[6536]) );
  DFF ram_reg_1234__7_ ( .D(n10752), .CP(wclk), .Q(ram[6511]) );
  DFF ram_reg_1234__6_ ( .D(n10751), .CP(wclk), .Q(ram[6510]) );
  DFF ram_reg_1234__5_ ( .D(n10750), .CP(wclk), .Q(ram[6509]) );
  DFF ram_reg_1234__4_ ( .D(n10749), .CP(wclk), .Q(ram[6508]) );
  DFF ram_reg_1234__3_ ( .D(n10748), .CP(wclk), .Q(ram[6507]) );
  DFF ram_reg_1234__2_ ( .D(n10747), .CP(wclk), .Q(ram[6506]) );
  DFF ram_reg_1234__1_ ( .D(n10746), .CP(wclk), .Q(ram[6505]) );
  DFF ram_reg_1234__0_ ( .D(n10745), .CP(wclk), .Q(ram[6504]) );
  DFF ram_reg_1238__7_ ( .D(n10720), .CP(wclk), .Q(ram[6479]) );
  DFF ram_reg_1238__6_ ( .D(n10719), .CP(wclk), .Q(ram[6478]) );
  DFF ram_reg_1238__5_ ( .D(n10718), .CP(wclk), .Q(ram[6477]) );
  DFF ram_reg_1238__4_ ( .D(n10717), .CP(wclk), .Q(ram[6476]) );
  DFF ram_reg_1238__3_ ( .D(n10716), .CP(wclk), .Q(ram[6475]) );
  DFF ram_reg_1238__2_ ( .D(n10715), .CP(wclk), .Q(ram[6474]) );
  DFF ram_reg_1238__1_ ( .D(n10714), .CP(wclk), .Q(ram[6473]) );
  DFF ram_reg_1238__0_ ( .D(n10713), .CP(wclk), .Q(ram[6472]) );
  DFF ram_reg_1246__7_ ( .D(n10656), .CP(wclk), .Q(ram[6415]) );
  DFF ram_reg_1246__6_ ( .D(n10655), .CP(wclk), .Q(ram[6414]) );
  DFF ram_reg_1246__5_ ( .D(n10654), .CP(wclk), .Q(ram[6413]) );
  DFF ram_reg_1246__4_ ( .D(n10653), .CP(wclk), .Q(ram[6412]) );
  DFF ram_reg_1246__3_ ( .D(n10652), .CP(wclk), .Q(ram[6411]) );
  DFF ram_reg_1246__2_ ( .D(n10651), .CP(wclk), .Q(ram[6410]) );
  DFF ram_reg_1246__1_ ( .D(n10650), .CP(wclk), .Q(ram[6409]) );
  DFF ram_reg_1246__0_ ( .D(n10649), .CP(wclk), .Q(ram[6408]) );
  DFF ram_reg_1250__7_ ( .D(n10624), .CP(wclk), .Q(ram[6383]) );
  DFF ram_reg_1250__6_ ( .D(n10623), .CP(wclk), .Q(ram[6382]) );
  DFF ram_reg_1250__5_ ( .D(n10622), .CP(wclk), .Q(ram[6381]) );
  DFF ram_reg_1250__4_ ( .D(n10621), .CP(wclk), .Q(ram[6380]) );
  DFF ram_reg_1250__3_ ( .D(n10620), .CP(wclk), .Q(ram[6379]) );
  DFF ram_reg_1250__2_ ( .D(n10619), .CP(wclk), .Q(ram[6378]) );
  DFF ram_reg_1250__1_ ( .D(n10618), .CP(wclk), .Q(ram[6377]) );
  DFF ram_reg_1250__0_ ( .D(n10617), .CP(wclk), .Q(ram[6376]) );
  DFF ram_reg_1254__7_ ( .D(n10592), .CP(wclk), .Q(ram[6351]) );
  DFF ram_reg_1254__6_ ( .D(n10591), .CP(wclk), .Q(ram[6350]) );
  DFF ram_reg_1254__5_ ( .D(n10590), .CP(wclk), .Q(ram[6349]) );
  DFF ram_reg_1254__4_ ( .D(n10589), .CP(wclk), .Q(ram[6348]) );
  DFF ram_reg_1254__3_ ( .D(n10588), .CP(wclk), .Q(ram[6347]) );
  DFF ram_reg_1254__2_ ( .D(n10587), .CP(wclk), .Q(ram[6346]) );
  DFF ram_reg_1254__1_ ( .D(n10586), .CP(wclk), .Q(ram[6345]) );
  DFF ram_reg_1254__0_ ( .D(n10585), .CP(wclk), .Q(ram[6344]) );
  DFF ram_reg_1266__7_ ( .D(n10496), .CP(wclk), .Q(ram[6255]) );
  DFF ram_reg_1266__6_ ( .D(n10495), .CP(wclk), .Q(ram[6254]) );
  DFF ram_reg_1266__5_ ( .D(n10494), .CP(wclk), .Q(ram[6253]) );
  DFF ram_reg_1266__4_ ( .D(n10493), .CP(wclk), .Q(ram[6252]) );
  DFF ram_reg_1266__3_ ( .D(n10492), .CP(wclk), .Q(ram[6251]) );
  DFF ram_reg_1266__2_ ( .D(n10491), .CP(wclk), .Q(ram[6250]) );
  DFF ram_reg_1266__1_ ( .D(n10490), .CP(wclk), .Q(ram[6249]) );
  DFF ram_reg_1266__0_ ( .D(n10489), .CP(wclk), .Q(ram[6248]) );
  DFF ram_reg_1270__7_ ( .D(n10464), .CP(wclk), .Q(ram[6223]) );
  DFF ram_reg_1270__6_ ( .D(n10463), .CP(wclk), .Q(ram[6222]) );
  DFF ram_reg_1270__5_ ( .D(n10462), .CP(wclk), .Q(ram[6221]) );
  DFF ram_reg_1270__4_ ( .D(n10461), .CP(wclk), .Q(ram[6220]) );
  DFF ram_reg_1270__3_ ( .D(n10460), .CP(wclk), .Q(ram[6219]) );
  DFF ram_reg_1270__2_ ( .D(n10459), .CP(wclk), .Q(ram[6218]) );
  DFF ram_reg_1270__1_ ( .D(n10458), .CP(wclk), .Q(ram[6217]) );
  DFF ram_reg_1270__0_ ( .D(n10457), .CP(wclk), .Q(ram[6216]) );
  DFF ram_reg_1282__7_ ( .D(n10368), .CP(wclk), .Q(ram[6127]) );
  DFF ram_reg_1282__6_ ( .D(n10367), .CP(wclk), .Q(ram[6126]) );
  DFF ram_reg_1282__5_ ( .D(n10366), .CP(wclk), .Q(ram[6125]) );
  DFF ram_reg_1282__4_ ( .D(n10365), .CP(wclk), .Q(ram[6124]) );
  DFF ram_reg_1282__3_ ( .D(n10364), .CP(wclk), .Q(ram[6123]) );
  DFF ram_reg_1282__2_ ( .D(n10363), .CP(wclk), .Q(ram[6122]) );
  DFF ram_reg_1282__1_ ( .D(n10362), .CP(wclk), .Q(ram[6121]) );
  DFF ram_reg_1282__0_ ( .D(n10361), .CP(wclk), .Q(ram[6120]) );
  DFF ram_reg_1286__7_ ( .D(n10336), .CP(wclk), .Q(ram[6095]) );
  DFF ram_reg_1286__6_ ( .D(n10335), .CP(wclk), .Q(ram[6094]) );
  DFF ram_reg_1286__5_ ( .D(n10334), .CP(wclk), .Q(ram[6093]) );
  DFF ram_reg_1286__4_ ( .D(n10333), .CP(wclk), .Q(ram[6092]) );
  DFF ram_reg_1286__3_ ( .D(n10332), .CP(wclk), .Q(ram[6091]) );
  DFF ram_reg_1286__2_ ( .D(n10331), .CP(wclk), .Q(ram[6090]) );
  DFF ram_reg_1286__1_ ( .D(n10330), .CP(wclk), .Q(ram[6089]) );
  DFF ram_reg_1286__0_ ( .D(n10329), .CP(wclk), .Q(ram[6088]) );
  DFF ram_reg_1298__7_ ( .D(n10240), .CP(wclk), .Q(ram[5999]) );
  DFF ram_reg_1298__6_ ( .D(n10239), .CP(wclk), .Q(ram[5998]) );
  DFF ram_reg_1298__5_ ( .D(n10238), .CP(wclk), .Q(ram[5997]) );
  DFF ram_reg_1298__4_ ( .D(n10237), .CP(wclk), .Q(ram[5996]) );
  DFF ram_reg_1298__3_ ( .D(n10236), .CP(wclk), .Q(ram[5995]) );
  DFF ram_reg_1298__2_ ( .D(n10235), .CP(wclk), .Q(ram[5994]) );
  DFF ram_reg_1298__1_ ( .D(n10234), .CP(wclk), .Q(ram[5993]) );
  DFF ram_reg_1298__0_ ( .D(n10233), .CP(wclk), .Q(ram[5992]) );
  DFF ram_reg_1302__7_ ( .D(n10208), .CP(wclk), .Q(ram[5967]) );
  DFF ram_reg_1302__6_ ( .D(n10207), .CP(wclk), .Q(ram[5966]) );
  DFF ram_reg_1302__5_ ( .D(n10206), .CP(wclk), .Q(ram[5965]) );
  DFF ram_reg_1302__4_ ( .D(n10205), .CP(wclk), .Q(ram[5964]) );
  DFF ram_reg_1302__3_ ( .D(n10204), .CP(wclk), .Q(ram[5963]) );
  DFF ram_reg_1302__2_ ( .D(n10203), .CP(wclk), .Q(ram[5962]) );
  DFF ram_reg_1302__1_ ( .D(n10202), .CP(wclk), .Q(ram[5961]) );
  DFF ram_reg_1302__0_ ( .D(n10201), .CP(wclk), .Q(ram[5960]) );
  DFF ram_reg_1310__7_ ( .D(n10144), .CP(wclk), .Q(ram[5903]) );
  DFF ram_reg_1310__6_ ( .D(n10143), .CP(wclk), .Q(ram[5902]) );
  DFF ram_reg_1310__5_ ( .D(n10142), .CP(wclk), .Q(ram[5901]) );
  DFF ram_reg_1310__4_ ( .D(n10141), .CP(wclk), .Q(ram[5900]) );
  DFF ram_reg_1310__3_ ( .D(n10140), .CP(wclk), .Q(ram[5899]) );
  DFF ram_reg_1310__2_ ( .D(n10139), .CP(wclk), .Q(ram[5898]) );
  DFF ram_reg_1310__1_ ( .D(n10138), .CP(wclk), .Q(ram[5897]) );
  DFF ram_reg_1310__0_ ( .D(n10137), .CP(wclk), .Q(ram[5896]) );
  DFF ram_reg_1314__7_ ( .D(n10112), .CP(wclk), .Q(ram[5871]) );
  DFF ram_reg_1314__6_ ( .D(n10111), .CP(wclk), .Q(ram[5870]) );
  DFF ram_reg_1314__5_ ( .D(n10110), .CP(wclk), .Q(ram[5869]) );
  DFF ram_reg_1314__4_ ( .D(n10109), .CP(wclk), .Q(ram[5868]) );
  DFF ram_reg_1314__3_ ( .D(n10108), .CP(wclk), .Q(ram[5867]) );
  DFF ram_reg_1314__2_ ( .D(n10107), .CP(wclk), .Q(ram[5866]) );
  DFF ram_reg_1314__1_ ( .D(n10106), .CP(wclk), .Q(ram[5865]) );
  DFF ram_reg_1314__0_ ( .D(n10105), .CP(wclk), .Q(ram[5864]) );
  DFF ram_reg_1318__7_ ( .D(n10080), .CP(wclk), .Q(ram[5839]) );
  DFF ram_reg_1318__6_ ( .D(n10079), .CP(wclk), .Q(ram[5838]) );
  DFF ram_reg_1318__5_ ( .D(n10078), .CP(wclk), .Q(ram[5837]) );
  DFF ram_reg_1318__4_ ( .D(n10077), .CP(wclk), .Q(ram[5836]) );
  DFF ram_reg_1318__3_ ( .D(n10076), .CP(wclk), .Q(ram[5835]) );
  DFF ram_reg_1318__2_ ( .D(n10075), .CP(wclk), .Q(ram[5834]) );
  DFF ram_reg_1318__1_ ( .D(n10074), .CP(wclk), .Q(ram[5833]) );
  DFF ram_reg_1318__0_ ( .D(n10073), .CP(wclk), .Q(ram[5832]) );
  DFF ram_reg_1330__7_ ( .D(n9984), .CP(wclk), .Q(ram[5743]) );
  DFF ram_reg_1330__6_ ( .D(n9983), .CP(wclk), .Q(ram[5742]) );
  DFF ram_reg_1330__5_ ( .D(n9982), .CP(wclk), .Q(ram[5741]) );
  DFF ram_reg_1330__4_ ( .D(n9981), .CP(wclk), .Q(ram[5740]) );
  DFF ram_reg_1330__3_ ( .D(n9980), .CP(wclk), .Q(ram[5739]) );
  DFF ram_reg_1330__2_ ( .D(n9979), .CP(wclk), .Q(ram[5738]) );
  DFF ram_reg_1330__1_ ( .D(n9978), .CP(wclk), .Q(ram[5737]) );
  DFF ram_reg_1330__0_ ( .D(n9977), .CP(wclk), .Q(ram[5736]) );
  DFF ram_reg_1334__7_ ( .D(n9952), .CP(wclk), .Q(ram[5711]) );
  DFF ram_reg_1334__6_ ( .D(n9951), .CP(wclk), .Q(ram[5710]) );
  DFF ram_reg_1334__5_ ( .D(n9950), .CP(wclk), .Q(ram[5709]) );
  DFF ram_reg_1334__4_ ( .D(n9949), .CP(wclk), .Q(ram[5708]) );
  DFF ram_reg_1334__3_ ( .D(n9948), .CP(wclk), .Q(ram[5707]) );
  DFF ram_reg_1334__2_ ( .D(n9947), .CP(wclk), .Q(ram[5706]) );
  DFF ram_reg_1334__1_ ( .D(n9946), .CP(wclk), .Q(ram[5705]) );
  DFF ram_reg_1334__0_ ( .D(n9945), .CP(wclk), .Q(ram[5704]) );
  DFF ram_reg_1346__7_ ( .D(n9856), .CP(wclk), .Q(ram[5615]) );
  DFF ram_reg_1346__6_ ( .D(n9855), .CP(wclk), .Q(ram[5614]) );
  DFF ram_reg_1346__5_ ( .D(n9854), .CP(wclk), .Q(ram[5613]) );
  DFF ram_reg_1346__4_ ( .D(n9853), .CP(wclk), .Q(ram[5612]) );
  DFF ram_reg_1346__3_ ( .D(n9852), .CP(wclk), .Q(ram[5611]) );
  DFF ram_reg_1346__2_ ( .D(n9851), .CP(wclk), .Q(ram[5610]) );
  DFF ram_reg_1346__1_ ( .D(n9850), .CP(wclk), .Q(ram[5609]) );
  DFF ram_reg_1346__0_ ( .D(n9849), .CP(wclk), .Q(ram[5608]) );
  DFF ram_reg_1350__7_ ( .D(n9824), .CP(wclk), .Q(ram[5583]) );
  DFF ram_reg_1350__6_ ( .D(n9823), .CP(wclk), .Q(ram[5582]) );
  DFF ram_reg_1350__5_ ( .D(n9822), .CP(wclk), .Q(ram[5581]) );
  DFF ram_reg_1350__4_ ( .D(n9821), .CP(wclk), .Q(ram[5580]) );
  DFF ram_reg_1350__3_ ( .D(n9820), .CP(wclk), .Q(ram[5579]) );
  DFF ram_reg_1350__2_ ( .D(n9819), .CP(wclk), .Q(ram[5578]) );
  DFF ram_reg_1350__1_ ( .D(n9818), .CP(wclk), .Q(ram[5577]) );
  DFF ram_reg_1350__0_ ( .D(n9817), .CP(wclk), .Q(ram[5576]) );
  DFF ram_reg_1354__7_ ( .D(n9792), .CP(wclk), .Q(ram[5551]) );
  DFF ram_reg_1354__6_ ( .D(n9791), .CP(wclk), .Q(ram[5550]) );
  DFF ram_reg_1354__5_ ( .D(n9790), .CP(wclk), .Q(ram[5549]) );
  DFF ram_reg_1354__4_ ( .D(n9789), .CP(wclk), .Q(ram[5548]) );
  DFF ram_reg_1354__3_ ( .D(n9788), .CP(wclk), .Q(ram[5547]) );
  DFF ram_reg_1354__2_ ( .D(n9787), .CP(wclk), .Q(ram[5546]) );
  DFF ram_reg_1354__1_ ( .D(n9786), .CP(wclk), .Q(ram[5545]) );
  DFF ram_reg_1354__0_ ( .D(n9785), .CP(wclk), .Q(ram[5544]) );
  DFF ram_reg_1358__7_ ( .D(n9760), .CP(wclk), .Q(ram[5519]) );
  DFF ram_reg_1358__6_ ( .D(n9759), .CP(wclk), .Q(ram[5518]) );
  DFF ram_reg_1358__5_ ( .D(n9758), .CP(wclk), .Q(ram[5517]) );
  DFF ram_reg_1358__4_ ( .D(n9757), .CP(wclk), .Q(ram[5516]) );
  DFF ram_reg_1358__3_ ( .D(n9756), .CP(wclk), .Q(ram[5515]) );
  DFF ram_reg_1358__2_ ( .D(n9755), .CP(wclk), .Q(ram[5514]) );
  DFF ram_reg_1358__1_ ( .D(n9754), .CP(wclk), .Q(ram[5513]) );
  DFF ram_reg_1358__0_ ( .D(n9753), .CP(wclk), .Q(ram[5512]) );
  DFF ram_reg_1362__7_ ( .D(n9728), .CP(wclk), .Q(ram[5487]) );
  DFF ram_reg_1362__6_ ( .D(n9727), .CP(wclk), .Q(ram[5486]) );
  DFF ram_reg_1362__5_ ( .D(n9726), .CP(wclk), .Q(ram[5485]) );
  DFF ram_reg_1362__4_ ( .D(n9725), .CP(wclk), .Q(ram[5484]) );
  DFF ram_reg_1362__3_ ( .D(n9724), .CP(wclk), .Q(ram[5483]) );
  DFF ram_reg_1362__2_ ( .D(n9723), .CP(wclk), .Q(ram[5482]) );
  DFF ram_reg_1362__1_ ( .D(n9722), .CP(wclk), .Q(ram[5481]) );
  DFF ram_reg_1362__0_ ( .D(n9721), .CP(wclk), .Q(ram[5480]) );
  DFF ram_reg_1366__7_ ( .D(n9696), .CP(wclk), .Q(ram[5455]) );
  DFF ram_reg_1366__6_ ( .D(n9695), .CP(wclk), .Q(ram[5454]) );
  DFF ram_reg_1366__5_ ( .D(n9694), .CP(wclk), .Q(ram[5453]) );
  DFF ram_reg_1366__4_ ( .D(n9693), .CP(wclk), .Q(ram[5452]) );
  DFF ram_reg_1366__3_ ( .D(n9692), .CP(wclk), .Q(ram[5451]) );
  DFF ram_reg_1366__2_ ( .D(n9691), .CP(wclk), .Q(ram[5450]) );
  DFF ram_reg_1366__1_ ( .D(n9690), .CP(wclk), .Q(ram[5449]) );
  DFF ram_reg_1366__0_ ( .D(n9689), .CP(wclk), .Q(ram[5448]) );
  DFF ram_reg_1370__7_ ( .D(n9664), .CP(wclk), .Q(ram[5423]) );
  DFF ram_reg_1370__6_ ( .D(n9663), .CP(wclk), .Q(ram[5422]) );
  DFF ram_reg_1370__5_ ( .D(n9662), .CP(wclk), .Q(ram[5421]) );
  DFF ram_reg_1370__4_ ( .D(n9661), .CP(wclk), .Q(ram[5420]) );
  DFF ram_reg_1370__3_ ( .D(n9660), .CP(wclk), .Q(ram[5419]) );
  DFF ram_reg_1370__2_ ( .D(n9659), .CP(wclk), .Q(ram[5418]) );
  DFF ram_reg_1370__1_ ( .D(n9658), .CP(wclk), .Q(ram[5417]) );
  DFF ram_reg_1370__0_ ( .D(n9657), .CP(wclk), .Q(ram[5416]) );
  DFF ram_reg_1374__7_ ( .D(n9632), .CP(wclk), .Q(ram[5391]) );
  DFF ram_reg_1374__6_ ( .D(n9631), .CP(wclk), .Q(ram[5390]) );
  DFF ram_reg_1374__5_ ( .D(n9630), .CP(wclk), .Q(ram[5389]) );
  DFF ram_reg_1374__4_ ( .D(n9629), .CP(wclk), .Q(ram[5388]) );
  DFF ram_reg_1374__3_ ( .D(n9628), .CP(wclk), .Q(ram[5387]) );
  DFF ram_reg_1374__2_ ( .D(n9627), .CP(wclk), .Q(ram[5386]) );
  DFF ram_reg_1374__1_ ( .D(n9626), .CP(wclk), .Q(ram[5385]) );
  DFF ram_reg_1374__0_ ( .D(n9625), .CP(wclk), .Q(ram[5384]) );
  DFF ram_reg_1378__7_ ( .D(n9600), .CP(wclk), .Q(ram[5359]) );
  DFF ram_reg_1378__6_ ( .D(n9599), .CP(wclk), .Q(ram[5358]) );
  DFF ram_reg_1378__5_ ( .D(n9598), .CP(wclk), .Q(ram[5357]) );
  DFF ram_reg_1378__4_ ( .D(n9597), .CP(wclk), .Q(ram[5356]) );
  DFF ram_reg_1378__3_ ( .D(n9596), .CP(wclk), .Q(ram[5355]) );
  DFF ram_reg_1378__2_ ( .D(n9595), .CP(wclk), .Q(ram[5354]) );
  DFF ram_reg_1378__1_ ( .D(n9594), .CP(wclk), .Q(ram[5353]) );
  DFF ram_reg_1378__0_ ( .D(n9593), .CP(wclk), .Q(ram[5352]) );
  DFF ram_reg_1382__7_ ( .D(n9568), .CP(wclk), .Q(ram[5327]) );
  DFF ram_reg_1382__6_ ( .D(n9567), .CP(wclk), .Q(ram[5326]) );
  DFF ram_reg_1382__5_ ( .D(n9566), .CP(wclk), .Q(ram[5325]) );
  DFF ram_reg_1382__4_ ( .D(n9565), .CP(wclk), .Q(ram[5324]) );
  DFF ram_reg_1382__3_ ( .D(n9564), .CP(wclk), .Q(ram[5323]) );
  DFF ram_reg_1382__2_ ( .D(n9563), .CP(wclk), .Q(ram[5322]) );
  DFF ram_reg_1382__1_ ( .D(n9562), .CP(wclk), .Q(ram[5321]) );
  DFF ram_reg_1382__0_ ( .D(n9561), .CP(wclk), .Q(ram[5320]) );
  DFF ram_reg_1390__7_ ( .D(n9504), .CP(wclk), .Q(ram[5263]) );
  DFF ram_reg_1390__6_ ( .D(n9503), .CP(wclk), .Q(ram[5262]) );
  DFF ram_reg_1390__5_ ( .D(n9502), .CP(wclk), .Q(ram[5261]) );
  DFF ram_reg_1390__4_ ( .D(n9501), .CP(wclk), .Q(ram[5260]) );
  DFF ram_reg_1390__3_ ( .D(n9500), .CP(wclk), .Q(ram[5259]) );
  DFF ram_reg_1390__2_ ( .D(n9499), .CP(wclk), .Q(ram[5258]) );
  DFF ram_reg_1390__1_ ( .D(n9498), .CP(wclk), .Q(ram[5257]) );
  DFF ram_reg_1390__0_ ( .D(n9497), .CP(wclk), .Q(ram[5256]) );
  DFF ram_reg_1394__7_ ( .D(n9472), .CP(wclk), .Q(ram[5231]) );
  DFF ram_reg_1394__6_ ( .D(n9471), .CP(wclk), .Q(ram[5230]) );
  DFF ram_reg_1394__5_ ( .D(n9470), .CP(wclk), .Q(ram[5229]) );
  DFF ram_reg_1394__4_ ( .D(n9469), .CP(wclk), .Q(ram[5228]) );
  DFF ram_reg_1394__3_ ( .D(n9468), .CP(wclk), .Q(ram[5227]) );
  DFF ram_reg_1394__2_ ( .D(n9467), .CP(wclk), .Q(ram[5226]) );
  DFF ram_reg_1394__1_ ( .D(n9466), .CP(wclk), .Q(ram[5225]) );
  DFF ram_reg_1394__0_ ( .D(n9465), .CP(wclk), .Q(ram[5224]) );
  DFF ram_reg_1398__7_ ( .D(n9440), .CP(wclk), .Q(ram[5199]) );
  DFF ram_reg_1398__6_ ( .D(n9439), .CP(wclk), .Q(ram[5198]) );
  DFF ram_reg_1398__5_ ( .D(n9438), .CP(wclk), .Q(ram[5197]) );
  DFF ram_reg_1398__4_ ( .D(n9437), .CP(wclk), .Q(ram[5196]) );
  DFF ram_reg_1398__3_ ( .D(n9436), .CP(wclk), .Q(ram[5195]) );
  DFF ram_reg_1398__2_ ( .D(n9435), .CP(wclk), .Q(ram[5194]) );
  DFF ram_reg_1398__1_ ( .D(n9434), .CP(wclk), .Q(ram[5193]) );
  DFF ram_reg_1398__0_ ( .D(n9433), .CP(wclk), .Q(ram[5192]) );
  DFF ram_reg_1406__7_ ( .D(n9376), .CP(wclk), .Q(ram[5135]) );
  DFF ram_reg_1406__6_ ( .D(n9375), .CP(wclk), .Q(ram[5134]) );
  DFF ram_reg_1406__5_ ( .D(n9374), .CP(wclk), .Q(ram[5133]) );
  DFF ram_reg_1406__4_ ( .D(n9373), .CP(wclk), .Q(ram[5132]) );
  DFF ram_reg_1406__3_ ( .D(n9372), .CP(wclk), .Q(ram[5131]) );
  DFF ram_reg_1406__2_ ( .D(n9371), .CP(wclk), .Q(ram[5130]) );
  DFF ram_reg_1406__1_ ( .D(n9370), .CP(wclk), .Q(ram[5129]) );
  DFF ram_reg_1406__0_ ( .D(n9369), .CP(wclk), .Q(ram[5128]) );
  DFF ram_reg_1414__7_ ( .D(n9312), .CP(wclk), .Q(ram[5071]) );
  DFF ram_reg_1414__6_ ( .D(n9311), .CP(wclk), .Q(ram[5070]) );
  DFF ram_reg_1414__5_ ( .D(n9310), .CP(wclk), .Q(ram[5069]) );
  DFF ram_reg_1414__4_ ( .D(n9309), .CP(wclk), .Q(ram[5068]) );
  DFF ram_reg_1414__3_ ( .D(n9308), .CP(wclk), .Q(ram[5067]) );
  DFF ram_reg_1414__2_ ( .D(n9307), .CP(wclk), .Q(ram[5066]) );
  DFF ram_reg_1414__1_ ( .D(n9306), .CP(wclk), .Q(ram[5065]) );
  DFF ram_reg_1414__0_ ( .D(n9305), .CP(wclk), .Q(ram[5064]) );
  DFF ram_reg_1430__7_ ( .D(n9184), .CP(wclk), .Q(ram[4943]) );
  DFF ram_reg_1430__6_ ( .D(n9183), .CP(wclk), .Q(ram[4942]) );
  DFF ram_reg_1430__5_ ( .D(n9182), .CP(wclk), .Q(ram[4941]) );
  DFF ram_reg_1430__4_ ( .D(n9181), .CP(wclk), .Q(ram[4940]) );
  DFF ram_reg_1430__3_ ( .D(n9180), .CP(wclk), .Q(ram[4939]) );
  DFF ram_reg_1430__2_ ( .D(n9179), .CP(wclk), .Q(ram[4938]) );
  DFF ram_reg_1430__1_ ( .D(n9178), .CP(wclk), .Q(ram[4937]) );
  DFF ram_reg_1430__0_ ( .D(n9177), .CP(wclk), .Q(ram[4936]) );
  DFF ram_reg_1478__7_ ( .D(n8800), .CP(wclk), .Q(ram[4559]) );
  DFF ram_reg_1478__6_ ( .D(n8799), .CP(wclk), .Q(ram[4558]) );
  DFF ram_reg_1478__5_ ( .D(n8798), .CP(wclk), .Q(ram[4557]) );
  DFF ram_reg_1478__4_ ( .D(n8797), .CP(wclk), .Q(ram[4556]) );
  DFF ram_reg_1478__3_ ( .D(n8796), .CP(wclk), .Q(ram[4555]) );
  DFF ram_reg_1478__2_ ( .D(n8795), .CP(wclk), .Q(ram[4554]) );
  DFF ram_reg_1478__1_ ( .D(n8794), .CP(wclk), .Q(ram[4553]) );
  DFF ram_reg_1478__0_ ( .D(n8793), .CP(wclk), .Q(ram[4552]) );
  DFF ram_reg_1490__7_ ( .D(n8704), .CP(wclk), .Q(ram[4463]) );
  DFF ram_reg_1490__6_ ( .D(n8703), .CP(wclk), .Q(ram[4462]) );
  DFF ram_reg_1490__5_ ( .D(n8702), .CP(wclk), .Q(ram[4461]) );
  DFF ram_reg_1490__4_ ( .D(n8701), .CP(wclk), .Q(ram[4460]) );
  DFF ram_reg_1490__3_ ( .D(n8700), .CP(wclk), .Q(ram[4459]) );
  DFF ram_reg_1490__2_ ( .D(n8699), .CP(wclk), .Q(ram[4458]) );
  DFF ram_reg_1490__1_ ( .D(n8698), .CP(wclk), .Q(ram[4457]) );
  DFF ram_reg_1490__0_ ( .D(n8697), .CP(wclk), .Q(ram[4456]) );
  DFF ram_reg_1494__7_ ( .D(n8672), .CP(wclk), .Q(ram[4431]) );
  DFF ram_reg_1494__6_ ( .D(n8671), .CP(wclk), .Q(ram[4430]) );
  DFF ram_reg_1494__5_ ( .D(n8670), .CP(wclk), .Q(ram[4429]) );
  DFF ram_reg_1494__4_ ( .D(n8669), .CP(wclk), .Q(ram[4428]) );
  DFF ram_reg_1494__3_ ( .D(n8668), .CP(wclk), .Q(ram[4427]) );
  DFF ram_reg_1494__2_ ( .D(n8667), .CP(wclk), .Q(ram[4426]) );
  DFF ram_reg_1494__1_ ( .D(n8666), .CP(wclk), .Q(ram[4425]) );
  DFF ram_reg_1494__0_ ( .D(n8665), .CP(wclk), .Q(ram[4424]) );
  DFF ram_reg_1510__7_ ( .D(n8544), .CP(wclk), .Q(ram[4303]) );
  DFF ram_reg_1510__6_ ( .D(n8543), .CP(wclk), .Q(ram[4302]) );
  DFF ram_reg_1510__5_ ( .D(n8542), .CP(wclk), .Q(ram[4301]) );
  DFF ram_reg_1510__4_ ( .D(n8541), .CP(wclk), .Q(ram[4300]) );
  DFF ram_reg_1510__3_ ( .D(n8540), .CP(wclk), .Q(ram[4299]) );
  DFF ram_reg_1510__2_ ( .D(n8539), .CP(wclk), .Q(ram[4298]) );
  DFF ram_reg_1510__1_ ( .D(n8538), .CP(wclk), .Q(ram[4297]) );
  DFF ram_reg_1510__0_ ( .D(n8537), .CP(wclk), .Q(ram[4296]) );
  DFF ram_reg_1526__7_ ( .D(n8416), .CP(wclk), .Q(ram[4175]) );
  DFF ram_reg_1526__6_ ( .D(n8415), .CP(wclk), .Q(ram[4174]) );
  DFF ram_reg_1526__5_ ( .D(n8414), .CP(wclk), .Q(ram[4173]) );
  DFF ram_reg_1526__4_ ( .D(n8413), .CP(wclk), .Q(ram[4172]) );
  DFF ram_reg_1526__3_ ( .D(n8412), .CP(wclk), .Q(ram[4171]) );
  DFF ram_reg_1526__2_ ( .D(n8411), .CP(wclk), .Q(ram[4170]) );
  DFF ram_reg_1526__1_ ( .D(n8410), .CP(wclk), .Q(ram[4169]) );
  DFF ram_reg_1526__0_ ( .D(n8409), .CP(wclk), .Q(ram[4168]) );
  DFF ram_reg_1538__7_ ( .D(n8320), .CP(wclk), .Q(ram[4079]) );
  DFF ram_reg_1538__6_ ( .D(n8319), .CP(wclk), .Q(ram[4078]) );
  DFF ram_reg_1538__5_ ( .D(n8318), .CP(wclk), .Q(ram[4077]) );
  DFF ram_reg_1538__4_ ( .D(n8317), .CP(wclk), .Q(ram[4076]) );
  DFF ram_reg_1538__3_ ( .D(n8316), .CP(wclk), .Q(ram[4075]) );
  DFF ram_reg_1538__2_ ( .D(n8315), .CP(wclk), .Q(ram[4074]) );
  DFF ram_reg_1538__1_ ( .D(n8314), .CP(wclk), .Q(ram[4073]) );
  DFF ram_reg_1538__0_ ( .D(n8313), .CP(wclk), .Q(ram[4072]) );
  DFF ram_reg_1542__7_ ( .D(n8288), .CP(wclk), .Q(ram[4047]) );
  DFF ram_reg_1542__6_ ( .D(n8287), .CP(wclk), .Q(ram[4046]) );
  DFF ram_reg_1542__5_ ( .D(n8286), .CP(wclk), .Q(ram[4045]) );
  DFF ram_reg_1542__4_ ( .D(n8285), .CP(wclk), .Q(ram[4044]) );
  DFF ram_reg_1542__3_ ( .D(n8284), .CP(wclk), .Q(ram[4043]) );
  DFF ram_reg_1542__2_ ( .D(n8283), .CP(wclk), .Q(ram[4042]) );
  DFF ram_reg_1542__1_ ( .D(n8282), .CP(wclk), .Q(ram[4041]) );
  DFF ram_reg_1542__0_ ( .D(n8281), .CP(wclk), .Q(ram[4040]) );
  DFF ram_reg_1546__7_ ( .D(n8256), .CP(wclk), .Q(ram[4015]) );
  DFF ram_reg_1546__6_ ( .D(n8255), .CP(wclk), .Q(ram[4014]) );
  DFF ram_reg_1546__5_ ( .D(n8254), .CP(wclk), .Q(ram[4013]) );
  DFF ram_reg_1546__4_ ( .D(n8253), .CP(wclk), .Q(ram[4012]) );
  DFF ram_reg_1546__3_ ( .D(n8252), .CP(wclk), .Q(ram[4011]) );
  DFF ram_reg_1546__2_ ( .D(n8251), .CP(wclk), .Q(ram[4010]) );
  DFF ram_reg_1546__1_ ( .D(n8250), .CP(wclk), .Q(ram[4009]) );
  DFF ram_reg_1546__0_ ( .D(n8249), .CP(wclk), .Q(ram[4008]) );
  DFF ram_reg_1550__7_ ( .D(n8224), .CP(wclk), .Q(ram[3983]) );
  DFF ram_reg_1550__6_ ( .D(n8223), .CP(wclk), .Q(ram[3982]) );
  DFF ram_reg_1550__5_ ( .D(n8222), .CP(wclk), .Q(ram[3981]) );
  DFF ram_reg_1550__4_ ( .D(n8221), .CP(wclk), .Q(ram[3980]) );
  DFF ram_reg_1550__3_ ( .D(n8220), .CP(wclk), .Q(ram[3979]) );
  DFF ram_reg_1550__2_ ( .D(n8219), .CP(wclk), .Q(ram[3978]) );
  DFF ram_reg_1550__1_ ( .D(n8218), .CP(wclk), .Q(ram[3977]) );
  DFF ram_reg_1550__0_ ( .D(n8217), .CP(wclk), .Q(ram[3976]) );
  DFF ram_reg_1554__7_ ( .D(n8192), .CP(wclk), .Q(ram[3951]) );
  DFF ram_reg_1554__6_ ( .D(n8191), .CP(wclk), .Q(ram[3950]) );
  DFF ram_reg_1554__5_ ( .D(n8190), .CP(wclk), .Q(ram[3949]) );
  DFF ram_reg_1554__4_ ( .D(n8189), .CP(wclk), .Q(ram[3948]) );
  DFF ram_reg_1554__3_ ( .D(n8188), .CP(wclk), .Q(ram[3947]) );
  DFF ram_reg_1554__2_ ( .D(n8187), .CP(wclk), .Q(ram[3946]) );
  DFF ram_reg_1554__1_ ( .D(n8186), .CP(wclk), .Q(ram[3945]) );
  DFF ram_reg_1554__0_ ( .D(n8185), .CP(wclk), .Q(ram[3944]) );
  DFF ram_reg_1558__7_ ( .D(n8160), .CP(wclk), .Q(ram[3919]) );
  DFF ram_reg_1558__6_ ( .D(n8159), .CP(wclk), .Q(ram[3918]) );
  DFF ram_reg_1558__5_ ( .D(n8158), .CP(wclk), .Q(ram[3917]) );
  DFF ram_reg_1558__4_ ( .D(n8157), .CP(wclk), .Q(ram[3916]) );
  DFF ram_reg_1558__3_ ( .D(n8156), .CP(wclk), .Q(ram[3915]) );
  DFF ram_reg_1558__2_ ( .D(n8155), .CP(wclk), .Q(ram[3914]) );
  DFF ram_reg_1558__1_ ( .D(n8154), .CP(wclk), .Q(ram[3913]) );
  DFF ram_reg_1558__0_ ( .D(n8153), .CP(wclk), .Q(ram[3912]) );
  DFF ram_reg_1562__7_ ( .D(n8128), .CP(wclk), .Q(ram[3887]) );
  DFF ram_reg_1562__6_ ( .D(n8127), .CP(wclk), .Q(ram[3886]) );
  DFF ram_reg_1562__5_ ( .D(n8126), .CP(wclk), .Q(ram[3885]) );
  DFF ram_reg_1562__4_ ( .D(n8125), .CP(wclk), .Q(ram[3884]) );
  DFF ram_reg_1562__3_ ( .D(n8124), .CP(wclk), .Q(ram[3883]) );
  DFF ram_reg_1562__2_ ( .D(n8123), .CP(wclk), .Q(ram[3882]) );
  DFF ram_reg_1562__1_ ( .D(n8122), .CP(wclk), .Q(ram[3881]) );
  DFF ram_reg_1562__0_ ( .D(n8121), .CP(wclk), .Q(ram[3880]) );
  DFF ram_reg_1566__7_ ( .D(n8096), .CP(wclk), .Q(ram[3855]) );
  DFF ram_reg_1566__6_ ( .D(n8095), .CP(wclk), .Q(ram[3854]) );
  DFF ram_reg_1566__5_ ( .D(n8094), .CP(wclk), .Q(ram[3853]) );
  DFF ram_reg_1566__4_ ( .D(n8093), .CP(wclk), .Q(ram[3852]) );
  DFF ram_reg_1566__3_ ( .D(n8092), .CP(wclk), .Q(ram[3851]) );
  DFF ram_reg_1566__2_ ( .D(n8091), .CP(wclk), .Q(ram[3850]) );
  DFF ram_reg_1566__1_ ( .D(n8090), .CP(wclk), .Q(ram[3849]) );
  DFF ram_reg_1566__0_ ( .D(n8089), .CP(wclk), .Q(ram[3848]) );
  DFF ram_reg_1570__7_ ( .D(n8064), .CP(wclk), .Q(ram[3823]) );
  DFF ram_reg_1570__6_ ( .D(n8063), .CP(wclk), .Q(ram[3822]) );
  DFF ram_reg_1570__5_ ( .D(n8062), .CP(wclk), .Q(ram[3821]) );
  DFF ram_reg_1570__4_ ( .D(n8061), .CP(wclk), .Q(ram[3820]) );
  DFF ram_reg_1570__3_ ( .D(n8060), .CP(wclk), .Q(ram[3819]) );
  DFF ram_reg_1570__2_ ( .D(n8059), .CP(wclk), .Q(ram[3818]) );
  DFF ram_reg_1570__1_ ( .D(n8058), .CP(wclk), .Q(ram[3817]) );
  DFF ram_reg_1570__0_ ( .D(n8057), .CP(wclk), .Q(ram[3816]) );
  DFF ram_reg_1574__7_ ( .D(n8032), .CP(wclk), .Q(ram[3791]) );
  DFF ram_reg_1574__6_ ( .D(n8031), .CP(wclk), .Q(ram[3790]) );
  DFF ram_reg_1574__5_ ( .D(n8030), .CP(wclk), .Q(ram[3789]) );
  DFF ram_reg_1574__4_ ( .D(n8029), .CP(wclk), .Q(ram[3788]) );
  DFF ram_reg_1574__3_ ( .D(n8028), .CP(wclk), .Q(ram[3787]) );
  DFF ram_reg_1574__2_ ( .D(n8027), .CP(wclk), .Q(ram[3786]) );
  DFF ram_reg_1574__1_ ( .D(n8026), .CP(wclk), .Q(ram[3785]) );
  DFF ram_reg_1574__0_ ( .D(n8025), .CP(wclk), .Q(ram[3784]) );
  DFF ram_reg_1582__7_ ( .D(n7968), .CP(wclk), .Q(ram[3727]) );
  DFF ram_reg_1582__6_ ( .D(n7967), .CP(wclk), .Q(ram[3726]) );
  DFF ram_reg_1582__5_ ( .D(n7966), .CP(wclk), .Q(ram[3725]) );
  DFF ram_reg_1582__4_ ( .D(n7965), .CP(wclk), .Q(ram[3724]) );
  DFF ram_reg_1582__3_ ( .D(n7964), .CP(wclk), .Q(ram[3723]) );
  DFF ram_reg_1582__2_ ( .D(n7963), .CP(wclk), .Q(ram[3722]) );
  DFF ram_reg_1582__1_ ( .D(n7962), .CP(wclk), .Q(ram[3721]) );
  DFF ram_reg_1582__0_ ( .D(n7961), .CP(wclk), .Q(ram[3720]) );
  DFF ram_reg_1586__7_ ( .D(n7936), .CP(wclk), .Q(ram[3695]) );
  DFF ram_reg_1586__6_ ( .D(n7935), .CP(wclk), .Q(ram[3694]) );
  DFF ram_reg_1586__5_ ( .D(n7934), .CP(wclk), .Q(ram[3693]) );
  DFF ram_reg_1586__4_ ( .D(n7933), .CP(wclk), .Q(ram[3692]) );
  DFF ram_reg_1586__3_ ( .D(n7932), .CP(wclk), .Q(ram[3691]) );
  DFF ram_reg_1586__2_ ( .D(n7931), .CP(wclk), .Q(ram[3690]) );
  DFF ram_reg_1586__1_ ( .D(n7930), .CP(wclk), .Q(ram[3689]) );
  DFF ram_reg_1586__0_ ( .D(n7929), .CP(wclk), .Q(ram[3688]) );
  DFF ram_reg_1590__7_ ( .D(n7904), .CP(wclk), .Q(ram[3663]) );
  DFF ram_reg_1590__6_ ( .D(n7903), .CP(wclk), .Q(ram[3662]) );
  DFF ram_reg_1590__5_ ( .D(n7902), .CP(wclk), .Q(ram[3661]) );
  DFF ram_reg_1590__4_ ( .D(n7901), .CP(wclk), .Q(ram[3660]) );
  DFF ram_reg_1590__3_ ( .D(n7900), .CP(wclk), .Q(ram[3659]) );
  DFF ram_reg_1590__2_ ( .D(n7899), .CP(wclk), .Q(ram[3658]) );
  DFF ram_reg_1590__1_ ( .D(n7898), .CP(wclk), .Q(ram[3657]) );
  DFF ram_reg_1590__0_ ( .D(n7897), .CP(wclk), .Q(ram[3656]) );
  DFF ram_reg_1598__7_ ( .D(n7840), .CP(wclk), .Q(ram[3599]) );
  DFF ram_reg_1598__6_ ( .D(n7839), .CP(wclk), .Q(ram[3598]) );
  DFF ram_reg_1598__5_ ( .D(n7838), .CP(wclk), .Q(ram[3597]) );
  DFF ram_reg_1598__4_ ( .D(n7837), .CP(wclk), .Q(ram[3596]) );
  DFF ram_reg_1598__3_ ( .D(n7836), .CP(wclk), .Q(ram[3595]) );
  DFF ram_reg_1598__2_ ( .D(n7835), .CP(wclk), .Q(ram[3594]) );
  DFF ram_reg_1598__1_ ( .D(n7834), .CP(wclk), .Q(ram[3593]) );
  DFF ram_reg_1598__0_ ( .D(n7833), .CP(wclk), .Q(ram[3592]) );
  DFF ram_reg_1602__7_ ( .D(n7808), .CP(wclk), .Q(ram[3567]) );
  DFF ram_reg_1602__6_ ( .D(n7807), .CP(wclk), .Q(ram[3566]) );
  DFF ram_reg_1602__5_ ( .D(n7806), .CP(wclk), .Q(ram[3565]) );
  DFF ram_reg_1602__4_ ( .D(n7805), .CP(wclk), .Q(ram[3564]) );
  DFF ram_reg_1602__3_ ( .D(n7804), .CP(wclk), .Q(ram[3563]) );
  DFF ram_reg_1602__2_ ( .D(n7803), .CP(wclk), .Q(ram[3562]) );
  DFF ram_reg_1602__1_ ( .D(n7802), .CP(wclk), .Q(ram[3561]) );
  DFF ram_reg_1602__0_ ( .D(n7801), .CP(wclk), .Q(ram[3560]) );
  DFF ram_reg_1606__7_ ( .D(n7776), .CP(wclk), .Q(ram[3535]) );
  DFF ram_reg_1606__6_ ( .D(n7775), .CP(wclk), .Q(ram[3534]) );
  DFF ram_reg_1606__5_ ( .D(n7774), .CP(wclk), .Q(ram[3533]) );
  DFF ram_reg_1606__4_ ( .D(n7773), .CP(wclk), .Q(ram[3532]) );
  DFF ram_reg_1606__3_ ( .D(n7772), .CP(wclk), .Q(ram[3531]) );
  DFF ram_reg_1606__2_ ( .D(n7771), .CP(wclk), .Q(ram[3530]) );
  DFF ram_reg_1606__1_ ( .D(n7770), .CP(wclk), .Q(ram[3529]) );
  DFF ram_reg_1606__0_ ( .D(n7769), .CP(wclk), .Q(ram[3528]) );
  DFF ram_reg_1610__7_ ( .D(n7744), .CP(wclk), .Q(ram[3503]) );
  DFF ram_reg_1610__6_ ( .D(n7743), .CP(wclk), .Q(ram[3502]) );
  DFF ram_reg_1610__5_ ( .D(n7742), .CP(wclk), .Q(ram[3501]) );
  DFF ram_reg_1610__4_ ( .D(n7741), .CP(wclk), .Q(ram[3500]) );
  DFF ram_reg_1610__3_ ( .D(n7740), .CP(wclk), .Q(ram[3499]) );
  DFF ram_reg_1610__2_ ( .D(n7739), .CP(wclk), .Q(ram[3498]) );
  DFF ram_reg_1610__1_ ( .D(n7738), .CP(wclk), .Q(ram[3497]) );
  DFF ram_reg_1610__0_ ( .D(n7737), .CP(wclk), .Q(ram[3496]) );
  DFF ram_reg_1614__7_ ( .D(n7712), .CP(wclk), .Q(ram[3471]) );
  DFF ram_reg_1614__6_ ( .D(n7711), .CP(wclk), .Q(ram[3470]) );
  DFF ram_reg_1614__5_ ( .D(n7710), .CP(wclk), .Q(ram[3469]) );
  DFF ram_reg_1614__4_ ( .D(n7709), .CP(wclk), .Q(ram[3468]) );
  DFF ram_reg_1614__3_ ( .D(n7708), .CP(wclk), .Q(ram[3467]) );
  DFF ram_reg_1614__2_ ( .D(n7707), .CP(wclk), .Q(ram[3466]) );
  DFF ram_reg_1614__1_ ( .D(n7706), .CP(wclk), .Q(ram[3465]) );
  DFF ram_reg_1614__0_ ( .D(n7705), .CP(wclk), .Q(ram[3464]) );
  DFF ram_reg_1618__7_ ( .D(n7680), .CP(wclk), .Q(ram[3439]) );
  DFF ram_reg_1618__6_ ( .D(n7679), .CP(wclk), .Q(ram[3438]) );
  DFF ram_reg_1618__5_ ( .D(n7678), .CP(wclk), .Q(ram[3437]) );
  DFF ram_reg_1618__4_ ( .D(n7677), .CP(wclk), .Q(ram[3436]) );
  DFF ram_reg_1618__3_ ( .D(n7676), .CP(wclk), .Q(ram[3435]) );
  DFF ram_reg_1618__2_ ( .D(n7675), .CP(wclk), .Q(ram[3434]) );
  DFF ram_reg_1618__1_ ( .D(n7674), .CP(wclk), .Q(ram[3433]) );
  DFF ram_reg_1618__0_ ( .D(n7673), .CP(wclk), .Q(ram[3432]) );
  DFF ram_reg_1622__7_ ( .D(n7648), .CP(wclk), .Q(ram[3407]) );
  DFF ram_reg_1622__6_ ( .D(n7647), .CP(wclk), .Q(ram[3406]) );
  DFF ram_reg_1622__5_ ( .D(n7646), .CP(wclk), .Q(ram[3405]) );
  DFF ram_reg_1622__4_ ( .D(n7645), .CP(wclk), .Q(ram[3404]) );
  DFF ram_reg_1622__3_ ( .D(n7644), .CP(wclk), .Q(ram[3403]) );
  DFF ram_reg_1622__2_ ( .D(n7643), .CP(wclk), .Q(ram[3402]) );
  DFF ram_reg_1622__1_ ( .D(n7642), .CP(wclk), .Q(ram[3401]) );
  DFF ram_reg_1622__0_ ( .D(n7641), .CP(wclk), .Q(ram[3400]) );
  DFF ram_reg_1626__7_ ( .D(n7616), .CP(wclk), .Q(ram[3375]) );
  DFF ram_reg_1626__6_ ( .D(n7615), .CP(wclk), .Q(ram[3374]) );
  DFF ram_reg_1626__5_ ( .D(n7614), .CP(wclk), .Q(ram[3373]) );
  DFF ram_reg_1626__4_ ( .D(n7613), .CP(wclk), .Q(ram[3372]) );
  DFF ram_reg_1626__3_ ( .D(n7612), .CP(wclk), .Q(ram[3371]) );
  DFF ram_reg_1626__2_ ( .D(n7611), .CP(wclk), .Q(ram[3370]) );
  DFF ram_reg_1626__1_ ( .D(n7610), .CP(wclk), .Q(ram[3369]) );
  DFF ram_reg_1626__0_ ( .D(n7609), .CP(wclk), .Q(ram[3368]) );
  DFF ram_reg_1630__7_ ( .D(n7584), .CP(wclk), .Q(ram[3343]) );
  DFF ram_reg_1630__6_ ( .D(n7583), .CP(wclk), .Q(ram[3342]) );
  DFF ram_reg_1630__5_ ( .D(n7582), .CP(wclk), .Q(ram[3341]) );
  DFF ram_reg_1630__4_ ( .D(n7581), .CP(wclk), .Q(ram[3340]) );
  DFF ram_reg_1630__3_ ( .D(n7580), .CP(wclk), .Q(ram[3339]) );
  DFF ram_reg_1630__2_ ( .D(n7579), .CP(wclk), .Q(ram[3338]) );
  DFF ram_reg_1630__1_ ( .D(n7578), .CP(wclk), .Q(ram[3337]) );
  DFF ram_reg_1630__0_ ( .D(n7577), .CP(wclk), .Q(ram[3336]) );
  DFF ram_reg_1634__7_ ( .D(n7552), .CP(wclk), .Q(ram[3311]) );
  DFF ram_reg_1634__6_ ( .D(n7551), .CP(wclk), .Q(ram[3310]) );
  DFF ram_reg_1634__5_ ( .D(n7550), .CP(wclk), .Q(ram[3309]) );
  DFF ram_reg_1634__4_ ( .D(n7549), .CP(wclk), .Q(ram[3308]) );
  DFF ram_reg_1634__3_ ( .D(n7548), .CP(wclk), .Q(ram[3307]) );
  DFF ram_reg_1634__2_ ( .D(n7547), .CP(wclk), .Q(ram[3306]) );
  DFF ram_reg_1634__1_ ( .D(n7546), .CP(wclk), .Q(ram[3305]) );
  DFF ram_reg_1634__0_ ( .D(n7545), .CP(wclk), .Q(ram[3304]) );
  DFF ram_reg_1638__7_ ( .D(n7520), .CP(wclk), .Q(ram[3279]) );
  DFF ram_reg_1638__6_ ( .D(n7519), .CP(wclk), .Q(ram[3278]) );
  DFF ram_reg_1638__5_ ( .D(n7518), .CP(wclk), .Q(ram[3277]) );
  DFF ram_reg_1638__4_ ( .D(n7517), .CP(wclk), .Q(ram[3276]) );
  DFF ram_reg_1638__3_ ( .D(n7516), .CP(wclk), .Q(ram[3275]) );
  DFF ram_reg_1638__2_ ( .D(n7515), .CP(wclk), .Q(ram[3274]) );
  DFF ram_reg_1638__1_ ( .D(n7514), .CP(wclk), .Q(ram[3273]) );
  DFF ram_reg_1638__0_ ( .D(n7513), .CP(wclk), .Q(ram[3272]) );
  DFF ram_reg_1642__7_ ( .D(n7488), .CP(wclk), .Q(ram[3247]) );
  DFF ram_reg_1642__6_ ( .D(n7487), .CP(wclk), .Q(ram[3246]) );
  DFF ram_reg_1642__5_ ( .D(n7486), .CP(wclk), .Q(ram[3245]) );
  DFF ram_reg_1642__4_ ( .D(n7485), .CP(wclk), .Q(ram[3244]) );
  DFF ram_reg_1642__3_ ( .D(n7484), .CP(wclk), .Q(ram[3243]) );
  DFF ram_reg_1642__2_ ( .D(n7483), .CP(wclk), .Q(ram[3242]) );
  DFF ram_reg_1642__1_ ( .D(n7482), .CP(wclk), .Q(ram[3241]) );
  DFF ram_reg_1642__0_ ( .D(n7481), .CP(wclk), .Q(ram[3240]) );
  DFF ram_reg_1646__7_ ( .D(n7456), .CP(wclk), .Q(ram[3215]) );
  DFF ram_reg_1646__6_ ( .D(n7455), .CP(wclk), .Q(ram[3214]) );
  DFF ram_reg_1646__5_ ( .D(n7454), .CP(wclk), .Q(ram[3213]) );
  DFF ram_reg_1646__4_ ( .D(n7453), .CP(wclk), .Q(ram[3212]) );
  DFF ram_reg_1646__3_ ( .D(n7452), .CP(wclk), .Q(ram[3211]) );
  DFF ram_reg_1646__2_ ( .D(n7451), .CP(wclk), .Q(ram[3210]) );
  DFF ram_reg_1646__1_ ( .D(n7450), .CP(wclk), .Q(ram[3209]) );
  DFF ram_reg_1646__0_ ( .D(n7449), .CP(wclk), .Q(ram[3208]) );
  DFF ram_reg_1650__7_ ( .D(n7424), .CP(wclk), .Q(ram[3183]) );
  DFF ram_reg_1650__6_ ( .D(n7423), .CP(wclk), .Q(ram[3182]) );
  DFF ram_reg_1650__5_ ( .D(n7422), .CP(wclk), .Q(ram[3181]) );
  DFF ram_reg_1650__4_ ( .D(n7421), .CP(wclk), .Q(ram[3180]) );
  DFF ram_reg_1650__3_ ( .D(n7420), .CP(wclk), .Q(ram[3179]) );
  DFF ram_reg_1650__2_ ( .D(n7419), .CP(wclk), .Q(ram[3178]) );
  DFF ram_reg_1650__1_ ( .D(n7418), .CP(wclk), .Q(ram[3177]) );
  DFF ram_reg_1650__0_ ( .D(n7417), .CP(wclk), .Q(ram[3176]) );
  DFF ram_reg_1654__7_ ( .D(n7392), .CP(wclk), .Q(ram[3151]) );
  DFF ram_reg_1654__6_ ( .D(n7391), .CP(wclk), .Q(ram[3150]) );
  DFF ram_reg_1654__5_ ( .D(n7390), .CP(wclk), .Q(ram[3149]) );
  DFF ram_reg_1654__4_ ( .D(n7389), .CP(wclk), .Q(ram[3148]) );
  DFF ram_reg_1654__3_ ( .D(n7388), .CP(wclk), .Q(ram[3147]) );
  DFF ram_reg_1654__2_ ( .D(n7387), .CP(wclk), .Q(ram[3146]) );
  DFF ram_reg_1654__1_ ( .D(n7386), .CP(wclk), .Q(ram[3145]) );
  DFF ram_reg_1654__0_ ( .D(n7385), .CP(wclk), .Q(ram[3144]) );
  DFF ram_reg_1658__7_ ( .D(n7360), .CP(wclk), .Q(ram[3119]) );
  DFF ram_reg_1658__6_ ( .D(n7359), .CP(wclk), .Q(ram[3118]) );
  DFF ram_reg_1658__5_ ( .D(n7358), .CP(wclk), .Q(ram[3117]) );
  DFF ram_reg_1658__4_ ( .D(n7357), .CP(wclk), .Q(ram[3116]) );
  DFF ram_reg_1658__3_ ( .D(n7356), .CP(wclk), .Q(ram[3115]) );
  DFF ram_reg_1658__2_ ( .D(n7355), .CP(wclk), .Q(ram[3114]) );
  DFF ram_reg_1658__1_ ( .D(n7354), .CP(wclk), .Q(ram[3113]) );
  DFF ram_reg_1658__0_ ( .D(n7353), .CP(wclk), .Q(ram[3112]) );
  DFF ram_reg_1662__7_ ( .D(n7328), .CP(wclk), .Q(ram[3087]) );
  DFF ram_reg_1662__6_ ( .D(n7327), .CP(wclk), .Q(ram[3086]) );
  DFF ram_reg_1662__5_ ( .D(n7326), .CP(wclk), .Q(ram[3085]) );
  DFF ram_reg_1662__4_ ( .D(n7325), .CP(wclk), .Q(ram[3084]) );
  DFF ram_reg_1662__3_ ( .D(n7324), .CP(wclk), .Q(ram[3083]) );
  DFF ram_reg_1662__2_ ( .D(n7323), .CP(wclk), .Q(ram[3082]) );
  DFF ram_reg_1662__1_ ( .D(n7322), .CP(wclk), .Q(ram[3081]) );
  DFF ram_reg_1662__0_ ( .D(n7321), .CP(wclk), .Q(ram[3080]) );
  DFF ram_reg_1666__7_ ( .D(n7296), .CP(wclk), .Q(ram[3055]) );
  DFF ram_reg_1666__6_ ( .D(n7295), .CP(wclk), .Q(ram[3054]) );
  DFF ram_reg_1666__5_ ( .D(n7294), .CP(wclk), .Q(ram[3053]) );
  DFF ram_reg_1666__4_ ( .D(n7293), .CP(wclk), .Q(ram[3052]) );
  DFF ram_reg_1666__3_ ( .D(n7292), .CP(wclk), .Q(ram[3051]) );
  DFF ram_reg_1666__2_ ( .D(n7291), .CP(wclk), .Q(ram[3050]) );
  DFF ram_reg_1666__1_ ( .D(n7290), .CP(wclk), .Q(ram[3049]) );
  DFF ram_reg_1666__0_ ( .D(n7289), .CP(wclk), .Q(ram[3048]) );
  DFF ram_reg_1670__7_ ( .D(n7264), .CP(wclk), .Q(ram[3023]) );
  DFF ram_reg_1670__6_ ( .D(n7263), .CP(wclk), .Q(ram[3022]) );
  DFF ram_reg_1670__5_ ( .D(n7262), .CP(wclk), .Q(ram[3021]) );
  DFF ram_reg_1670__4_ ( .D(n7261), .CP(wclk), .Q(ram[3020]) );
  DFF ram_reg_1670__3_ ( .D(n7260), .CP(wclk), .Q(ram[3019]) );
  DFF ram_reg_1670__2_ ( .D(n7259), .CP(wclk), .Q(ram[3018]) );
  DFF ram_reg_1670__1_ ( .D(n7258), .CP(wclk), .Q(ram[3017]) );
  DFF ram_reg_1670__0_ ( .D(n7257), .CP(wclk), .Q(ram[3016]) );
  DFF ram_reg_1682__7_ ( .D(n7168), .CP(wclk), .Q(ram[2927]) );
  DFF ram_reg_1682__6_ ( .D(n7167), .CP(wclk), .Q(ram[2926]) );
  DFF ram_reg_1682__5_ ( .D(n7166), .CP(wclk), .Q(ram[2925]) );
  DFF ram_reg_1682__4_ ( .D(n7165), .CP(wclk), .Q(ram[2924]) );
  DFF ram_reg_1682__3_ ( .D(n7164), .CP(wclk), .Q(ram[2923]) );
  DFF ram_reg_1682__2_ ( .D(n7163), .CP(wclk), .Q(ram[2922]) );
  DFF ram_reg_1682__1_ ( .D(n7162), .CP(wclk), .Q(ram[2921]) );
  DFF ram_reg_1682__0_ ( .D(n7161), .CP(wclk), .Q(ram[2920]) );
  DFF ram_reg_1686__7_ ( .D(n7136), .CP(wclk), .Q(ram[2895]) );
  DFF ram_reg_1686__6_ ( .D(n7135), .CP(wclk), .Q(ram[2894]) );
  DFF ram_reg_1686__5_ ( .D(n7134), .CP(wclk), .Q(ram[2893]) );
  DFF ram_reg_1686__4_ ( .D(n7133), .CP(wclk), .Q(ram[2892]) );
  DFF ram_reg_1686__3_ ( .D(n7132), .CP(wclk), .Q(ram[2891]) );
  DFF ram_reg_1686__2_ ( .D(n7131), .CP(wclk), .Q(ram[2890]) );
  DFF ram_reg_1686__1_ ( .D(n7130), .CP(wclk), .Q(ram[2889]) );
  DFF ram_reg_1686__0_ ( .D(n7129), .CP(wclk), .Q(ram[2888]) );
  DFF ram_reg_1694__7_ ( .D(n7072), .CP(wclk), .Q(ram[2831]) );
  DFF ram_reg_1694__6_ ( .D(n7071), .CP(wclk), .Q(ram[2830]) );
  DFF ram_reg_1694__5_ ( .D(n7070), .CP(wclk), .Q(ram[2829]) );
  DFF ram_reg_1694__4_ ( .D(n7069), .CP(wclk), .Q(ram[2828]) );
  DFF ram_reg_1694__3_ ( .D(n7068), .CP(wclk), .Q(ram[2827]) );
  DFF ram_reg_1694__2_ ( .D(n7067), .CP(wclk), .Q(ram[2826]) );
  DFF ram_reg_1694__1_ ( .D(n7066), .CP(wclk), .Q(ram[2825]) );
  DFF ram_reg_1694__0_ ( .D(n7065), .CP(wclk), .Q(ram[2824]) );
  DFF ram_reg_1702__7_ ( .D(n7008), .CP(wclk), .Q(ram[2767]) );
  DFF ram_reg_1702__6_ ( .D(n7007), .CP(wclk), .Q(ram[2766]) );
  DFF ram_reg_1702__5_ ( .D(n7006), .CP(wclk), .Q(ram[2765]) );
  DFF ram_reg_1702__4_ ( .D(n7005), .CP(wclk), .Q(ram[2764]) );
  DFF ram_reg_1702__3_ ( .D(n7004), .CP(wclk), .Q(ram[2763]) );
  DFF ram_reg_1702__2_ ( .D(n7003), .CP(wclk), .Q(ram[2762]) );
  DFF ram_reg_1702__1_ ( .D(n7002), .CP(wclk), .Q(ram[2761]) );
  DFF ram_reg_1702__0_ ( .D(n7001), .CP(wclk), .Q(ram[2760]) );
  DFF ram_reg_1718__7_ ( .D(n6880), .CP(wclk), .Q(ram[2639]) );
  DFF ram_reg_1718__6_ ( .D(n6879), .CP(wclk), .Q(ram[2638]) );
  DFF ram_reg_1718__5_ ( .D(n6878), .CP(wclk), .Q(ram[2637]) );
  DFF ram_reg_1718__4_ ( .D(n6877), .CP(wclk), .Q(ram[2636]) );
  DFF ram_reg_1718__3_ ( .D(n6876), .CP(wclk), .Q(ram[2635]) );
  DFF ram_reg_1718__2_ ( .D(n6875), .CP(wclk), .Q(ram[2634]) );
  DFF ram_reg_1718__1_ ( .D(n6874), .CP(wclk), .Q(ram[2633]) );
  DFF ram_reg_1718__0_ ( .D(n6873), .CP(wclk), .Q(ram[2632]) );
  DFF ram_reg_1730__7_ ( .D(n6784), .CP(wclk), .Q(ram[2543]) );
  DFF ram_reg_1730__6_ ( .D(n6783), .CP(wclk), .Q(ram[2542]) );
  DFF ram_reg_1730__5_ ( .D(n6782), .CP(wclk), .Q(ram[2541]) );
  DFF ram_reg_1730__4_ ( .D(n6781), .CP(wclk), .Q(ram[2540]) );
  DFF ram_reg_1730__3_ ( .D(n6780), .CP(wclk), .Q(ram[2539]) );
  DFF ram_reg_1730__2_ ( .D(n6779), .CP(wclk), .Q(ram[2538]) );
  DFF ram_reg_1730__1_ ( .D(n6778), .CP(wclk), .Q(ram[2537]) );
  DFF ram_reg_1730__0_ ( .D(n6777), .CP(wclk), .Q(ram[2536]) );
  DFF ram_reg_1734__7_ ( .D(n6752), .CP(wclk), .Q(ram[2511]) );
  DFF ram_reg_1734__6_ ( .D(n6751), .CP(wclk), .Q(ram[2510]) );
  DFF ram_reg_1734__5_ ( .D(n6750), .CP(wclk), .Q(ram[2509]) );
  DFF ram_reg_1734__4_ ( .D(n6749), .CP(wclk), .Q(ram[2508]) );
  DFF ram_reg_1734__3_ ( .D(n6748), .CP(wclk), .Q(ram[2507]) );
  DFF ram_reg_1734__2_ ( .D(n6747), .CP(wclk), .Q(ram[2506]) );
  DFF ram_reg_1734__1_ ( .D(n6746), .CP(wclk), .Q(ram[2505]) );
  DFF ram_reg_1734__0_ ( .D(n6745), .CP(wclk), .Q(ram[2504]) );
  DFF ram_reg_1742__7_ ( .D(n6688), .CP(wclk), .Q(ram[2447]) );
  DFF ram_reg_1742__6_ ( .D(n6687), .CP(wclk), .Q(ram[2446]) );
  DFF ram_reg_1742__5_ ( .D(n6686), .CP(wclk), .Q(ram[2445]) );
  DFF ram_reg_1742__4_ ( .D(n6685), .CP(wclk), .Q(ram[2444]) );
  DFF ram_reg_1742__3_ ( .D(n6684), .CP(wclk), .Q(ram[2443]) );
  DFF ram_reg_1742__2_ ( .D(n6683), .CP(wclk), .Q(ram[2442]) );
  DFF ram_reg_1742__1_ ( .D(n6682), .CP(wclk), .Q(ram[2441]) );
  DFF ram_reg_1742__0_ ( .D(n6681), .CP(wclk), .Q(ram[2440]) );
  DFF ram_reg_1746__7_ ( .D(n6656), .CP(wclk), .Q(ram[2415]) );
  DFF ram_reg_1746__6_ ( .D(n6655), .CP(wclk), .Q(ram[2414]) );
  DFF ram_reg_1746__5_ ( .D(n6654), .CP(wclk), .Q(ram[2413]) );
  DFF ram_reg_1746__4_ ( .D(n6653), .CP(wclk), .Q(ram[2412]) );
  DFF ram_reg_1746__3_ ( .D(n6652), .CP(wclk), .Q(ram[2411]) );
  DFF ram_reg_1746__2_ ( .D(n6651), .CP(wclk), .Q(ram[2410]) );
  DFF ram_reg_1746__1_ ( .D(n6650), .CP(wclk), .Q(ram[2409]) );
  DFF ram_reg_1746__0_ ( .D(n6649), .CP(wclk), .Q(ram[2408]) );
  DFF ram_reg_1750__7_ ( .D(n6624), .CP(wclk), .Q(ram[2383]) );
  DFF ram_reg_1750__6_ ( .D(n6623), .CP(wclk), .Q(ram[2382]) );
  DFF ram_reg_1750__5_ ( .D(n6622), .CP(wclk), .Q(ram[2381]) );
  DFF ram_reg_1750__4_ ( .D(n6621), .CP(wclk), .Q(ram[2380]) );
  DFF ram_reg_1750__3_ ( .D(n6620), .CP(wclk), .Q(ram[2379]) );
  DFF ram_reg_1750__2_ ( .D(n6619), .CP(wclk), .Q(ram[2378]) );
  DFF ram_reg_1750__1_ ( .D(n6618), .CP(wclk), .Q(ram[2377]) );
  DFF ram_reg_1750__0_ ( .D(n6617), .CP(wclk), .Q(ram[2376]) );
  DFF ram_reg_1754__7_ ( .D(n6592), .CP(wclk), .Q(ram[2351]) );
  DFF ram_reg_1754__6_ ( .D(n6591), .CP(wclk), .Q(ram[2350]) );
  DFF ram_reg_1754__5_ ( .D(n6590), .CP(wclk), .Q(ram[2349]) );
  DFF ram_reg_1754__4_ ( .D(n6589), .CP(wclk), .Q(ram[2348]) );
  DFF ram_reg_1754__3_ ( .D(n6588), .CP(wclk), .Q(ram[2347]) );
  DFF ram_reg_1754__2_ ( .D(n6587), .CP(wclk), .Q(ram[2346]) );
  DFF ram_reg_1754__1_ ( .D(n6586), .CP(wclk), .Q(ram[2345]) );
  DFF ram_reg_1754__0_ ( .D(n6585), .CP(wclk), .Q(ram[2344]) );
  DFF ram_reg_1758__7_ ( .D(n6560), .CP(wclk), .Q(ram[2319]) );
  DFF ram_reg_1758__6_ ( .D(n6559), .CP(wclk), .Q(ram[2318]) );
  DFF ram_reg_1758__5_ ( .D(n6558), .CP(wclk), .Q(ram[2317]) );
  DFF ram_reg_1758__4_ ( .D(n6557), .CP(wclk), .Q(ram[2316]) );
  DFF ram_reg_1758__3_ ( .D(n6556), .CP(wclk), .Q(ram[2315]) );
  DFF ram_reg_1758__2_ ( .D(n6555), .CP(wclk), .Q(ram[2314]) );
  DFF ram_reg_1758__1_ ( .D(n6554), .CP(wclk), .Q(ram[2313]) );
  DFF ram_reg_1758__0_ ( .D(n6553), .CP(wclk), .Q(ram[2312]) );
  DFF ram_reg_1762__7_ ( .D(n6528), .CP(wclk), .Q(ram[2287]) );
  DFF ram_reg_1762__6_ ( .D(n6527), .CP(wclk), .Q(ram[2286]) );
  DFF ram_reg_1762__5_ ( .D(n6526), .CP(wclk), .Q(ram[2285]) );
  DFF ram_reg_1762__4_ ( .D(n6525), .CP(wclk), .Q(ram[2284]) );
  DFF ram_reg_1762__3_ ( .D(n6524), .CP(wclk), .Q(ram[2283]) );
  DFF ram_reg_1762__2_ ( .D(n6523), .CP(wclk), .Q(ram[2282]) );
  DFF ram_reg_1762__1_ ( .D(n6522), .CP(wclk), .Q(ram[2281]) );
  DFF ram_reg_1762__0_ ( .D(n6521), .CP(wclk), .Q(ram[2280]) );
  DFF ram_reg_1766__7_ ( .D(n6496), .CP(wclk), .Q(ram[2255]) );
  DFF ram_reg_1766__6_ ( .D(n6495), .CP(wclk), .Q(ram[2254]) );
  DFF ram_reg_1766__5_ ( .D(n6494), .CP(wclk), .Q(ram[2253]) );
  DFF ram_reg_1766__4_ ( .D(n6493), .CP(wclk), .Q(ram[2252]) );
  DFF ram_reg_1766__3_ ( .D(n6492), .CP(wclk), .Q(ram[2251]) );
  DFF ram_reg_1766__2_ ( .D(n6491), .CP(wclk), .Q(ram[2250]) );
  DFF ram_reg_1766__1_ ( .D(n6490), .CP(wclk), .Q(ram[2249]) );
  DFF ram_reg_1766__0_ ( .D(n6489), .CP(wclk), .Q(ram[2248]) );
  DFF ram_reg_1778__7_ ( .D(n6400), .CP(wclk), .Q(ram[2159]) );
  DFF ram_reg_1778__6_ ( .D(n6399), .CP(wclk), .Q(ram[2158]) );
  DFF ram_reg_1778__5_ ( .D(n6398), .CP(wclk), .Q(ram[2157]) );
  DFF ram_reg_1778__4_ ( .D(n6397), .CP(wclk), .Q(ram[2156]) );
  DFF ram_reg_1778__3_ ( .D(n6396), .CP(wclk), .Q(ram[2155]) );
  DFF ram_reg_1778__2_ ( .D(n6395), .CP(wclk), .Q(ram[2154]) );
  DFF ram_reg_1778__1_ ( .D(n6394), .CP(wclk), .Q(ram[2153]) );
  DFF ram_reg_1778__0_ ( .D(n6393), .CP(wclk), .Q(ram[2152]) );
  DFF ram_reg_1782__7_ ( .D(n6368), .CP(wclk), .Q(ram[2127]) );
  DFF ram_reg_1782__6_ ( .D(n6367), .CP(wclk), .Q(ram[2126]) );
  DFF ram_reg_1782__5_ ( .D(n6366), .CP(wclk), .Q(ram[2125]) );
  DFF ram_reg_1782__4_ ( .D(n6365), .CP(wclk), .Q(ram[2124]) );
  DFF ram_reg_1782__3_ ( .D(n6364), .CP(wclk), .Q(ram[2123]) );
  DFF ram_reg_1782__2_ ( .D(n6363), .CP(wclk), .Q(ram[2122]) );
  DFF ram_reg_1782__1_ ( .D(n6362), .CP(wclk), .Q(ram[2121]) );
  DFF ram_reg_1782__0_ ( .D(n6361), .CP(wclk), .Q(ram[2120]) );
  DFF ram_reg_1794__7_ ( .D(n6272), .CP(wclk), .Q(ram[2031]) );
  DFF ram_reg_1794__6_ ( .D(n6271), .CP(wclk), .Q(ram[2030]) );
  DFF ram_reg_1794__5_ ( .D(n6270), .CP(wclk), .Q(ram[2029]) );
  DFF ram_reg_1794__4_ ( .D(n6269), .CP(wclk), .Q(ram[2028]) );
  DFF ram_reg_1794__3_ ( .D(n6268), .CP(wclk), .Q(ram[2027]) );
  DFF ram_reg_1794__2_ ( .D(n6267), .CP(wclk), .Q(ram[2026]) );
  DFF ram_reg_1794__1_ ( .D(n6266), .CP(wclk), .Q(ram[2025]) );
  DFF ram_reg_1794__0_ ( .D(n6265), .CP(wclk), .Q(ram[2024]) );
  DFF ram_reg_1798__7_ ( .D(n6240), .CP(wclk), .Q(ram[1999]) );
  DFF ram_reg_1798__6_ ( .D(n6239), .CP(wclk), .Q(ram[1998]) );
  DFF ram_reg_1798__5_ ( .D(n6238), .CP(wclk), .Q(ram[1997]) );
  DFF ram_reg_1798__4_ ( .D(n6237), .CP(wclk), .Q(ram[1996]) );
  DFF ram_reg_1798__3_ ( .D(n6236), .CP(wclk), .Q(ram[1995]) );
  DFF ram_reg_1798__2_ ( .D(n6235), .CP(wclk), .Q(ram[1994]) );
  DFF ram_reg_1798__1_ ( .D(n6234), .CP(wclk), .Q(ram[1993]) );
  DFF ram_reg_1798__0_ ( .D(n6233), .CP(wclk), .Q(ram[1992]) );
  DFF ram_reg_1802__7_ ( .D(n6208), .CP(wclk), .Q(ram[1967]) );
  DFF ram_reg_1802__6_ ( .D(n6207), .CP(wclk), .Q(ram[1966]) );
  DFF ram_reg_1802__5_ ( .D(n6206), .CP(wclk), .Q(ram[1965]) );
  DFF ram_reg_1802__4_ ( .D(n6205), .CP(wclk), .Q(ram[1964]) );
  DFF ram_reg_1802__3_ ( .D(n6204), .CP(wclk), .Q(ram[1963]) );
  DFF ram_reg_1802__2_ ( .D(n6203), .CP(wclk), .Q(ram[1962]) );
  DFF ram_reg_1802__1_ ( .D(n6202), .CP(wclk), .Q(ram[1961]) );
  DFF ram_reg_1802__0_ ( .D(n6201), .CP(wclk), .Q(ram[1960]) );
  DFF ram_reg_1806__7_ ( .D(n6176), .CP(wclk), .Q(ram[1935]) );
  DFF ram_reg_1806__6_ ( .D(n6175), .CP(wclk), .Q(ram[1934]) );
  DFF ram_reg_1806__5_ ( .D(n6174), .CP(wclk), .Q(ram[1933]) );
  DFF ram_reg_1806__4_ ( .D(n6173), .CP(wclk), .Q(ram[1932]) );
  DFF ram_reg_1806__3_ ( .D(n6172), .CP(wclk), .Q(ram[1931]) );
  DFF ram_reg_1806__2_ ( .D(n6171), .CP(wclk), .Q(ram[1930]) );
  DFF ram_reg_1806__1_ ( .D(n6170), .CP(wclk), .Q(ram[1929]) );
  DFF ram_reg_1806__0_ ( .D(n6169), .CP(wclk), .Q(ram[1928]) );
  DFF ram_reg_1810__7_ ( .D(n6144), .CP(wclk), .Q(ram[1903]) );
  DFF ram_reg_1810__6_ ( .D(n6143), .CP(wclk), .Q(ram[1902]) );
  DFF ram_reg_1810__5_ ( .D(n6142), .CP(wclk), .Q(ram[1901]) );
  DFF ram_reg_1810__4_ ( .D(n6141), .CP(wclk), .Q(ram[1900]) );
  DFF ram_reg_1810__3_ ( .D(n6140), .CP(wclk), .Q(ram[1899]) );
  DFF ram_reg_1810__2_ ( .D(n6139), .CP(wclk), .Q(ram[1898]) );
  DFF ram_reg_1810__1_ ( .D(n6138), .CP(wclk), .Q(ram[1897]) );
  DFF ram_reg_1810__0_ ( .D(n6137), .CP(wclk), .Q(ram[1896]) );
  DFF ram_reg_1814__7_ ( .D(n6112), .CP(wclk), .Q(ram[1871]) );
  DFF ram_reg_1814__6_ ( .D(n6111), .CP(wclk), .Q(ram[1870]) );
  DFF ram_reg_1814__5_ ( .D(n6110), .CP(wclk), .Q(ram[1869]) );
  DFF ram_reg_1814__4_ ( .D(n6109), .CP(wclk), .Q(ram[1868]) );
  DFF ram_reg_1814__3_ ( .D(n6108), .CP(wclk), .Q(ram[1867]) );
  DFF ram_reg_1814__2_ ( .D(n6107), .CP(wclk), .Q(ram[1866]) );
  DFF ram_reg_1814__1_ ( .D(n6106), .CP(wclk), .Q(ram[1865]) );
  DFF ram_reg_1814__0_ ( .D(n6105), .CP(wclk), .Q(ram[1864]) );
  DFF ram_reg_1818__7_ ( .D(n6080), .CP(wclk), .Q(ram[1839]) );
  DFF ram_reg_1818__6_ ( .D(n6079), .CP(wclk), .Q(ram[1838]) );
  DFF ram_reg_1818__5_ ( .D(n6078), .CP(wclk), .Q(ram[1837]) );
  DFF ram_reg_1818__4_ ( .D(n6077), .CP(wclk), .Q(ram[1836]) );
  DFF ram_reg_1818__3_ ( .D(n6076), .CP(wclk), .Q(ram[1835]) );
  DFF ram_reg_1818__2_ ( .D(n6075), .CP(wclk), .Q(ram[1834]) );
  DFF ram_reg_1818__1_ ( .D(n6074), .CP(wclk), .Q(ram[1833]) );
  DFF ram_reg_1818__0_ ( .D(n6073), .CP(wclk), .Q(ram[1832]) );
  DFF ram_reg_1822__7_ ( .D(n6048), .CP(wclk), .Q(ram[1807]) );
  DFF ram_reg_1822__6_ ( .D(n6047), .CP(wclk), .Q(ram[1806]) );
  DFF ram_reg_1822__5_ ( .D(n6046), .CP(wclk), .Q(ram[1805]) );
  DFF ram_reg_1822__4_ ( .D(n6045), .CP(wclk), .Q(ram[1804]) );
  DFF ram_reg_1822__3_ ( .D(n6044), .CP(wclk), .Q(ram[1803]) );
  DFF ram_reg_1822__2_ ( .D(n6043), .CP(wclk), .Q(ram[1802]) );
  DFF ram_reg_1822__1_ ( .D(n6042), .CP(wclk), .Q(ram[1801]) );
  DFF ram_reg_1822__0_ ( .D(n6041), .CP(wclk), .Q(ram[1800]) );
  DFF ram_reg_1826__7_ ( .D(n6016), .CP(wclk), .Q(ram[1775]) );
  DFF ram_reg_1826__6_ ( .D(n6015), .CP(wclk), .Q(ram[1774]) );
  DFF ram_reg_1826__5_ ( .D(n6014), .CP(wclk), .Q(ram[1773]) );
  DFF ram_reg_1826__4_ ( .D(n6013), .CP(wclk), .Q(ram[1772]) );
  DFF ram_reg_1826__3_ ( .D(n6012), .CP(wclk), .Q(ram[1771]) );
  DFF ram_reg_1826__2_ ( .D(n6011), .CP(wclk), .Q(ram[1770]) );
  DFF ram_reg_1826__1_ ( .D(n6010), .CP(wclk), .Q(ram[1769]) );
  DFF ram_reg_1826__0_ ( .D(n6009), .CP(wclk), .Q(ram[1768]) );
  DFF ram_reg_1830__7_ ( .D(n5984), .CP(wclk), .Q(ram[1743]) );
  DFF ram_reg_1830__6_ ( .D(n5983), .CP(wclk), .Q(ram[1742]) );
  DFF ram_reg_1830__5_ ( .D(n5982), .CP(wclk), .Q(ram[1741]) );
  DFF ram_reg_1830__4_ ( .D(n5981), .CP(wclk), .Q(ram[1740]) );
  DFF ram_reg_1830__3_ ( .D(n5980), .CP(wclk), .Q(ram[1739]) );
  DFF ram_reg_1830__2_ ( .D(n5979), .CP(wclk), .Q(ram[1738]) );
  DFF ram_reg_1830__1_ ( .D(n5978), .CP(wclk), .Q(ram[1737]) );
  DFF ram_reg_1830__0_ ( .D(n5977), .CP(wclk), .Q(ram[1736]) );
  DFF ram_reg_1838__7_ ( .D(n5920), .CP(wclk), .Q(ram[1679]) );
  DFF ram_reg_1838__6_ ( .D(n5919), .CP(wclk), .Q(ram[1678]) );
  DFF ram_reg_1838__5_ ( .D(n5918), .CP(wclk), .Q(ram[1677]) );
  DFF ram_reg_1838__4_ ( .D(n5917), .CP(wclk), .Q(ram[1676]) );
  DFF ram_reg_1838__3_ ( .D(n5916), .CP(wclk), .Q(ram[1675]) );
  DFF ram_reg_1838__2_ ( .D(n5915), .CP(wclk), .Q(ram[1674]) );
  DFF ram_reg_1838__1_ ( .D(n5914), .CP(wclk), .Q(ram[1673]) );
  DFF ram_reg_1838__0_ ( .D(n5913), .CP(wclk), .Q(ram[1672]) );
  DFF ram_reg_1842__7_ ( .D(n5888), .CP(wclk), .Q(ram[1647]) );
  DFF ram_reg_1842__6_ ( .D(n5887), .CP(wclk), .Q(ram[1646]) );
  DFF ram_reg_1842__5_ ( .D(n5886), .CP(wclk), .Q(ram[1645]) );
  DFF ram_reg_1842__4_ ( .D(n5885), .CP(wclk), .Q(ram[1644]) );
  DFF ram_reg_1842__3_ ( .D(n5884), .CP(wclk), .Q(ram[1643]) );
  DFF ram_reg_1842__2_ ( .D(n5883), .CP(wclk), .Q(ram[1642]) );
  DFF ram_reg_1842__1_ ( .D(n5882), .CP(wclk), .Q(ram[1641]) );
  DFF ram_reg_1842__0_ ( .D(n5881), .CP(wclk), .Q(ram[1640]) );
  DFF ram_reg_1846__7_ ( .D(n5856), .CP(wclk), .Q(ram[1615]) );
  DFF ram_reg_1846__6_ ( .D(n5855), .CP(wclk), .Q(ram[1614]) );
  DFF ram_reg_1846__5_ ( .D(n5854), .CP(wclk), .Q(ram[1613]) );
  DFF ram_reg_1846__4_ ( .D(n5853), .CP(wclk), .Q(ram[1612]) );
  DFF ram_reg_1846__3_ ( .D(n5852), .CP(wclk), .Q(ram[1611]) );
  DFF ram_reg_1846__2_ ( .D(n5851), .CP(wclk), .Q(ram[1610]) );
  DFF ram_reg_1846__1_ ( .D(n5850), .CP(wclk), .Q(ram[1609]) );
  DFF ram_reg_1846__0_ ( .D(n5849), .CP(wclk), .Q(ram[1608]) );
  DFF ram_reg_1858__7_ ( .D(n5760), .CP(wclk), .Q(ram[1519]) );
  DFF ram_reg_1858__6_ ( .D(n5759), .CP(wclk), .Q(ram[1518]) );
  DFF ram_reg_1858__5_ ( .D(n5758), .CP(wclk), .Q(ram[1517]) );
  DFF ram_reg_1858__4_ ( .D(n5757), .CP(wclk), .Q(ram[1516]) );
  DFF ram_reg_1858__3_ ( .D(n5756), .CP(wclk), .Q(ram[1515]) );
  DFF ram_reg_1858__2_ ( .D(n5755), .CP(wclk), .Q(ram[1514]) );
  DFF ram_reg_1858__1_ ( .D(n5754), .CP(wclk), .Q(ram[1513]) );
  DFF ram_reg_1858__0_ ( .D(n5753), .CP(wclk), .Q(ram[1512]) );
  DFF ram_reg_1862__7_ ( .D(n5728), .CP(wclk), .Q(ram[1487]) );
  DFF ram_reg_1862__6_ ( .D(n5727), .CP(wclk), .Q(ram[1486]) );
  DFF ram_reg_1862__5_ ( .D(n5726), .CP(wclk), .Q(ram[1485]) );
  DFF ram_reg_1862__4_ ( .D(n5725), .CP(wclk), .Q(ram[1484]) );
  DFF ram_reg_1862__3_ ( .D(n5724), .CP(wclk), .Q(ram[1483]) );
  DFF ram_reg_1862__2_ ( .D(n5723), .CP(wclk), .Q(ram[1482]) );
  DFF ram_reg_1862__1_ ( .D(n5722), .CP(wclk), .Q(ram[1481]) );
  DFF ram_reg_1862__0_ ( .D(n5721), .CP(wclk), .Q(ram[1480]) );
  DFF ram_reg_1866__7_ ( .D(n5696), .CP(wclk), .Q(ram[1455]) );
  DFF ram_reg_1866__6_ ( .D(n5695), .CP(wclk), .Q(ram[1454]) );
  DFF ram_reg_1866__5_ ( .D(n5694), .CP(wclk), .Q(ram[1453]) );
  DFF ram_reg_1866__4_ ( .D(n5693), .CP(wclk), .Q(ram[1452]) );
  DFF ram_reg_1866__3_ ( .D(n5692), .CP(wclk), .Q(ram[1451]) );
  DFF ram_reg_1866__2_ ( .D(n5691), .CP(wclk), .Q(ram[1450]) );
  DFF ram_reg_1866__1_ ( .D(n5690), .CP(wclk), .Q(ram[1449]) );
  DFF ram_reg_1866__0_ ( .D(n5689), .CP(wclk), .Q(ram[1448]) );
  DFF ram_reg_1870__7_ ( .D(n5664), .CP(wclk), .Q(ram[1423]) );
  DFF ram_reg_1870__6_ ( .D(n5663), .CP(wclk), .Q(ram[1422]) );
  DFF ram_reg_1870__5_ ( .D(n5662), .CP(wclk), .Q(ram[1421]) );
  DFF ram_reg_1870__4_ ( .D(n5661), .CP(wclk), .Q(ram[1420]) );
  DFF ram_reg_1870__3_ ( .D(n5660), .CP(wclk), .Q(ram[1419]) );
  DFF ram_reg_1870__2_ ( .D(n5659), .CP(wclk), .Q(ram[1418]) );
  DFF ram_reg_1870__1_ ( .D(n5658), .CP(wclk), .Q(ram[1417]) );
  DFF ram_reg_1870__0_ ( .D(n5657), .CP(wclk), .Q(ram[1416]) );
  DFF ram_reg_1874__7_ ( .D(n5632), .CP(wclk), .Q(ram[1391]) );
  DFF ram_reg_1874__6_ ( .D(n5631), .CP(wclk), .Q(ram[1390]) );
  DFF ram_reg_1874__5_ ( .D(n5630), .CP(wclk), .Q(ram[1389]) );
  DFF ram_reg_1874__4_ ( .D(n5629), .CP(wclk), .Q(ram[1388]) );
  DFF ram_reg_1874__3_ ( .D(n5628), .CP(wclk), .Q(ram[1387]) );
  DFF ram_reg_1874__2_ ( .D(n5627), .CP(wclk), .Q(ram[1386]) );
  DFF ram_reg_1874__1_ ( .D(n5626), .CP(wclk), .Q(ram[1385]) );
  DFF ram_reg_1874__0_ ( .D(n5625), .CP(wclk), .Q(ram[1384]) );
  DFF ram_reg_1878__7_ ( .D(n5600), .CP(wclk), .Q(ram[1359]) );
  DFF ram_reg_1878__6_ ( .D(n5599), .CP(wclk), .Q(ram[1358]) );
  DFF ram_reg_1878__5_ ( .D(n5598), .CP(wclk), .Q(ram[1357]) );
  DFF ram_reg_1878__4_ ( .D(n5597), .CP(wclk), .Q(ram[1356]) );
  DFF ram_reg_1878__3_ ( .D(n5596), .CP(wclk), .Q(ram[1355]) );
  DFF ram_reg_1878__2_ ( .D(n5595), .CP(wclk), .Q(ram[1354]) );
  DFF ram_reg_1878__1_ ( .D(n5594), .CP(wclk), .Q(ram[1353]) );
  DFF ram_reg_1878__0_ ( .D(n5593), .CP(wclk), .Q(ram[1352]) );
  DFF ram_reg_1882__7_ ( .D(n5568), .CP(wclk), .Q(ram[1327]) );
  DFF ram_reg_1882__6_ ( .D(n5567), .CP(wclk), .Q(ram[1326]) );
  DFF ram_reg_1882__5_ ( .D(n5566), .CP(wclk), .Q(ram[1325]) );
  DFF ram_reg_1882__4_ ( .D(n5565), .CP(wclk), .Q(ram[1324]) );
  DFF ram_reg_1882__3_ ( .D(n5564), .CP(wclk), .Q(ram[1323]) );
  DFF ram_reg_1882__2_ ( .D(n5563), .CP(wclk), .Q(ram[1322]) );
  DFF ram_reg_1882__1_ ( .D(n5562), .CP(wclk), .Q(ram[1321]) );
  DFF ram_reg_1882__0_ ( .D(n5561), .CP(wclk), .Q(ram[1320]) );
  DFF ram_reg_1886__7_ ( .D(n5536), .CP(wclk), .Q(ram[1295]) );
  DFF ram_reg_1886__6_ ( .D(n5535), .CP(wclk), .Q(ram[1294]) );
  DFF ram_reg_1886__5_ ( .D(n5534), .CP(wclk), .Q(ram[1293]) );
  DFF ram_reg_1886__4_ ( .D(n5533), .CP(wclk), .Q(ram[1292]) );
  DFF ram_reg_1886__3_ ( .D(n5532), .CP(wclk), .Q(ram[1291]) );
  DFF ram_reg_1886__2_ ( .D(n5531), .CP(wclk), .Q(ram[1290]) );
  DFF ram_reg_1886__1_ ( .D(n5530), .CP(wclk), .Q(ram[1289]) );
  DFF ram_reg_1886__0_ ( .D(n5529), .CP(wclk), .Q(ram[1288]) );
  DFF ram_reg_1890__7_ ( .D(n5504), .CP(wclk), .Q(ram[1263]) );
  DFF ram_reg_1890__6_ ( .D(n5503), .CP(wclk), .Q(ram[1262]) );
  DFF ram_reg_1890__5_ ( .D(n5502), .CP(wclk), .Q(ram[1261]) );
  DFF ram_reg_1890__4_ ( .D(n5501), .CP(wclk), .Q(ram[1260]) );
  DFF ram_reg_1890__3_ ( .D(n5500), .CP(wclk), .Q(ram[1259]) );
  DFF ram_reg_1890__2_ ( .D(n5499), .CP(wclk), .Q(ram[1258]) );
  DFF ram_reg_1890__1_ ( .D(n5498), .CP(wclk), .Q(ram[1257]) );
  DFF ram_reg_1890__0_ ( .D(n5497), .CP(wclk), .Q(ram[1256]) );
  DFF ram_reg_1894__7_ ( .D(n5472), .CP(wclk), .Q(ram[1231]) );
  DFF ram_reg_1894__6_ ( .D(n5471), .CP(wclk), .Q(ram[1230]) );
  DFF ram_reg_1894__5_ ( .D(n5470), .CP(wclk), .Q(ram[1229]) );
  DFF ram_reg_1894__4_ ( .D(n5469), .CP(wclk), .Q(ram[1228]) );
  DFF ram_reg_1894__3_ ( .D(n5468), .CP(wclk), .Q(ram[1227]) );
  DFF ram_reg_1894__2_ ( .D(n5467), .CP(wclk), .Q(ram[1226]) );
  DFF ram_reg_1894__1_ ( .D(n5466), .CP(wclk), .Q(ram[1225]) );
  DFF ram_reg_1894__0_ ( .D(n5465), .CP(wclk), .Q(ram[1224]) );
  DFF ram_reg_1898__7_ ( .D(n5440), .CP(wclk), .Q(ram[1199]) );
  DFF ram_reg_1898__6_ ( .D(n5439), .CP(wclk), .Q(ram[1198]) );
  DFF ram_reg_1898__5_ ( .D(n5438), .CP(wclk), .Q(ram[1197]) );
  DFF ram_reg_1898__4_ ( .D(n5437), .CP(wclk), .Q(ram[1196]) );
  DFF ram_reg_1898__3_ ( .D(n5436), .CP(wclk), .Q(ram[1195]) );
  DFF ram_reg_1898__2_ ( .D(n5435), .CP(wclk), .Q(ram[1194]) );
  DFF ram_reg_1898__1_ ( .D(n5434), .CP(wclk), .Q(ram[1193]) );
  DFF ram_reg_1898__0_ ( .D(n5433), .CP(wclk), .Q(ram[1192]) );
  DFF ram_reg_1902__7_ ( .D(n5408), .CP(wclk), .Q(ram[1167]) );
  DFF ram_reg_1902__6_ ( .D(n5407), .CP(wclk), .Q(ram[1166]) );
  DFF ram_reg_1902__5_ ( .D(n5406), .CP(wclk), .Q(ram[1165]) );
  DFF ram_reg_1902__4_ ( .D(n5405), .CP(wclk), .Q(ram[1164]) );
  DFF ram_reg_1902__3_ ( .D(n5404), .CP(wclk), .Q(ram[1163]) );
  DFF ram_reg_1902__2_ ( .D(n5403), .CP(wclk), .Q(ram[1162]) );
  DFF ram_reg_1902__1_ ( .D(n5402), .CP(wclk), .Q(ram[1161]) );
  DFF ram_reg_1902__0_ ( .D(n5401), .CP(wclk), .Q(ram[1160]) );
  DFF ram_reg_1906__7_ ( .D(n5376), .CP(wclk), .Q(ram[1135]) );
  DFF ram_reg_1906__6_ ( .D(n5375), .CP(wclk), .Q(ram[1134]) );
  DFF ram_reg_1906__5_ ( .D(n5374), .CP(wclk), .Q(ram[1133]) );
  DFF ram_reg_1906__4_ ( .D(n5373), .CP(wclk), .Q(ram[1132]) );
  DFF ram_reg_1906__3_ ( .D(n5372), .CP(wclk), .Q(ram[1131]) );
  DFF ram_reg_1906__2_ ( .D(n5371), .CP(wclk), .Q(ram[1130]) );
  DFF ram_reg_1906__1_ ( .D(n5370), .CP(wclk), .Q(ram[1129]) );
  DFF ram_reg_1906__0_ ( .D(n5369), .CP(wclk), .Q(ram[1128]) );
  DFF ram_reg_1910__7_ ( .D(n5344), .CP(wclk), .Q(ram[1103]) );
  DFF ram_reg_1910__6_ ( .D(n5343), .CP(wclk), .Q(ram[1102]) );
  DFF ram_reg_1910__5_ ( .D(n5342), .CP(wclk), .Q(ram[1101]) );
  DFF ram_reg_1910__4_ ( .D(n5341), .CP(wclk), .Q(ram[1100]) );
  DFF ram_reg_1910__3_ ( .D(n5340), .CP(wclk), .Q(ram[1099]) );
  DFF ram_reg_1910__2_ ( .D(n5339), .CP(wclk), .Q(ram[1098]) );
  DFF ram_reg_1910__1_ ( .D(n5338), .CP(wclk), .Q(ram[1097]) );
  DFF ram_reg_1910__0_ ( .D(n5337), .CP(wclk), .Q(ram[1096]) );
  DFF ram_reg_1914__7_ ( .D(n5312), .CP(wclk), .Q(ram[1071]) );
  DFF ram_reg_1914__6_ ( .D(n5311), .CP(wclk), .Q(ram[1070]) );
  DFF ram_reg_1914__5_ ( .D(n5310), .CP(wclk), .Q(ram[1069]) );
  DFF ram_reg_1914__4_ ( .D(n5309), .CP(wclk), .Q(ram[1068]) );
  DFF ram_reg_1914__3_ ( .D(n5308), .CP(wclk), .Q(ram[1067]) );
  DFF ram_reg_1914__2_ ( .D(n5307), .CP(wclk), .Q(ram[1066]) );
  DFF ram_reg_1914__1_ ( .D(n5306), .CP(wclk), .Q(ram[1065]) );
  DFF ram_reg_1914__0_ ( .D(n5305), .CP(wclk), .Q(ram[1064]) );
  DFF ram_reg_1918__7_ ( .D(n5280), .CP(wclk), .Q(ram[1039]) );
  DFF ram_reg_1918__6_ ( .D(n5279), .CP(wclk), .Q(ram[1038]) );
  DFF ram_reg_1918__5_ ( .D(n5278), .CP(wclk), .Q(ram[1037]) );
  DFF ram_reg_1918__4_ ( .D(n5277), .CP(wclk), .Q(ram[1036]) );
  DFF ram_reg_1918__3_ ( .D(n5276), .CP(wclk), .Q(ram[1035]) );
  DFF ram_reg_1918__2_ ( .D(n5275), .CP(wclk), .Q(ram[1034]) );
  DFF ram_reg_1918__1_ ( .D(n5274), .CP(wclk), .Q(ram[1033]) );
  DFF ram_reg_1918__0_ ( .D(n5273), .CP(wclk), .Q(ram[1032]) );
  DFF ram_reg_1922__7_ ( .D(n5248), .CP(wclk), .Q(ram[1007]) );
  DFF ram_reg_1922__6_ ( .D(n5247), .CP(wclk), .Q(ram[1006]) );
  DFF ram_reg_1922__5_ ( .D(n5246), .CP(wclk), .Q(ram[1005]) );
  DFF ram_reg_1922__4_ ( .D(n5245), .CP(wclk), .Q(ram[1004]) );
  DFF ram_reg_1922__3_ ( .D(n5244), .CP(wclk), .Q(ram[1003]) );
  DFF ram_reg_1922__2_ ( .D(n5243), .CP(wclk), .Q(ram[1002]) );
  DFF ram_reg_1922__1_ ( .D(n5242), .CP(wclk), .Q(ram[1001]) );
  DFF ram_reg_1922__0_ ( .D(n5241), .CP(wclk), .Q(ram[1000]) );
  DFF ram_reg_1926__7_ ( .D(n5216), .CP(wclk), .Q(ram[975]) );
  DFF ram_reg_1926__6_ ( .D(n5215), .CP(wclk), .Q(ram[974]) );
  DFF ram_reg_1926__5_ ( .D(n5214), .CP(wclk), .Q(ram[973]) );
  DFF ram_reg_1926__4_ ( .D(n5213), .CP(wclk), .Q(ram[972]) );
  DFF ram_reg_1926__3_ ( .D(n5212), .CP(wclk), .Q(ram[971]) );
  DFF ram_reg_1926__2_ ( .D(n5211), .CP(wclk), .Q(ram[970]) );
  DFF ram_reg_1926__1_ ( .D(n5210), .CP(wclk), .Q(ram[969]) );
  DFF ram_reg_1926__0_ ( .D(n5209), .CP(wclk), .Q(ram[968]) );
  DFF ram_reg_1938__7_ ( .D(n5120), .CP(wclk), .Q(ram[879]) );
  DFF ram_reg_1938__6_ ( .D(n5119), .CP(wclk), .Q(ram[878]) );
  DFF ram_reg_1938__5_ ( .D(n5118), .CP(wclk), .Q(ram[877]) );
  DFF ram_reg_1938__4_ ( .D(n5117), .CP(wclk), .Q(ram[876]) );
  DFF ram_reg_1938__3_ ( .D(n5116), .CP(wclk), .Q(ram[875]) );
  DFF ram_reg_1938__2_ ( .D(n5115), .CP(wclk), .Q(ram[874]) );
  DFF ram_reg_1938__1_ ( .D(n5114), .CP(wclk), .Q(ram[873]) );
  DFF ram_reg_1938__0_ ( .D(n5113), .CP(wclk), .Q(ram[872]) );
  DFF ram_reg_1942__7_ ( .D(n5088), .CP(wclk), .Q(ram[847]) );
  DFF ram_reg_1942__6_ ( .D(n5087), .CP(wclk), .Q(ram[846]) );
  DFF ram_reg_1942__5_ ( .D(n5086), .CP(wclk), .Q(ram[845]) );
  DFF ram_reg_1942__4_ ( .D(n5085), .CP(wclk), .Q(ram[844]) );
  DFF ram_reg_1942__3_ ( .D(n5084), .CP(wclk), .Q(ram[843]) );
  DFF ram_reg_1942__2_ ( .D(n5083), .CP(wclk), .Q(ram[842]) );
  DFF ram_reg_1942__1_ ( .D(n5082), .CP(wclk), .Q(ram[841]) );
  DFF ram_reg_1942__0_ ( .D(n5081), .CP(wclk), .Q(ram[840]) );
  DFF ram_reg_1958__7_ ( .D(n4960), .CP(wclk), .Q(ram[719]) );
  DFF ram_reg_1958__6_ ( .D(n4959), .CP(wclk), .Q(ram[718]) );
  DFF ram_reg_1958__5_ ( .D(n4958), .CP(wclk), .Q(ram[717]) );
  DFF ram_reg_1958__4_ ( .D(n4957), .CP(wclk), .Q(ram[716]) );
  DFF ram_reg_1958__3_ ( .D(n4956), .CP(wclk), .Q(ram[715]) );
  DFF ram_reg_1958__2_ ( .D(n4955), .CP(wclk), .Q(ram[714]) );
  DFF ram_reg_1958__1_ ( .D(n4954), .CP(wclk), .Q(ram[713]) );
  DFF ram_reg_1958__0_ ( .D(n4953), .CP(wclk), .Q(ram[712]) );
  DFF ram_reg_1974__7_ ( .D(n4832), .CP(wclk), .Q(ram[591]) );
  DFF ram_reg_1974__6_ ( .D(n4831), .CP(wclk), .Q(ram[590]) );
  DFF ram_reg_1974__5_ ( .D(n4830), .CP(wclk), .Q(ram[589]) );
  DFF ram_reg_1974__4_ ( .D(n4829), .CP(wclk), .Q(ram[588]) );
  DFF ram_reg_1974__3_ ( .D(n4828), .CP(wclk), .Q(ram[587]) );
  DFF ram_reg_1974__2_ ( .D(n4827), .CP(wclk), .Q(ram[586]) );
  DFF ram_reg_1974__1_ ( .D(n4826), .CP(wclk), .Q(ram[585]) );
  DFF ram_reg_1974__0_ ( .D(n4825), .CP(wclk), .Q(ram[584]) );
  DFF ram_reg_1986__7_ ( .D(n4736), .CP(wclk), .Q(ram[495]) );
  DFF ram_reg_1986__6_ ( .D(n4735), .CP(wclk), .Q(ram[494]) );
  DFF ram_reg_1986__5_ ( .D(n4734), .CP(wclk), .Q(ram[493]) );
  DFF ram_reg_1986__4_ ( .D(n4733), .CP(wclk), .Q(ram[492]) );
  DFF ram_reg_1986__3_ ( .D(n4732), .CP(wclk), .Q(ram[491]) );
  DFF ram_reg_1986__2_ ( .D(n4731), .CP(wclk), .Q(ram[490]) );
  DFF ram_reg_1986__1_ ( .D(n4730), .CP(wclk), .Q(ram[489]) );
  DFF ram_reg_1986__0_ ( .D(n4729), .CP(wclk), .Q(ram[488]) );
  DFF ram_reg_1990__7_ ( .D(n4704), .CP(wclk), .Q(ram[463]) );
  DFF ram_reg_1990__6_ ( .D(n4703), .CP(wclk), .Q(ram[462]) );
  DFF ram_reg_1990__5_ ( .D(n4702), .CP(wclk), .Q(ram[461]) );
  DFF ram_reg_1990__4_ ( .D(n4701), .CP(wclk), .Q(ram[460]) );
  DFF ram_reg_1990__3_ ( .D(n4700), .CP(wclk), .Q(ram[459]) );
  DFF ram_reg_1990__2_ ( .D(n4699), .CP(wclk), .Q(ram[458]) );
  DFF ram_reg_1990__1_ ( .D(n4698), .CP(wclk), .Q(ram[457]) );
  DFF ram_reg_1990__0_ ( .D(n4697), .CP(wclk), .Q(ram[456]) );
  DFF ram_reg_2002__7_ ( .D(n4608), .CP(wclk), .Q(ram[367]) );
  DFF ram_reg_2002__6_ ( .D(n4607), .CP(wclk), .Q(ram[366]) );
  DFF ram_reg_2002__5_ ( .D(n4606), .CP(wclk), .Q(ram[365]) );
  DFF ram_reg_2002__4_ ( .D(n4605), .CP(wclk), .Q(ram[364]) );
  DFF ram_reg_2002__3_ ( .D(n4604), .CP(wclk), .Q(ram[363]) );
  DFF ram_reg_2002__2_ ( .D(n4603), .CP(wclk), .Q(ram[362]) );
  DFF ram_reg_2002__1_ ( .D(n4602), .CP(wclk), .Q(ram[361]) );
  DFF ram_reg_2002__0_ ( .D(n4601), .CP(wclk), .Q(ram[360]) );
  DFF ram_reg_2006__7_ ( .D(n4576), .CP(wclk), .Q(ram[335]) );
  DFF ram_reg_2006__6_ ( .D(n4575), .CP(wclk), .Q(ram[334]) );
  DFF ram_reg_2006__5_ ( .D(n4574), .CP(wclk), .Q(ram[333]) );
  DFF ram_reg_2006__4_ ( .D(n4573), .CP(wclk), .Q(ram[332]) );
  DFF ram_reg_2006__3_ ( .D(n4572), .CP(wclk), .Q(ram[331]) );
  DFF ram_reg_2006__2_ ( .D(n4571), .CP(wclk), .Q(ram[330]) );
  DFF ram_reg_2006__1_ ( .D(n4570), .CP(wclk), .Q(ram[329]) );
  DFF ram_reg_2006__0_ ( .D(n4569), .CP(wclk), .Q(ram[328]) );
  DFF ram_reg_2014__7_ ( .D(n4512), .CP(wclk), .Q(ram[271]) );
  DFF ram_reg_2014__6_ ( .D(n4511), .CP(wclk), .Q(ram[270]) );
  DFF ram_reg_2014__5_ ( .D(n4510), .CP(wclk), .Q(ram[269]) );
  DFF ram_reg_2014__4_ ( .D(n4509), .CP(wclk), .Q(ram[268]) );
  DFF ram_reg_2014__3_ ( .D(n4508), .CP(wclk), .Q(ram[267]) );
  DFF ram_reg_2014__2_ ( .D(n4507), .CP(wclk), .Q(ram[266]) );
  DFF ram_reg_2014__1_ ( .D(n4506), .CP(wclk), .Q(ram[265]) );
  DFF ram_reg_2014__0_ ( .D(n4505), .CP(wclk), .Q(ram[264]) );
  DFF ram_reg_2018__7_ ( .D(n4480), .CP(wclk), .Q(ram[239]) );
  DFF ram_reg_2018__6_ ( .D(n4479), .CP(wclk), .Q(ram[238]) );
  DFF ram_reg_2018__5_ ( .D(n4478), .CP(wclk), .Q(ram[237]) );
  DFF ram_reg_2018__4_ ( .D(n4477), .CP(wclk), .Q(ram[236]) );
  DFF ram_reg_2018__3_ ( .D(n4476), .CP(wclk), .Q(ram[235]) );
  DFF ram_reg_2018__2_ ( .D(n4475), .CP(wclk), .Q(ram[234]) );
  DFF ram_reg_2018__1_ ( .D(n4474), .CP(wclk), .Q(ram[233]) );
  DFF ram_reg_2018__0_ ( .D(n4473), .CP(wclk), .Q(ram[232]) );
  DFF ram_reg_2022__7_ ( .D(n4448), .CP(wclk), .Q(ram[207]) );
  DFF ram_reg_2022__6_ ( .D(n4447), .CP(wclk), .Q(ram[206]) );
  DFF ram_reg_2022__5_ ( .D(n4446), .CP(wclk), .Q(ram[205]) );
  DFF ram_reg_2022__4_ ( .D(n4445), .CP(wclk), .Q(ram[204]) );
  DFF ram_reg_2022__3_ ( .D(n4444), .CP(wclk), .Q(ram[203]) );
  DFF ram_reg_2022__2_ ( .D(n4443), .CP(wclk), .Q(ram[202]) );
  DFF ram_reg_2022__1_ ( .D(n4442), .CP(wclk), .Q(ram[201]) );
  DFF ram_reg_2022__0_ ( .D(n4441), .CP(wclk), .Q(ram[200]) );
  DFF ram_reg_2038__7_ ( .D(n4320), .CP(wclk), .Q(ram[79]) );
  DFF ram_reg_2038__6_ ( .D(n4319), .CP(wclk), .Q(ram[78]) );
  DFF ram_reg_2038__5_ ( .D(n4318), .CP(wclk), .Q(ram[77]) );
  DFF ram_reg_2038__4_ ( .D(n4317), .CP(wclk), .Q(ram[76]) );
  DFF ram_reg_2038__3_ ( .D(n4316), .CP(wclk), .Q(ram[75]) );
  DFF ram_reg_2038__2_ ( .D(n4315), .CP(wclk), .Q(ram[74]) );
  DFF ram_reg_2038__1_ ( .D(n4314), .CP(wclk), .Q(ram[73]) );
  DFF ram_reg_2038__0_ ( .D(n4313), .CP(wclk), .Q(ram[72]) );
  DFF ram_reg_1__7_ ( .D(n20616), .CP(wclk), .Q(ram[16375]) );
  DFF ram_reg_1__6_ ( .D(n20615), .CP(wclk), .Q(ram[16374]) );
  DFF ram_reg_1__5_ ( .D(n20614), .CP(wclk), .Q(ram[16373]) );
  DFF ram_reg_1__4_ ( .D(n20613), .CP(wclk), .Q(ram[16372]) );
  DFF ram_reg_1__3_ ( .D(n20612), .CP(wclk), .Q(ram[16371]) );
  DFF ram_reg_1__2_ ( .D(n20611), .CP(wclk), .Q(ram[16370]) );
  DFF ram_reg_1__1_ ( .D(n20610), .CP(wclk), .Q(ram[16369]) );
  DFF ram_reg_1__0_ ( .D(n20609), .CP(wclk), .Q(ram[16368]) );
  DFF ram_reg_5__7_ ( .D(n20584), .CP(wclk), .Q(ram[16343]) );
  DFF ram_reg_5__6_ ( .D(n20583), .CP(wclk), .Q(ram[16342]) );
  DFF ram_reg_5__5_ ( .D(n20582), .CP(wclk), .Q(ram[16341]) );
  DFF ram_reg_5__4_ ( .D(n20581), .CP(wclk), .Q(ram[16340]) );
  DFF ram_reg_5__3_ ( .D(n20580), .CP(wclk), .Q(ram[16339]) );
  DFF ram_reg_5__2_ ( .D(n20579), .CP(wclk), .Q(ram[16338]) );
  DFF ram_reg_5__1_ ( .D(n20578), .CP(wclk), .Q(ram[16337]) );
  DFF ram_reg_5__0_ ( .D(n20577), .CP(wclk), .Q(ram[16336]) );
  DFF ram_reg_13__7_ ( .D(n20520), .CP(wclk), .Q(ram[16279]) );
  DFF ram_reg_13__6_ ( .D(n20519), .CP(wclk), .Q(ram[16278]) );
  DFF ram_reg_13__5_ ( .D(n20518), .CP(wclk), .Q(ram[16277]) );
  DFF ram_reg_13__4_ ( .D(n20517), .CP(wclk), .Q(ram[16276]) );
  DFF ram_reg_13__3_ ( .D(n20516), .CP(wclk), .Q(ram[16275]) );
  DFF ram_reg_13__2_ ( .D(n20515), .CP(wclk), .Q(ram[16274]) );
  DFF ram_reg_13__1_ ( .D(n20514), .CP(wclk), .Q(ram[16273]) );
  DFF ram_reg_13__0_ ( .D(n20513), .CP(wclk), .Q(ram[16272]) );
  DFF ram_reg_17__7_ ( .D(n20488), .CP(wclk), .Q(ram[16247]) );
  DFF ram_reg_17__6_ ( .D(n20487), .CP(wclk), .Q(ram[16246]) );
  DFF ram_reg_17__5_ ( .D(n20486), .CP(wclk), .Q(ram[16245]) );
  DFF ram_reg_17__4_ ( .D(n20485), .CP(wclk), .Q(ram[16244]) );
  DFF ram_reg_17__3_ ( .D(n20484), .CP(wclk), .Q(ram[16243]) );
  DFF ram_reg_17__2_ ( .D(n20483), .CP(wclk), .Q(ram[16242]) );
  DFF ram_reg_17__1_ ( .D(n20482), .CP(wclk), .Q(ram[16241]) );
  DFF ram_reg_17__0_ ( .D(n20481), .CP(wclk), .Q(ram[16240]) );
  DFF ram_reg_21__7_ ( .D(n20456), .CP(wclk), .Q(ram[16215]) );
  DFF ram_reg_21__6_ ( .D(n20455), .CP(wclk), .Q(ram[16214]) );
  DFF ram_reg_21__5_ ( .D(n20454), .CP(wclk), .Q(ram[16213]) );
  DFF ram_reg_21__4_ ( .D(n20453), .CP(wclk), .Q(ram[16212]) );
  DFF ram_reg_21__3_ ( .D(n20452), .CP(wclk), .Q(ram[16211]) );
  DFF ram_reg_21__2_ ( .D(n20451), .CP(wclk), .Q(ram[16210]) );
  DFF ram_reg_21__1_ ( .D(n20450), .CP(wclk), .Q(ram[16209]) );
  DFF ram_reg_21__0_ ( .D(n20449), .CP(wclk), .Q(ram[16208]) );
  DFF ram_reg_25__7_ ( .D(n20424), .CP(wclk), .Q(ram[16183]) );
  DFF ram_reg_25__6_ ( .D(n20423), .CP(wclk), .Q(ram[16182]) );
  DFF ram_reg_25__5_ ( .D(n20422), .CP(wclk), .Q(ram[16181]) );
  DFF ram_reg_25__4_ ( .D(n20421), .CP(wclk), .Q(ram[16180]) );
  DFF ram_reg_25__3_ ( .D(n20420), .CP(wclk), .Q(ram[16179]) );
  DFF ram_reg_25__2_ ( .D(n20419), .CP(wclk), .Q(ram[16178]) );
  DFF ram_reg_25__1_ ( .D(n20418), .CP(wclk), .Q(ram[16177]) );
  DFF ram_reg_25__0_ ( .D(n20417), .CP(wclk), .Q(ram[16176]) );
  DFF ram_reg_29__7_ ( .D(n20392), .CP(wclk), .Q(ram[16151]) );
  DFF ram_reg_29__6_ ( .D(n20391), .CP(wclk), .Q(ram[16150]) );
  DFF ram_reg_29__5_ ( .D(n20390), .CP(wclk), .Q(ram[16149]) );
  DFF ram_reg_29__4_ ( .D(n20389), .CP(wclk), .Q(ram[16148]) );
  DFF ram_reg_29__3_ ( .D(n20388), .CP(wclk), .Q(ram[16147]) );
  DFF ram_reg_29__2_ ( .D(n20387), .CP(wclk), .Q(ram[16146]) );
  DFF ram_reg_29__1_ ( .D(n20386), .CP(wclk), .Q(ram[16145]) );
  DFF ram_reg_29__0_ ( .D(n20385), .CP(wclk), .Q(ram[16144]) );
  DFF ram_reg_33__7_ ( .D(n20360), .CP(wclk), .Q(ram[16119]) );
  DFF ram_reg_33__6_ ( .D(n20359), .CP(wclk), .Q(ram[16118]) );
  DFF ram_reg_33__5_ ( .D(n20358), .CP(wclk), .Q(ram[16117]) );
  DFF ram_reg_33__4_ ( .D(n20357), .CP(wclk), .Q(ram[16116]) );
  DFF ram_reg_33__3_ ( .D(n20356), .CP(wclk), .Q(ram[16115]) );
  DFF ram_reg_33__2_ ( .D(n20355), .CP(wclk), .Q(ram[16114]) );
  DFF ram_reg_33__1_ ( .D(n20354), .CP(wclk), .Q(ram[16113]) );
  DFF ram_reg_33__0_ ( .D(n20353), .CP(wclk), .Q(ram[16112]) );
  DFF ram_reg_37__7_ ( .D(n20328), .CP(wclk), .Q(ram[16087]) );
  DFF ram_reg_37__6_ ( .D(n20327), .CP(wclk), .Q(ram[16086]) );
  DFF ram_reg_37__5_ ( .D(n20326), .CP(wclk), .Q(ram[16085]) );
  DFF ram_reg_37__4_ ( .D(n20325), .CP(wclk), .Q(ram[16084]) );
  DFF ram_reg_37__3_ ( .D(n20324), .CP(wclk), .Q(ram[16083]) );
  DFF ram_reg_37__2_ ( .D(n20323), .CP(wclk), .Q(ram[16082]) );
  DFF ram_reg_37__1_ ( .D(n20322), .CP(wclk), .Q(ram[16081]) );
  DFF ram_reg_37__0_ ( .D(n20321), .CP(wclk), .Q(ram[16080]) );
  DFF ram_reg_49__7_ ( .D(n20232), .CP(wclk), .Q(ram[15991]) );
  DFF ram_reg_49__6_ ( .D(n20231), .CP(wclk), .Q(ram[15990]) );
  DFF ram_reg_49__5_ ( .D(n20230), .CP(wclk), .Q(ram[15989]) );
  DFF ram_reg_49__4_ ( .D(n20229), .CP(wclk), .Q(ram[15988]) );
  DFF ram_reg_49__3_ ( .D(n20228), .CP(wclk), .Q(ram[15987]) );
  DFF ram_reg_49__2_ ( .D(n20227), .CP(wclk), .Q(ram[15986]) );
  DFF ram_reg_49__1_ ( .D(n20226), .CP(wclk), .Q(ram[15985]) );
  DFF ram_reg_49__0_ ( .D(n20225), .CP(wclk), .Q(ram[15984]) );
  DFF ram_reg_53__7_ ( .D(n20200), .CP(wclk), .Q(ram[15959]) );
  DFF ram_reg_53__6_ ( .D(n20199), .CP(wclk), .Q(ram[15958]) );
  DFF ram_reg_53__5_ ( .D(n20198), .CP(wclk), .Q(ram[15957]) );
  DFF ram_reg_53__4_ ( .D(n20197), .CP(wclk), .Q(ram[15956]) );
  DFF ram_reg_53__3_ ( .D(n20196), .CP(wclk), .Q(ram[15955]) );
  DFF ram_reg_53__2_ ( .D(n20195), .CP(wclk), .Q(ram[15954]) );
  DFF ram_reg_53__1_ ( .D(n20194), .CP(wclk), .Q(ram[15953]) );
  DFF ram_reg_53__0_ ( .D(n20193), .CP(wclk), .Q(ram[15952]) );
  DFF ram_reg_65__7_ ( .D(n20104), .CP(wclk), .Q(ram[15863]) );
  DFF ram_reg_65__6_ ( .D(n20103), .CP(wclk), .Q(ram[15862]) );
  DFF ram_reg_65__5_ ( .D(n20102), .CP(wclk), .Q(ram[15861]) );
  DFF ram_reg_65__4_ ( .D(n20101), .CP(wclk), .Q(ram[15860]) );
  DFF ram_reg_65__3_ ( .D(n20100), .CP(wclk), .Q(ram[15859]) );
  DFF ram_reg_65__2_ ( .D(n20099), .CP(wclk), .Q(ram[15858]) );
  DFF ram_reg_65__1_ ( .D(n20098), .CP(wclk), .Q(ram[15857]) );
  DFF ram_reg_65__0_ ( .D(n20097), .CP(wclk), .Q(ram[15856]) );
  DFF ram_reg_69__7_ ( .D(n20072), .CP(wclk), .Q(ram[15831]) );
  DFF ram_reg_69__6_ ( .D(n20071), .CP(wclk), .Q(ram[15830]) );
  DFF ram_reg_69__5_ ( .D(n20070), .CP(wclk), .Q(ram[15829]) );
  DFF ram_reg_69__4_ ( .D(n20069), .CP(wclk), .Q(ram[15828]) );
  DFF ram_reg_69__3_ ( .D(n20068), .CP(wclk), .Q(ram[15827]) );
  DFF ram_reg_69__2_ ( .D(n20067), .CP(wclk), .Q(ram[15826]) );
  DFF ram_reg_69__1_ ( .D(n20066), .CP(wclk), .Q(ram[15825]) );
  DFF ram_reg_69__0_ ( .D(n20065), .CP(wclk), .Q(ram[15824]) );
  DFF ram_reg_73__7_ ( .D(n20040), .CP(wclk), .Q(ram[15799]) );
  DFF ram_reg_73__6_ ( .D(n20039), .CP(wclk), .Q(ram[15798]) );
  DFF ram_reg_73__5_ ( .D(n20038), .CP(wclk), .Q(ram[15797]) );
  DFF ram_reg_73__4_ ( .D(n20037), .CP(wclk), .Q(ram[15796]) );
  DFF ram_reg_73__3_ ( .D(n20036), .CP(wclk), .Q(ram[15795]) );
  DFF ram_reg_73__2_ ( .D(n20035), .CP(wclk), .Q(ram[15794]) );
  DFF ram_reg_73__1_ ( .D(n20034), .CP(wclk), .Q(ram[15793]) );
  DFF ram_reg_73__0_ ( .D(n20033), .CP(wclk), .Q(ram[15792]) );
  DFF ram_reg_77__7_ ( .D(n20008), .CP(wclk), .Q(ram[15767]) );
  DFF ram_reg_77__6_ ( .D(n20007), .CP(wclk), .Q(ram[15766]) );
  DFF ram_reg_77__5_ ( .D(n20006), .CP(wclk), .Q(ram[15765]) );
  DFF ram_reg_77__4_ ( .D(n20005), .CP(wclk), .Q(ram[15764]) );
  DFF ram_reg_77__3_ ( .D(n20004), .CP(wclk), .Q(ram[15763]) );
  DFF ram_reg_77__2_ ( .D(n20003), .CP(wclk), .Q(ram[15762]) );
  DFF ram_reg_77__1_ ( .D(n20002), .CP(wclk), .Q(ram[15761]) );
  DFF ram_reg_77__0_ ( .D(n20001), .CP(wclk), .Q(ram[15760]) );
  DFF ram_reg_81__7_ ( .D(n19976), .CP(wclk), .Q(ram[15735]) );
  DFF ram_reg_81__6_ ( .D(n19975), .CP(wclk), .Q(ram[15734]) );
  DFF ram_reg_81__5_ ( .D(n19974), .CP(wclk), .Q(ram[15733]) );
  DFF ram_reg_81__4_ ( .D(n19973), .CP(wclk), .Q(ram[15732]) );
  DFF ram_reg_81__3_ ( .D(n19972), .CP(wclk), .Q(ram[15731]) );
  DFF ram_reg_81__2_ ( .D(n19971), .CP(wclk), .Q(ram[15730]) );
  DFF ram_reg_81__1_ ( .D(n19970), .CP(wclk), .Q(ram[15729]) );
  DFF ram_reg_81__0_ ( .D(n19969), .CP(wclk), .Q(ram[15728]) );
  DFF ram_reg_85__7_ ( .D(n19944), .CP(wclk), .Q(ram[15703]) );
  DFF ram_reg_85__6_ ( .D(n19943), .CP(wclk), .Q(ram[15702]) );
  DFF ram_reg_85__5_ ( .D(n19942), .CP(wclk), .Q(ram[15701]) );
  DFF ram_reg_85__4_ ( .D(n19941), .CP(wclk), .Q(ram[15700]) );
  DFF ram_reg_85__3_ ( .D(n19940), .CP(wclk), .Q(ram[15699]) );
  DFF ram_reg_85__2_ ( .D(n19939), .CP(wclk), .Q(ram[15698]) );
  DFF ram_reg_85__1_ ( .D(n19938), .CP(wclk), .Q(ram[15697]) );
  DFF ram_reg_85__0_ ( .D(n19937), .CP(wclk), .Q(ram[15696]) );
  DFF ram_reg_89__7_ ( .D(n19912), .CP(wclk), .Q(ram[15671]) );
  DFF ram_reg_89__6_ ( .D(n19911), .CP(wclk), .Q(ram[15670]) );
  DFF ram_reg_89__5_ ( .D(n19910), .CP(wclk), .Q(ram[15669]) );
  DFF ram_reg_89__4_ ( .D(n19909), .CP(wclk), .Q(ram[15668]) );
  DFF ram_reg_89__3_ ( .D(n19908), .CP(wclk), .Q(ram[15667]) );
  DFF ram_reg_89__2_ ( .D(n19907), .CP(wclk), .Q(ram[15666]) );
  DFF ram_reg_89__1_ ( .D(n19906), .CP(wclk), .Q(ram[15665]) );
  DFF ram_reg_89__0_ ( .D(n19905), .CP(wclk), .Q(ram[15664]) );
  DFF ram_reg_93__7_ ( .D(n19880), .CP(wclk), .Q(ram[15639]) );
  DFF ram_reg_93__6_ ( .D(n19879), .CP(wclk), .Q(ram[15638]) );
  DFF ram_reg_93__5_ ( .D(n19878), .CP(wclk), .Q(ram[15637]) );
  DFF ram_reg_93__4_ ( .D(n19877), .CP(wclk), .Q(ram[15636]) );
  DFF ram_reg_93__3_ ( .D(n19876), .CP(wclk), .Q(ram[15635]) );
  DFF ram_reg_93__2_ ( .D(n19875), .CP(wclk), .Q(ram[15634]) );
  DFF ram_reg_93__1_ ( .D(n19874), .CP(wclk), .Q(ram[15633]) );
  DFF ram_reg_93__0_ ( .D(n19873), .CP(wclk), .Q(ram[15632]) );
  DFF ram_reg_97__7_ ( .D(n19848), .CP(wclk), .Q(ram[15607]) );
  DFF ram_reg_97__6_ ( .D(n19847), .CP(wclk), .Q(ram[15606]) );
  DFF ram_reg_97__5_ ( .D(n19846), .CP(wclk), .Q(ram[15605]) );
  DFF ram_reg_97__4_ ( .D(n19845), .CP(wclk), .Q(ram[15604]) );
  DFF ram_reg_97__3_ ( .D(n19844), .CP(wclk), .Q(ram[15603]) );
  DFF ram_reg_97__2_ ( .D(n19843), .CP(wclk), .Q(ram[15602]) );
  DFF ram_reg_97__1_ ( .D(n19842), .CP(wclk), .Q(ram[15601]) );
  DFF ram_reg_97__0_ ( .D(n19841), .CP(wclk), .Q(ram[15600]) );
  DFF ram_reg_101__7_ ( .D(n19816), .CP(wclk), .Q(ram[15575]) );
  DFF ram_reg_101__6_ ( .D(n19815), .CP(wclk), .Q(ram[15574]) );
  DFF ram_reg_101__5_ ( .D(n19814), .CP(wclk), .Q(ram[15573]) );
  DFF ram_reg_101__4_ ( .D(n19813), .CP(wclk), .Q(ram[15572]) );
  DFF ram_reg_101__3_ ( .D(n19812), .CP(wclk), .Q(ram[15571]) );
  DFF ram_reg_101__2_ ( .D(n19811), .CP(wclk), .Q(ram[15570]) );
  DFF ram_reg_101__1_ ( .D(n19810), .CP(wclk), .Q(ram[15569]) );
  DFF ram_reg_101__0_ ( .D(n19809), .CP(wclk), .Q(ram[15568]) );
  DFF ram_reg_105__7_ ( .D(n19784), .CP(wclk), .Q(ram[15543]) );
  DFF ram_reg_105__6_ ( .D(n19783), .CP(wclk), .Q(ram[15542]) );
  DFF ram_reg_105__5_ ( .D(n19782), .CP(wclk), .Q(ram[15541]) );
  DFF ram_reg_105__4_ ( .D(n19781), .CP(wclk), .Q(ram[15540]) );
  DFF ram_reg_105__3_ ( .D(n19780), .CP(wclk), .Q(ram[15539]) );
  DFF ram_reg_105__2_ ( .D(n19779), .CP(wclk), .Q(ram[15538]) );
  DFF ram_reg_105__1_ ( .D(n19778), .CP(wclk), .Q(ram[15537]) );
  DFF ram_reg_105__0_ ( .D(n19777), .CP(wclk), .Q(ram[15536]) );
  DFF ram_reg_109__7_ ( .D(n19752), .CP(wclk), .Q(ram[15511]) );
  DFF ram_reg_109__6_ ( .D(n19751), .CP(wclk), .Q(ram[15510]) );
  DFF ram_reg_109__5_ ( .D(n19750), .CP(wclk), .Q(ram[15509]) );
  DFF ram_reg_109__4_ ( .D(n19749), .CP(wclk), .Q(ram[15508]) );
  DFF ram_reg_109__3_ ( .D(n19748), .CP(wclk), .Q(ram[15507]) );
  DFF ram_reg_109__2_ ( .D(n19747), .CP(wclk), .Q(ram[15506]) );
  DFF ram_reg_109__1_ ( .D(n19746), .CP(wclk), .Q(ram[15505]) );
  DFF ram_reg_109__0_ ( .D(n19745), .CP(wclk), .Q(ram[15504]) );
  DFF ram_reg_113__7_ ( .D(n19720), .CP(wclk), .Q(ram[15479]) );
  DFF ram_reg_113__6_ ( .D(n19719), .CP(wclk), .Q(ram[15478]) );
  DFF ram_reg_113__5_ ( .D(n19718), .CP(wclk), .Q(ram[15477]) );
  DFF ram_reg_113__4_ ( .D(n19717), .CP(wclk), .Q(ram[15476]) );
  DFF ram_reg_113__3_ ( .D(n19716), .CP(wclk), .Q(ram[15475]) );
  DFF ram_reg_113__2_ ( .D(n19715), .CP(wclk), .Q(ram[15474]) );
  DFF ram_reg_113__1_ ( .D(n19714), .CP(wclk), .Q(ram[15473]) );
  DFF ram_reg_113__0_ ( .D(n19713), .CP(wclk), .Q(ram[15472]) );
  DFF ram_reg_117__7_ ( .D(n19688), .CP(wclk), .Q(ram[15447]) );
  DFF ram_reg_117__6_ ( .D(n19687), .CP(wclk), .Q(ram[15446]) );
  DFF ram_reg_117__5_ ( .D(n19686), .CP(wclk), .Q(ram[15445]) );
  DFF ram_reg_117__4_ ( .D(n19685), .CP(wclk), .Q(ram[15444]) );
  DFF ram_reg_117__3_ ( .D(n19684), .CP(wclk), .Q(ram[15443]) );
  DFF ram_reg_117__2_ ( .D(n19683), .CP(wclk), .Q(ram[15442]) );
  DFF ram_reg_117__1_ ( .D(n19682), .CP(wclk), .Q(ram[15441]) );
  DFF ram_reg_117__0_ ( .D(n19681), .CP(wclk), .Q(ram[15440]) );
  DFF ram_reg_121__7_ ( .D(n19656), .CP(wclk), .Q(ram[15415]) );
  DFF ram_reg_121__6_ ( .D(n19655), .CP(wclk), .Q(ram[15414]) );
  DFF ram_reg_121__5_ ( .D(n19654), .CP(wclk), .Q(ram[15413]) );
  DFF ram_reg_121__4_ ( .D(n19653), .CP(wclk), .Q(ram[15412]) );
  DFF ram_reg_121__3_ ( .D(n19652), .CP(wclk), .Q(ram[15411]) );
  DFF ram_reg_121__2_ ( .D(n19651), .CP(wclk), .Q(ram[15410]) );
  DFF ram_reg_121__1_ ( .D(n19650), .CP(wclk), .Q(ram[15409]) );
  DFF ram_reg_121__0_ ( .D(n19649), .CP(wclk), .Q(ram[15408]) );
  DFF ram_reg_125__7_ ( .D(n19624), .CP(wclk), .Q(ram[15383]) );
  DFF ram_reg_125__6_ ( .D(n19623), .CP(wclk), .Q(ram[15382]) );
  DFF ram_reg_125__5_ ( .D(n19622), .CP(wclk), .Q(ram[15381]) );
  DFF ram_reg_125__4_ ( .D(n19621), .CP(wclk), .Q(ram[15380]) );
  DFF ram_reg_125__3_ ( .D(n19620), .CP(wclk), .Q(ram[15379]) );
  DFF ram_reg_125__2_ ( .D(n19619), .CP(wclk), .Q(ram[15378]) );
  DFF ram_reg_125__1_ ( .D(n19618), .CP(wclk), .Q(ram[15377]) );
  DFF ram_reg_125__0_ ( .D(n19617), .CP(wclk), .Q(ram[15376]) );
  DFF ram_reg_133__7_ ( .D(n19560), .CP(wclk), .Q(ram[15319]) );
  DFF ram_reg_133__6_ ( .D(n19559), .CP(wclk), .Q(ram[15318]) );
  DFF ram_reg_133__5_ ( .D(n19558), .CP(wclk), .Q(ram[15317]) );
  DFF ram_reg_133__4_ ( .D(n19557), .CP(wclk), .Q(ram[15316]) );
  DFF ram_reg_133__3_ ( .D(n19556), .CP(wclk), .Q(ram[15315]) );
  DFF ram_reg_133__2_ ( .D(n19555), .CP(wclk), .Q(ram[15314]) );
  DFF ram_reg_133__1_ ( .D(n19554), .CP(wclk), .Q(ram[15313]) );
  DFF ram_reg_133__0_ ( .D(n19553), .CP(wclk), .Q(ram[15312]) );
  DFF ram_reg_145__7_ ( .D(n19464), .CP(wclk), .Q(ram[15223]) );
  DFF ram_reg_145__6_ ( .D(n19463), .CP(wclk), .Q(ram[15222]) );
  DFF ram_reg_145__5_ ( .D(n19462), .CP(wclk), .Q(ram[15221]) );
  DFF ram_reg_145__4_ ( .D(n19461), .CP(wclk), .Q(ram[15220]) );
  DFF ram_reg_145__3_ ( .D(n19460), .CP(wclk), .Q(ram[15219]) );
  DFF ram_reg_145__2_ ( .D(n19459), .CP(wclk), .Q(ram[15218]) );
  DFF ram_reg_145__1_ ( .D(n19458), .CP(wclk), .Q(ram[15217]) );
  DFF ram_reg_145__0_ ( .D(n19457), .CP(wclk), .Q(ram[15216]) );
  DFF ram_reg_149__7_ ( .D(n19432), .CP(wclk), .Q(ram[15191]) );
  DFF ram_reg_149__6_ ( .D(n19431), .CP(wclk), .Q(ram[15190]) );
  DFF ram_reg_149__5_ ( .D(n19430), .CP(wclk), .Q(ram[15189]) );
  DFF ram_reg_149__4_ ( .D(n19429), .CP(wclk), .Q(ram[15188]) );
  DFF ram_reg_149__3_ ( .D(n19428), .CP(wclk), .Q(ram[15187]) );
  DFF ram_reg_149__2_ ( .D(n19427), .CP(wclk), .Q(ram[15186]) );
  DFF ram_reg_149__1_ ( .D(n19426), .CP(wclk), .Q(ram[15185]) );
  DFF ram_reg_149__0_ ( .D(n19425), .CP(wclk), .Q(ram[15184]) );
  DFF ram_reg_165__7_ ( .D(n19304), .CP(wclk), .Q(ram[15063]) );
  DFF ram_reg_165__6_ ( .D(n19303), .CP(wclk), .Q(ram[15062]) );
  DFF ram_reg_165__5_ ( .D(n19302), .CP(wclk), .Q(ram[15061]) );
  DFF ram_reg_165__4_ ( .D(n19301), .CP(wclk), .Q(ram[15060]) );
  DFF ram_reg_165__3_ ( .D(n19300), .CP(wclk), .Q(ram[15059]) );
  DFF ram_reg_165__2_ ( .D(n19299), .CP(wclk), .Q(ram[15058]) );
  DFF ram_reg_165__1_ ( .D(n19298), .CP(wclk), .Q(ram[15057]) );
  DFF ram_reg_165__0_ ( .D(n19297), .CP(wclk), .Q(ram[15056]) );
  DFF ram_reg_181__7_ ( .D(n19176), .CP(wclk), .Q(ram[14935]) );
  DFF ram_reg_181__6_ ( .D(n19175), .CP(wclk), .Q(ram[14934]) );
  DFF ram_reg_181__5_ ( .D(n19174), .CP(wclk), .Q(ram[14933]) );
  DFF ram_reg_181__4_ ( .D(n19173), .CP(wclk), .Q(ram[14932]) );
  DFF ram_reg_181__3_ ( .D(n19172), .CP(wclk), .Q(ram[14931]) );
  DFF ram_reg_181__2_ ( .D(n19171), .CP(wclk), .Q(ram[14930]) );
  DFF ram_reg_181__1_ ( .D(n19170), .CP(wclk), .Q(ram[14929]) );
  DFF ram_reg_181__0_ ( .D(n19169), .CP(wclk), .Q(ram[14928]) );
  DFF ram_reg_193__7_ ( .D(n19080), .CP(wclk), .Q(ram[14839]) );
  DFF ram_reg_193__6_ ( .D(n19079), .CP(wclk), .Q(ram[14838]) );
  DFF ram_reg_193__5_ ( .D(n19078), .CP(wclk), .Q(ram[14837]) );
  DFF ram_reg_193__4_ ( .D(n19077), .CP(wclk), .Q(ram[14836]) );
  DFF ram_reg_193__3_ ( .D(n19076), .CP(wclk), .Q(ram[14835]) );
  DFF ram_reg_193__2_ ( .D(n19075), .CP(wclk), .Q(ram[14834]) );
  DFF ram_reg_193__1_ ( .D(n19074), .CP(wclk), .Q(ram[14833]) );
  DFF ram_reg_193__0_ ( .D(n19073), .CP(wclk), .Q(ram[14832]) );
  DFF ram_reg_197__7_ ( .D(n19048), .CP(wclk), .Q(ram[14807]) );
  DFF ram_reg_197__6_ ( .D(n19047), .CP(wclk), .Q(ram[14806]) );
  DFF ram_reg_197__5_ ( .D(n19046), .CP(wclk), .Q(ram[14805]) );
  DFF ram_reg_197__4_ ( .D(n19045), .CP(wclk), .Q(ram[14804]) );
  DFF ram_reg_197__3_ ( .D(n19044), .CP(wclk), .Q(ram[14803]) );
  DFF ram_reg_197__2_ ( .D(n19043), .CP(wclk), .Q(ram[14802]) );
  DFF ram_reg_197__1_ ( .D(n19042), .CP(wclk), .Q(ram[14801]) );
  DFF ram_reg_197__0_ ( .D(n19041), .CP(wclk), .Q(ram[14800]) );
  DFF ram_reg_209__7_ ( .D(n18952), .CP(wclk), .Q(ram[14711]) );
  DFF ram_reg_209__6_ ( .D(n18951), .CP(wclk), .Q(ram[14710]) );
  DFF ram_reg_209__5_ ( .D(n18950), .CP(wclk), .Q(ram[14709]) );
  DFF ram_reg_209__4_ ( .D(n18949), .CP(wclk), .Q(ram[14708]) );
  DFF ram_reg_209__3_ ( .D(n18948), .CP(wclk), .Q(ram[14707]) );
  DFF ram_reg_209__2_ ( .D(n18947), .CP(wclk), .Q(ram[14706]) );
  DFF ram_reg_209__1_ ( .D(n18946), .CP(wclk), .Q(ram[14705]) );
  DFF ram_reg_209__0_ ( .D(n18945), .CP(wclk), .Q(ram[14704]) );
  DFF ram_reg_213__7_ ( .D(n18920), .CP(wclk), .Q(ram[14679]) );
  DFF ram_reg_213__6_ ( .D(n18919), .CP(wclk), .Q(ram[14678]) );
  DFF ram_reg_213__5_ ( .D(n18918), .CP(wclk), .Q(ram[14677]) );
  DFF ram_reg_213__4_ ( .D(n18917), .CP(wclk), .Q(ram[14676]) );
  DFF ram_reg_213__3_ ( .D(n18916), .CP(wclk), .Q(ram[14675]) );
  DFF ram_reg_213__2_ ( .D(n18915), .CP(wclk), .Q(ram[14674]) );
  DFF ram_reg_213__1_ ( .D(n18914), .CP(wclk), .Q(ram[14673]) );
  DFF ram_reg_213__0_ ( .D(n18913), .CP(wclk), .Q(ram[14672]) );
  DFF ram_reg_229__7_ ( .D(n18792), .CP(wclk), .Q(ram[14551]) );
  DFF ram_reg_229__6_ ( .D(n18791), .CP(wclk), .Q(ram[14550]) );
  DFF ram_reg_229__5_ ( .D(n18790), .CP(wclk), .Q(ram[14549]) );
  DFF ram_reg_229__4_ ( .D(n18789), .CP(wclk), .Q(ram[14548]) );
  DFF ram_reg_229__3_ ( .D(n18788), .CP(wclk), .Q(ram[14547]) );
  DFF ram_reg_229__2_ ( .D(n18787), .CP(wclk), .Q(ram[14546]) );
  DFF ram_reg_229__1_ ( .D(n18786), .CP(wclk), .Q(ram[14545]) );
  DFF ram_reg_229__0_ ( .D(n18785), .CP(wclk), .Q(ram[14544]) );
  DFF ram_reg_245__7_ ( .D(n18664), .CP(wclk), .Q(ram[14423]) );
  DFF ram_reg_245__6_ ( .D(n18663), .CP(wclk), .Q(ram[14422]) );
  DFF ram_reg_245__5_ ( .D(n18662), .CP(wclk), .Q(ram[14421]) );
  DFF ram_reg_245__4_ ( .D(n18661), .CP(wclk), .Q(ram[14420]) );
  DFF ram_reg_245__3_ ( .D(n18660), .CP(wclk), .Q(ram[14419]) );
  DFF ram_reg_245__2_ ( .D(n18659), .CP(wclk), .Q(ram[14418]) );
  DFF ram_reg_245__1_ ( .D(n18658), .CP(wclk), .Q(ram[14417]) );
  DFF ram_reg_245__0_ ( .D(n18657), .CP(wclk), .Q(ram[14416]) );
  DFF ram_reg_257__7_ ( .D(n18568), .CP(wclk), .Q(ram[14327]) );
  DFF ram_reg_257__6_ ( .D(n18567), .CP(wclk), .Q(ram[14326]) );
  DFF ram_reg_257__5_ ( .D(n18566), .CP(wclk), .Q(ram[14325]) );
  DFF ram_reg_257__4_ ( .D(n18565), .CP(wclk), .Q(ram[14324]) );
  DFF ram_reg_257__3_ ( .D(n18564), .CP(wclk), .Q(ram[14323]) );
  DFF ram_reg_257__2_ ( .D(n18563), .CP(wclk), .Q(ram[14322]) );
  DFF ram_reg_257__1_ ( .D(n18562), .CP(wclk), .Q(ram[14321]) );
  DFF ram_reg_257__0_ ( .D(n18561), .CP(wclk), .Q(ram[14320]) );
  DFF ram_reg_261__7_ ( .D(n18536), .CP(wclk), .Q(ram[14295]) );
  DFF ram_reg_261__6_ ( .D(n18535), .CP(wclk), .Q(ram[14294]) );
  DFF ram_reg_261__5_ ( .D(n18534), .CP(wclk), .Q(ram[14293]) );
  DFF ram_reg_261__4_ ( .D(n18533), .CP(wclk), .Q(ram[14292]) );
  DFF ram_reg_261__3_ ( .D(n18532), .CP(wclk), .Q(ram[14291]) );
  DFF ram_reg_261__2_ ( .D(n18531), .CP(wclk), .Q(ram[14290]) );
  DFF ram_reg_261__1_ ( .D(n18530), .CP(wclk), .Q(ram[14289]) );
  DFF ram_reg_261__0_ ( .D(n18529), .CP(wclk), .Q(ram[14288]) );
  DFF ram_reg_269__7_ ( .D(n18472), .CP(wclk), .Q(ram[14231]) );
  DFF ram_reg_269__6_ ( .D(n18471), .CP(wclk), .Q(ram[14230]) );
  DFF ram_reg_269__5_ ( .D(n18470), .CP(wclk), .Q(ram[14229]) );
  DFF ram_reg_269__4_ ( .D(n18469), .CP(wclk), .Q(ram[14228]) );
  DFF ram_reg_269__3_ ( .D(n18468), .CP(wclk), .Q(ram[14227]) );
  DFF ram_reg_269__2_ ( .D(n18467), .CP(wclk), .Q(ram[14226]) );
  DFF ram_reg_269__1_ ( .D(n18466), .CP(wclk), .Q(ram[14225]) );
  DFF ram_reg_269__0_ ( .D(n18465), .CP(wclk), .Q(ram[14224]) );
  DFF ram_reg_273__7_ ( .D(n18440), .CP(wclk), .Q(ram[14199]) );
  DFF ram_reg_273__6_ ( .D(n18439), .CP(wclk), .Q(ram[14198]) );
  DFF ram_reg_273__5_ ( .D(n18438), .CP(wclk), .Q(ram[14197]) );
  DFF ram_reg_273__4_ ( .D(n18437), .CP(wclk), .Q(ram[14196]) );
  DFF ram_reg_273__3_ ( .D(n18436), .CP(wclk), .Q(ram[14195]) );
  DFF ram_reg_273__2_ ( .D(n18435), .CP(wclk), .Q(ram[14194]) );
  DFF ram_reg_273__1_ ( .D(n18434), .CP(wclk), .Q(ram[14193]) );
  DFF ram_reg_273__0_ ( .D(n18433), .CP(wclk), .Q(ram[14192]) );
  DFF ram_reg_277__7_ ( .D(n18408), .CP(wclk), .Q(ram[14167]) );
  DFF ram_reg_277__6_ ( .D(n18407), .CP(wclk), .Q(ram[14166]) );
  DFF ram_reg_277__5_ ( .D(n18406), .CP(wclk), .Q(ram[14165]) );
  DFF ram_reg_277__4_ ( .D(n18405), .CP(wclk), .Q(ram[14164]) );
  DFF ram_reg_277__3_ ( .D(n18404), .CP(wclk), .Q(ram[14163]) );
  DFF ram_reg_277__2_ ( .D(n18403), .CP(wclk), .Q(ram[14162]) );
  DFF ram_reg_277__1_ ( .D(n18402), .CP(wclk), .Q(ram[14161]) );
  DFF ram_reg_277__0_ ( .D(n18401), .CP(wclk), .Q(ram[14160]) );
  DFF ram_reg_281__7_ ( .D(n18376), .CP(wclk), .Q(ram[14135]) );
  DFF ram_reg_281__6_ ( .D(n18375), .CP(wclk), .Q(ram[14134]) );
  DFF ram_reg_281__5_ ( .D(n18374), .CP(wclk), .Q(ram[14133]) );
  DFF ram_reg_281__4_ ( .D(n18373), .CP(wclk), .Q(ram[14132]) );
  DFF ram_reg_281__3_ ( .D(n18372), .CP(wclk), .Q(ram[14131]) );
  DFF ram_reg_281__2_ ( .D(n18371), .CP(wclk), .Q(ram[14130]) );
  DFF ram_reg_281__1_ ( .D(n18370), .CP(wclk), .Q(ram[14129]) );
  DFF ram_reg_281__0_ ( .D(n18369), .CP(wclk), .Q(ram[14128]) );
  DFF ram_reg_285__7_ ( .D(n18344), .CP(wclk), .Q(ram[14103]) );
  DFF ram_reg_285__6_ ( .D(n18343), .CP(wclk), .Q(ram[14102]) );
  DFF ram_reg_285__5_ ( .D(n18342), .CP(wclk), .Q(ram[14101]) );
  DFF ram_reg_285__4_ ( .D(n18341), .CP(wclk), .Q(ram[14100]) );
  DFF ram_reg_285__3_ ( .D(n18340), .CP(wclk), .Q(ram[14099]) );
  DFF ram_reg_285__2_ ( .D(n18339), .CP(wclk), .Q(ram[14098]) );
  DFF ram_reg_285__1_ ( .D(n18338), .CP(wclk), .Q(ram[14097]) );
  DFF ram_reg_285__0_ ( .D(n18337), .CP(wclk), .Q(ram[14096]) );
  DFF ram_reg_289__7_ ( .D(n18312), .CP(wclk), .Q(ram[14071]) );
  DFF ram_reg_289__6_ ( .D(n18311), .CP(wclk), .Q(ram[14070]) );
  DFF ram_reg_289__5_ ( .D(n18310), .CP(wclk), .Q(ram[14069]) );
  DFF ram_reg_289__4_ ( .D(n18309), .CP(wclk), .Q(ram[14068]) );
  DFF ram_reg_289__3_ ( .D(n18308), .CP(wclk), .Q(ram[14067]) );
  DFF ram_reg_289__2_ ( .D(n18307), .CP(wclk), .Q(ram[14066]) );
  DFF ram_reg_289__1_ ( .D(n18306), .CP(wclk), .Q(ram[14065]) );
  DFF ram_reg_289__0_ ( .D(n18305), .CP(wclk), .Q(ram[14064]) );
  DFF ram_reg_293__7_ ( .D(n18280), .CP(wclk), .Q(ram[14039]) );
  DFF ram_reg_293__6_ ( .D(n18279), .CP(wclk), .Q(ram[14038]) );
  DFF ram_reg_293__5_ ( .D(n18278), .CP(wclk), .Q(ram[14037]) );
  DFF ram_reg_293__4_ ( .D(n18277), .CP(wclk), .Q(ram[14036]) );
  DFF ram_reg_293__3_ ( .D(n18276), .CP(wclk), .Q(ram[14035]) );
  DFF ram_reg_293__2_ ( .D(n18275), .CP(wclk), .Q(ram[14034]) );
  DFF ram_reg_293__1_ ( .D(n18274), .CP(wclk), .Q(ram[14033]) );
  DFF ram_reg_293__0_ ( .D(n18273), .CP(wclk), .Q(ram[14032]) );
  DFF ram_reg_305__7_ ( .D(n18184), .CP(wclk), .Q(ram[13943]) );
  DFF ram_reg_305__6_ ( .D(n18183), .CP(wclk), .Q(ram[13942]) );
  DFF ram_reg_305__5_ ( .D(n18182), .CP(wclk), .Q(ram[13941]) );
  DFF ram_reg_305__4_ ( .D(n18181), .CP(wclk), .Q(ram[13940]) );
  DFF ram_reg_305__3_ ( .D(n18180), .CP(wclk), .Q(ram[13939]) );
  DFF ram_reg_305__2_ ( .D(n18179), .CP(wclk), .Q(ram[13938]) );
  DFF ram_reg_305__1_ ( .D(n18178), .CP(wclk), .Q(ram[13937]) );
  DFF ram_reg_305__0_ ( .D(n18177), .CP(wclk), .Q(ram[13936]) );
  DFF ram_reg_309__7_ ( .D(n18152), .CP(wclk), .Q(ram[13911]) );
  DFF ram_reg_309__6_ ( .D(n18151), .CP(wclk), .Q(ram[13910]) );
  DFF ram_reg_309__5_ ( .D(n18150), .CP(wclk), .Q(ram[13909]) );
  DFF ram_reg_309__4_ ( .D(n18149), .CP(wclk), .Q(ram[13908]) );
  DFF ram_reg_309__3_ ( .D(n18148), .CP(wclk), .Q(ram[13907]) );
  DFF ram_reg_309__2_ ( .D(n18147), .CP(wclk), .Q(ram[13906]) );
  DFF ram_reg_309__1_ ( .D(n18146), .CP(wclk), .Q(ram[13905]) );
  DFF ram_reg_309__0_ ( .D(n18145), .CP(wclk), .Q(ram[13904]) );
  DFF ram_reg_321__7_ ( .D(n18056), .CP(wclk), .Q(ram[13815]) );
  DFF ram_reg_321__6_ ( .D(n18055), .CP(wclk), .Q(ram[13814]) );
  DFF ram_reg_321__5_ ( .D(n18054), .CP(wclk), .Q(ram[13813]) );
  DFF ram_reg_321__4_ ( .D(n18053), .CP(wclk), .Q(ram[13812]) );
  DFF ram_reg_321__3_ ( .D(n18052), .CP(wclk), .Q(ram[13811]) );
  DFF ram_reg_321__2_ ( .D(n18051), .CP(wclk), .Q(ram[13810]) );
  DFF ram_reg_321__1_ ( .D(n18050), .CP(wclk), .Q(ram[13809]) );
  DFF ram_reg_321__0_ ( .D(n18049), .CP(wclk), .Q(ram[13808]) );
  DFF ram_reg_325__7_ ( .D(n18024), .CP(wclk), .Q(ram[13783]) );
  DFF ram_reg_325__6_ ( .D(n18023), .CP(wclk), .Q(ram[13782]) );
  DFF ram_reg_325__5_ ( .D(n18022), .CP(wclk), .Q(ram[13781]) );
  DFF ram_reg_325__4_ ( .D(n18021), .CP(wclk), .Q(ram[13780]) );
  DFF ram_reg_325__3_ ( .D(n18020), .CP(wclk), .Q(ram[13779]) );
  DFF ram_reg_325__2_ ( .D(n18019), .CP(wclk), .Q(ram[13778]) );
  DFF ram_reg_325__1_ ( .D(n18018), .CP(wclk), .Q(ram[13777]) );
  DFF ram_reg_325__0_ ( .D(n18017), .CP(wclk), .Q(ram[13776]) );
  DFF ram_reg_329__7_ ( .D(n17992), .CP(wclk), .Q(ram[13751]) );
  DFF ram_reg_329__6_ ( .D(n17991), .CP(wclk), .Q(ram[13750]) );
  DFF ram_reg_329__5_ ( .D(n17990), .CP(wclk), .Q(ram[13749]) );
  DFF ram_reg_329__4_ ( .D(n17989), .CP(wclk), .Q(ram[13748]) );
  DFF ram_reg_329__3_ ( .D(n17988), .CP(wclk), .Q(ram[13747]) );
  DFF ram_reg_329__2_ ( .D(n17987), .CP(wclk), .Q(ram[13746]) );
  DFF ram_reg_329__1_ ( .D(n17986), .CP(wclk), .Q(ram[13745]) );
  DFF ram_reg_329__0_ ( .D(n17985), .CP(wclk), .Q(ram[13744]) );
  DFF ram_reg_333__7_ ( .D(n17960), .CP(wclk), .Q(ram[13719]) );
  DFF ram_reg_333__6_ ( .D(n17959), .CP(wclk), .Q(ram[13718]) );
  DFF ram_reg_333__5_ ( .D(n17958), .CP(wclk), .Q(ram[13717]) );
  DFF ram_reg_333__4_ ( .D(n17957), .CP(wclk), .Q(ram[13716]) );
  DFF ram_reg_333__3_ ( .D(n17956), .CP(wclk), .Q(ram[13715]) );
  DFF ram_reg_333__2_ ( .D(n17955), .CP(wclk), .Q(ram[13714]) );
  DFF ram_reg_333__1_ ( .D(n17954), .CP(wclk), .Q(ram[13713]) );
  DFF ram_reg_333__0_ ( .D(n17953), .CP(wclk), .Q(ram[13712]) );
  DFF ram_reg_337__7_ ( .D(n17928), .CP(wclk), .Q(ram[13687]) );
  DFF ram_reg_337__6_ ( .D(n17927), .CP(wclk), .Q(ram[13686]) );
  DFF ram_reg_337__5_ ( .D(n17926), .CP(wclk), .Q(ram[13685]) );
  DFF ram_reg_337__4_ ( .D(n17925), .CP(wclk), .Q(ram[13684]) );
  DFF ram_reg_337__3_ ( .D(n17924), .CP(wclk), .Q(ram[13683]) );
  DFF ram_reg_337__2_ ( .D(n17923), .CP(wclk), .Q(ram[13682]) );
  DFF ram_reg_337__1_ ( .D(n17922), .CP(wclk), .Q(ram[13681]) );
  DFF ram_reg_337__0_ ( .D(n17921), .CP(wclk), .Q(ram[13680]) );
  DFF ram_reg_341__7_ ( .D(n17896), .CP(wclk), .Q(ram[13655]) );
  DFF ram_reg_341__6_ ( .D(n17895), .CP(wclk), .Q(ram[13654]) );
  DFF ram_reg_341__5_ ( .D(n17894), .CP(wclk), .Q(ram[13653]) );
  DFF ram_reg_341__4_ ( .D(n17893), .CP(wclk), .Q(ram[13652]) );
  DFF ram_reg_341__3_ ( .D(n17892), .CP(wclk), .Q(ram[13651]) );
  DFF ram_reg_341__2_ ( .D(n17891), .CP(wclk), .Q(ram[13650]) );
  DFF ram_reg_341__1_ ( .D(n17890), .CP(wclk), .Q(ram[13649]) );
  DFF ram_reg_341__0_ ( .D(n17889), .CP(wclk), .Q(ram[13648]) );
  DFF ram_reg_345__7_ ( .D(n17864), .CP(wclk), .Q(ram[13623]) );
  DFF ram_reg_345__6_ ( .D(n17863), .CP(wclk), .Q(ram[13622]) );
  DFF ram_reg_345__5_ ( .D(n17862), .CP(wclk), .Q(ram[13621]) );
  DFF ram_reg_345__4_ ( .D(n17861), .CP(wclk), .Q(ram[13620]) );
  DFF ram_reg_345__3_ ( .D(n17860), .CP(wclk), .Q(ram[13619]) );
  DFF ram_reg_345__2_ ( .D(n17859), .CP(wclk), .Q(ram[13618]) );
  DFF ram_reg_345__1_ ( .D(n17858), .CP(wclk), .Q(ram[13617]) );
  DFF ram_reg_345__0_ ( .D(n17857), .CP(wclk), .Q(ram[13616]) );
  DFF ram_reg_349__7_ ( .D(n17832), .CP(wclk), .Q(ram[13591]) );
  DFF ram_reg_349__6_ ( .D(n17831), .CP(wclk), .Q(ram[13590]) );
  DFF ram_reg_349__5_ ( .D(n17830), .CP(wclk), .Q(ram[13589]) );
  DFF ram_reg_349__4_ ( .D(n17829), .CP(wclk), .Q(ram[13588]) );
  DFF ram_reg_349__3_ ( .D(n17828), .CP(wclk), .Q(ram[13587]) );
  DFF ram_reg_349__2_ ( .D(n17827), .CP(wclk), .Q(ram[13586]) );
  DFF ram_reg_349__1_ ( .D(n17826), .CP(wclk), .Q(ram[13585]) );
  DFF ram_reg_349__0_ ( .D(n17825), .CP(wclk), .Q(ram[13584]) );
  DFF ram_reg_353__7_ ( .D(n17800), .CP(wclk), .Q(ram[13559]) );
  DFF ram_reg_353__6_ ( .D(n17799), .CP(wclk), .Q(ram[13558]) );
  DFF ram_reg_353__5_ ( .D(n17798), .CP(wclk), .Q(ram[13557]) );
  DFF ram_reg_353__4_ ( .D(n17797), .CP(wclk), .Q(ram[13556]) );
  DFF ram_reg_353__3_ ( .D(n17796), .CP(wclk), .Q(ram[13555]) );
  DFF ram_reg_353__2_ ( .D(n17795), .CP(wclk), .Q(ram[13554]) );
  DFF ram_reg_353__1_ ( .D(n17794), .CP(wclk), .Q(ram[13553]) );
  DFF ram_reg_353__0_ ( .D(n17793), .CP(wclk), .Q(ram[13552]) );
  DFF ram_reg_357__7_ ( .D(n17768), .CP(wclk), .Q(ram[13527]) );
  DFF ram_reg_357__6_ ( .D(n17767), .CP(wclk), .Q(ram[13526]) );
  DFF ram_reg_357__5_ ( .D(n17766), .CP(wclk), .Q(ram[13525]) );
  DFF ram_reg_357__4_ ( .D(n17765), .CP(wclk), .Q(ram[13524]) );
  DFF ram_reg_357__3_ ( .D(n17764), .CP(wclk), .Q(ram[13523]) );
  DFF ram_reg_357__2_ ( .D(n17763), .CP(wclk), .Q(ram[13522]) );
  DFF ram_reg_357__1_ ( .D(n17762), .CP(wclk), .Q(ram[13521]) );
  DFF ram_reg_357__0_ ( .D(n17761), .CP(wclk), .Q(ram[13520]) );
  DFF ram_reg_361__7_ ( .D(n17736), .CP(wclk), .Q(ram[13495]) );
  DFF ram_reg_361__6_ ( .D(n17735), .CP(wclk), .Q(ram[13494]) );
  DFF ram_reg_361__5_ ( .D(n17734), .CP(wclk), .Q(ram[13493]) );
  DFF ram_reg_361__4_ ( .D(n17733), .CP(wclk), .Q(ram[13492]) );
  DFF ram_reg_361__3_ ( .D(n17732), .CP(wclk), .Q(ram[13491]) );
  DFF ram_reg_361__2_ ( .D(n17731), .CP(wclk), .Q(ram[13490]) );
  DFF ram_reg_361__1_ ( .D(n17730), .CP(wclk), .Q(ram[13489]) );
  DFF ram_reg_361__0_ ( .D(n17729), .CP(wclk), .Q(ram[13488]) );
  DFF ram_reg_365__7_ ( .D(n17704), .CP(wclk), .Q(ram[13463]) );
  DFF ram_reg_365__6_ ( .D(n17703), .CP(wclk), .Q(ram[13462]) );
  DFF ram_reg_365__5_ ( .D(n17702), .CP(wclk), .Q(ram[13461]) );
  DFF ram_reg_365__4_ ( .D(n17701), .CP(wclk), .Q(ram[13460]) );
  DFF ram_reg_365__3_ ( .D(n17700), .CP(wclk), .Q(ram[13459]) );
  DFF ram_reg_365__2_ ( .D(n17699), .CP(wclk), .Q(ram[13458]) );
  DFF ram_reg_365__1_ ( .D(n17698), .CP(wclk), .Q(ram[13457]) );
  DFF ram_reg_365__0_ ( .D(n17697), .CP(wclk), .Q(ram[13456]) );
  DFF ram_reg_369__7_ ( .D(n17672), .CP(wclk), .Q(ram[13431]) );
  DFF ram_reg_369__6_ ( .D(n17671), .CP(wclk), .Q(ram[13430]) );
  DFF ram_reg_369__5_ ( .D(n17670), .CP(wclk), .Q(ram[13429]) );
  DFF ram_reg_369__4_ ( .D(n17669), .CP(wclk), .Q(ram[13428]) );
  DFF ram_reg_369__3_ ( .D(n17668), .CP(wclk), .Q(ram[13427]) );
  DFF ram_reg_369__2_ ( .D(n17667), .CP(wclk), .Q(ram[13426]) );
  DFF ram_reg_369__1_ ( .D(n17666), .CP(wclk), .Q(ram[13425]) );
  DFF ram_reg_369__0_ ( .D(n17665), .CP(wclk), .Q(ram[13424]) );
  DFF ram_reg_373__7_ ( .D(n17640), .CP(wclk), .Q(ram[13399]) );
  DFF ram_reg_373__6_ ( .D(n17639), .CP(wclk), .Q(ram[13398]) );
  DFF ram_reg_373__5_ ( .D(n17638), .CP(wclk), .Q(ram[13397]) );
  DFF ram_reg_373__4_ ( .D(n17637), .CP(wclk), .Q(ram[13396]) );
  DFF ram_reg_373__3_ ( .D(n17636), .CP(wclk), .Q(ram[13395]) );
  DFF ram_reg_373__2_ ( .D(n17635), .CP(wclk), .Q(ram[13394]) );
  DFF ram_reg_373__1_ ( .D(n17634), .CP(wclk), .Q(ram[13393]) );
  DFF ram_reg_373__0_ ( .D(n17633), .CP(wclk), .Q(ram[13392]) );
  DFF ram_reg_381__7_ ( .D(n17576), .CP(wclk), .Q(ram[13335]) );
  DFF ram_reg_381__6_ ( .D(n17575), .CP(wclk), .Q(ram[13334]) );
  DFF ram_reg_381__5_ ( .D(n17574), .CP(wclk), .Q(ram[13333]) );
  DFF ram_reg_381__4_ ( .D(n17573), .CP(wclk), .Q(ram[13332]) );
  DFF ram_reg_381__3_ ( .D(n17572), .CP(wclk), .Q(ram[13331]) );
  DFF ram_reg_381__2_ ( .D(n17571), .CP(wclk), .Q(ram[13330]) );
  DFF ram_reg_381__1_ ( .D(n17570), .CP(wclk), .Q(ram[13329]) );
  DFF ram_reg_381__0_ ( .D(n17569), .CP(wclk), .Q(ram[13328]) );
  DFF ram_reg_389__7_ ( .D(n17512), .CP(wclk), .Q(ram[13271]) );
  DFF ram_reg_389__6_ ( .D(n17511), .CP(wclk), .Q(ram[13270]) );
  DFF ram_reg_389__5_ ( .D(n17510), .CP(wclk), .Q(ram[13269]) );
  DFF ram_reg_389__4_ ( .D(n17509), .CP(wclk), .Q(ram[13268]) );
  DFF ram_reg_389__3_ ( .D(n17508), .CP(wclk), .Q(ram[13267]) );
  DFF ram_reg_389__2_ ( .D(n17507), .CP(wclk), .Q(ram[13266]) );
  DFF ram_reg_389__1_ ( .D(n17506), .CP(wclk), .Q(ram[13265]) );
  DFF ram_reg_389__0_ ( .D(n17505), .CP(wclk), .Q(ram[13264]) );
  DFF ram_reg_401__7_ ( .D(n17416), .CP(wclk), .Q(ram[13175]) );
  DFF ram_reg_401__6_ ( .D(n17415), .CP(wclk), .Q(ram[13174]) );
  DFF ram_reg_401__5_ ( .D(n17414), .CP(wclk), .Q(ram[13173]) );
  DFF ram_reg_401__4_ ( .D(n17413), .CP(wclk), .Q(ram[13172]) );
  DFF ram_reg_401__3_ ( .D(n17412), .CP(wclk), .Q(ram[13171]) );
  DFF ram_reg_401__2_ ( .D(n17411), .CP(wclk), .Q(ram[13170]) );
  DFF ram_reg_401__1_ ( .D(n17410), .CP(wclk), .Q(ram[13169]) );
  DFF ram_reg_401__0_ ( .D(n17409), .CP(wclk), .Q(ram[13168]) );
  DFF ram_reg_405__7_ ( .D(n17384), .CP(wclk), .Q(ram[13143]) );
  DFF ram_reg_405__6_ ( .D(n17383), .CP(wclk), .Q(ram[13142]) );
  DFF ram_reg_405__5_ ( .D(n17382), .CP(wclk), .Q(ram[13141]) );
  DFF ram_reg_405__4_ ( .D(n17381), .CP(wclk), .Q(ram[13140]) );
  DFF ram_reg_405__3_ ( .D(n17380), .CP(wclk), .Q(ram[13139]) );
  DFF ram_reg_405__2_ ( .D(n17379), .CP(wclk), .Q(ram[13138]) );
  DFF ram_reg_405__1_ ( .D(n17378), .CP(wclk), .Q(ram[13137]) );
  DFF ram_reg_405__0_ ( .D(n17377), .CP(wclk), .Q(ram[13136]) );
  DFF ram_reg_421__7_ ( .D(n17256), .CP(wclk), .Q(ram[13015]) );
  DFF ram_reg_421__6_ ( .D(n17255), .CP(wclk), .Q(ram[13014]) );
  DFF ram_reg_421__5_ ( .D(n17254), .CP(wclk), .Q(ram[13013]) );
  DFF ram_reg_421__4_ ( .D(n17253), .CP(wclk), .Q(ram[13012]) );
  DFF ram_reg_421__3_ ( .D(n17252), .CP(wclk), .Q(ram[13011]) );
  DFF ram_reg_421__2_ ( .D(n17251), .CP(wclk), .Q(ram[13010]) );
  DFF ram_reg_421__1_ ( .D(n17250), .CP(wclk), .Q(ram[13009]) );
  DFF ram_reg_421__0_ ( .D(n17249), .CP(wclk), .Q(ram[13008]) );
  DFF ram_reg_449__7_ ( .D(n17032), .CP(wclk), .Q(ram[12791]) );
  DFF ram_reg_449__6_ ( .D(n17031), .CP(wclk), .Q(ram[12790]) );
  DFF ram_reg_449__5_ ( .D(n17030), .CP(wclk), .Q(ram[12789]) );
  DFF ram_reg_449__4_ ( .D(n17029), .CP(wclk), .Q(ram[12788]) );
  DFF ram_reg_449__3_ ( .D(n17028), .CP(wclk), .Q(ram[12787]) );
  DFF ram_reg_449__2_ ( .D(n17027), .CP(wclk), .Q(ram[12786]) );
  DFF ram_reg_449__1_ ( .D(n17026), .CP(wclk), .Q(ram[12785]) );
  DFF ram_reg_449__0_ ( .D(n17025), .CP(wclk), .Q(ram[12784]) );
  DFF ram_reg_453__7_ ( .D(n17000), .CP(wclk), .Q(ram[12759]) );
  DFF ram_reg_453__6_ ( .D(n16999), .CP(wclk), .Q(ram[12758]) );
  DFF ram_reg_453__5_ ( .D(n16998), .CP(wclk), .Q(ram[12757]) );
  DFF ram_reg_453__4_ ( .D(n16997), .CP(wclk), .Q(ram[12756]) );
  DFF ram_reg_453__3_ ( .D(n16996), .CP(wclk), .Q(ram[12755]) );
  DFF ram_reg_453__2_ ( .D(n16995), .CP(wclk), .Q(ram[12754]) );
  DFF ram_reg_453__1_ ( .D(n16994), .CP(wclk), .Q(ram[12753]) );
  DFF ram_reg_453__0_ ( .D(n16993), .CP(wclk), .Q(ram[12752]) );
  DFF ram_reg_465__7_ ( .D(n16904), .CP(wclk), .Q(ram[12663]) );
  DFF ram_reg_465__6_ ( .D(n16903), .CP(wclk), .Q(ram[12662]) );
  DFF ram_reg_465__5_ ( .D(n16902), .CP(wclk), .Q(ram[12661]) );
  DFF ram_reg_465__4_ ( .D(n16901), .CP(wclk), .Q(ram[12660]) );
  DFF ram_reg_465__3_ ( .D(n16900), .CP(wclk), .Q(ram[12659]) );
  DFF ram_reg_465__2_ ( .D(n16899), .CP(wclk), .Q(ram[12658]) );
  DFF ram_reg_465__1_ ( .D(n16898), .CP(wclk), .Q(ram[12657]) );
  DFF ram_reg_465__0_ ( .D(n16897), .CP(wclk), .Q(ram[12656]) );
  DFF ram_reg_469__7_ ( .D(n16872), .CP(wclk), .Q(ram[12631]) );
  DFF ram_reg_469__6_ ( .D(n16871), .CP(wclk), .Q(ram[12630]) );
  DFF ram_reg_469__5_ ( .D(n16870), .CP(wclk), .Q(ram[12629]) );
  DFF ram_reg_469__4_ ( .D(n16869), .CP(wclk), .Q(ram[12628]) );
  DFF ram_reg_469__3_ ( .D(n16868), .CP(wclk), .Q(ram[12627]) );
  DFF ram_reg_469__2_ ( .D(n16867), .CP(wclk), .Q(ram[12626]) );
  DFF ram_reg_469__1_ ( .D(n16866), .CP(wclk), .Q(ram[12625]) );
  DFF ram_reg_469__0_ ( .D(n16865), .CP(wclk), .Q(ram[12624]) );
  DFF ram_reg_485__7_ ( .D(n16744), .CP(wclk), .Q(ram[12503]) );
  DFF ram_reg_485__6_ ( .D(n16743), .CP(wclk), .Q(ram[12502]) );
  DFF ram_reg_485__5_ ( .D(n16742), .CP(wclk), .Q(ram[12501]) );
  DFF ram_reg_485__4_ ( .D(n16741), .CP(wclk), .Q(ram[12500]) );
  DFF ram_reg_485__3_ ( .D(n16740), .CP(wclk), .Q(ram[12499]) );
  DFF ram_reg_485__2_ ( .D(n16739), .CP(wclk), .Q(ram[12498]) );
  DFF ram_reg_485__1_ ( .D(n16738), .CP(wclk), .Q(ram[12497]) );
  DFF ram_reg_485__0_ ( .D(n16737), .CP(wclk), .Q(ram[12496]) );
  DFF ram_reg_501__7_ ( .D(n16616), .CP(wclk), .Q(ram[12375]) );
  DFF ram_reg_501__6_ ( .D(n16615), .CP(wclk), .Q(ram[12374]) );
  DFF ram_reg_501__5_ ( .D(n16614), .CP(wclk), .Q(ram[12373]) );
  DFF ram_reg_501__4_ ( .D(n16613), .CP(wclk), .Q(ram[12372]) );
  DFF ram_reg_501__3_ ( .D(n16612), .CP(wclk), .Q(ram[12371]) );
  DFF ram_reg_501__2_ ( .D(n16611), .CP(wclk), .Q(ram[12370]) );
  DFF ram_reg_501__1_ ( .D(n16610), .CP(wclk), .Q(ram[12369]) );
  DFF ram_reg_501__0_ ( .D(n16609), .CP(wclk), .Q(ram[12368]) );
  DFF ram_reg_513__7_ ( .D(n16520), .CP(wclk), .Q(ram[12279]) );
  DFF ram_reg_513__6_ ( .D(n16519), .CP(wclk), .Q(ram[12278]) );
  DFF ram_reg_513__5_ ( .D(n16518), .CP(wclk), .Q(ram[12277]) );
  DFF ram_reg_513__4_ ( .D(n16517), .CP(wclk), .Q(ram[12276]) );
  DFF ram_reg_513__3_ ( .D(n16516), .CP(wclk), .Q(ram[12275]) );
  DFF ram_reg_513__2_ ( .D(n16515), .CP(wclk), .Q(ram[12274]) );
  DFF ram_reg_513__1_ ( .D(n16514), .CP(wclk), .Q(ram[12273]) );
  DFF ram_reg_513__0_ ( .D(n16513), .CP(wclk), .Q(ram[12272]) );
  DFF ram_reg_517__7_ ( .D(n16488), .CP(wclk), .Q(ram[12247]) );
  DFF ram_reg_517__6_ ( .D(n16487), .CP(wclk), .Q(ram[12246]) );
  DFF ram_reg_517__5_ ( .D(n16486), .CP(wclk), .Q(ram[12245]) );
  DFF ram_reg_517__4_ ( .D(n16485), .CP(wclk), .Q(ram[12244]) );
  DFF ram_reg_517__3_ ( .D(n16484), .CP(wclk), .Q(ram[12243]) );
  DFF ram_reg_517__2_ ( .D(n16483), .CP(wclk), .Q(ram[12242]) );
  DFF ram_reg_517__1_ ( .D(n16482), .CP(wclk), .Q(ram[12241]) );
  DFF ram_reg_517__0_ ( .D(n16481), .CP(wclk), .Q(ram[12240]) );
  DFF ram_reg_529__7_ ( .D(n16392), .CP(wclk), .Q(ram[12151]) );
  DFF ram_reg_529__6_ ( .D(n16391), .CP(wclk), .Q(ram[12150]) );
  DFF ram_reg_529__5_ ( .D(n16390), .CP(wclk), .Q(ram[12149]) );
  DFF ram_reg_529__4_ ( .D(n16389), .CP(wclk), .Q(ram[12148]) );
  DFF ram_reg_529__3_ ( .D(n16388), .CP(wclk), .Q(ram[12147]) );
  DFF ram_reg_529__2_ ( .D(n16387), .CP(wclk), .Q(ram[12146]) );
  DFF ram_reg_529__1_ ( .D(n16386), .CP(wclk), .Q(ram[12145]) );
  DFF ram_reg_529__0_ ( .D(n16385), .CP(wclk), .Q(ram[12144]) );
  DFF ram_reg_533__7_ ( .D(n16360), .CP(wclk), .Q(ram[12119]) );
  DFF ram_reg_533__6_ ( .D(n16359), .CP(wclk), .Q(ram[12118]) );
  DFF ram_reg_533__5_ ( .D(n16358), .CP(wclk), .Q(ram[12117]) );
  DFF ram_reg_533__4_ ( .D(n16357), .CP(wclk), .Q(ram[12116]) );
  DFF ram_reg_533__3_ ( .D(n16356), .CP(wclk), .Q(ram[12115]) );
  DFF ram_reg_533__2_ ( .D(n16355), .CP(wclk), .Q(ram[12114]) );
  DFF ram_reg_533__1_ ( .D(n16354), .CP(wclk), .Q(ram[12113]) );
  DFF ram_reg_533__0_ ( .D(n16353), .CP(wclk), .Q(ram[12112]) );
  DFF ram_reg_549__7_ ( .D(n16232), .CP(wclk), .Q(ram[11991]) );
  DFF ram_reg_549__6_ ( .D(n16231), .CP(wclk), .Q(ram[11990]) );
  DFF ram_reg_549__5_ ( .D(n16230), .CP(wclk), .Q(ram[11989]) );
  DFF ram_reg_549__4_ ( .D(n16229), .CP(wclk), .Q(ram[11988]) );
  DFF ram_reg_549__3_ ( .D(n16228), .CP(wclk), .Q(ram[11987]) );
  DFF ram_reg_549__2_ ( .D(n16227), .CP(wclk), .Q(ram[11986]) );
  DFF ram_reg_549__1_ ( .D(n16226), .CP(wclk), .Q(ram[11985]) );
  DFF ram_reg_549__0_ ( .D(n16225), .CP(wclk), .Q(ram[11984]) );
  DFF ram_reg_565__7_ ( .D(n16104), .CP(wclk), .Q(ram[11863]) );
  DFF ram_reg_565__6_ ( .D(n16103), .CP(wclk), .Q(ram[11862]) );
  DFF ram_reg_565__5_ ( .D(n16102), .CP(wclk), .Q(ram[11861]) );
  DFF ram_reg_565__4_ ( .D(n16101), .CP(wclk), .Q(ram[11860]) );
  DFF ram_reg_565__3_ ( .D(n16100), .CP(wclk), .Q(ram[11859]) );
  DFF ram_reg_565__2_ ( .D(n16099), .CP(wclk), .Q(ram[11858]) );
  DFF ram_reg_565__1_ ( .D(n16098), .CP(wclk), .Q(ram[11857]) );
  DFF ram_reg_565__0_ ( .D(n16097), .CP(wclk), .Q(ram[11856]) );
  DFF ram_reg_577__7_ ( .D(n16008), .CP(wclk), .Q(ram[11767]) );
  DFF ram_reg_577__6_ ( .D(n16007), .CP(wclk), .Q(ram[11766]) );
  DFF ram_reg_577__5_ ( .D(n16006), .CP(wclk), .Q(ram[11765]) );
  DFF ram_reg_577__4_ ( .D(n16005), .CP(wclk), .Q(ram[11764]) );
  DFF ram_reg_577__3_ ( .D(n16004), .CP(wclk), .Q(ram[11763]) );
  DFF ram_reg_577__2_ ( .D(n16003), .CP(wclk), .Q(ram[11762]) );
  DFF ram_reg_577__1_ ( .D(n16002), .CP(wclk), .Q(ram[11761]) );
  DFF ram_reg_577__0_ ( .D(n16001), .CP(wclk), .Q(ram[11760]) );
  DFF ram_reg_581__7_ ( .D(n15976), .CP(wclk), .Q(ram[11735]) );
  DFF ram_reg_581__6_ ( .D(n15975), .CP(wclk), .Q(ram[11734]) );
  DFF ram_reg_581__5_ ( .D(n15974), .CP(wclk), .Q(ram[11733]) );
  DFF ram_reg_581__4_ ( .D(n15973), .CP(wclk), .Q(ram[11732]) );
  DFF ram_reg_581__3_ ( .D(n15972), .CP(wclk), .Q(ram[11731]) );
  DFF ram_reg_581__2_ ( .D(n15971), .CP(wclk), .Q(ram[11730]) );
  DFF ram_reg_581__1_ ( .D(n15970), .CP(wclk), .Q(ram[11729]) );
  DFF ram_reg_581__0_ ( .D(n15969), .CP(wclk), .Q(ram[11728]) );
  DFF ram_reg_589__7_ ( .D(n15912), .CP(wclk), .Q(ram[11671]) );
  DFF ram_reg_589__6_ ( .D(n15911), .CP(wclk), .Q(ram[11670]) );
  DFF ram_reg_589__5_ ( .D(n15910), .CP(wclk), .Q(ram[11669]) );
  DFF ram_reg_589__4_ ( .D(n15909), .CP(wclk), .Q(ram[11668]) );
  DFF ram_reg_589__3_ ( .D(n15908), .CP(wclk), .Q(ram[11667]) );
  DFF ram_reg_589__2_ ( .D(n15907), .CP(wclk), .Q(ram[11666]) );
  DFF ram_reg_589__1_ ( .D(n15906), .CP(wclk), .Q(ram[11665]) );
  DFF ram_reg_589__0_ ( .D(n15905), .CP(wclk), .Q(ram[11664]) );
  DFF ram_reg_593__7_ ( .D(n15880), .CP(wclk), .Q(ram[11639]) );
  DFF ram_reg_593__6_ ( .D(n15879), .CP(wclk), .Q(ram[11638]) );
  DFF ram_reg_593__5_ ( .D(n15878), .CP(wclk), .Q(ram[11637]) );
  DFF ram_reg_593__4_ ( .D(n15877), .CP(wclk), .Q(ram[11636]) );
  DFF ram_reg_593__3_ ( .D(n15876), .CP(wclk), .Q(ram[11635]) );
  DFF ram_reg_593__2_ ( .D(n15875), .CP(wclk), .Q(ram[11634]) );
  DFF ram_reg_593__1_ ( .D(n15874), .CP(wclk), .Q(ram[11633]) );
  DFF ram_reg_593__0_ ( .D(n15873), .CP(wclk), .Q(ram[11632]) );
  DFF ram_reg_597__7_ ( .D(n15848), .CP(wclk), .Q(ram[11607]) );
  DFF ram_reg_597__6_ ( .D(n15847), .CP(wclk), .Q(ram[11606]) );
  DFF ram_reg_597__5_ ( .D(n15846), .CP(wclk), .Q(ram[11605]) );
  DFF ram_reg_597__4_ ( .D(n15845), .CP(wclk), .Q(ram[11604]) );
  DFF ram_reg_597__3_ ( .D(n15844), .CP(wclk), .Q(ram[11603]) );
  DFF ram_reg_597__2_ ( .D(n15843), .CP(wclk), .Q(ram[11602]) );
  DFF ram_reg_597__1_ ( .D(n15842), .CP(wclk), .Q(ram[11601]) );
  DFF ram_reg_597__0_ ( .D(n15841), .CP(wclk), .Q(ram[11600]) );
  DFF ram_reg_601__7_ ( .D(n15816), .CP(wclk), .Q(ram[11575]) );
  DFF ram_reg_601__6_ ( .D(n15815), .CP(wclk), .Q(ram[11574]) );
  DFF ram_reg_601__5_ ( .D(n15814), .CP(wclk), .Q(ram[11573]) );
  DFF ram_reg_601__4_ ( .D(n15813), .CP(wclk), .Q(ram[11572]) );
  DFF ram_reg_601__3_ ( .D(n15812), .CP(wclk), .Q(ram[11571]) );
  DFF ram_reg_601__2_ ( .D(n15811), .CP(wclk), .Q(ram[11570]) );
  DFF ram_reg_601__1_ ( .D(n15810), .CP(wclk), .Q(ram[11569]) );
  DFF ram_reg_601__0_ ( .D(n15809), .CP(wclk), .Q(ram[11568]) );
  DFF ram_reg_605__7_ ( .D(n15784), .CP(wclk), .Q(ram[11543]) );
  DFF ram_reg_605__6_ ( .D(n15783), .CP(wclk), .Q(ram[11542]) );
  DFF ram_reg_605__5_ ( .D(n15782), .CP(wclk), .Q(ram[11541]) );
  DFF ram_reg_605__4_ ( .D(n15781), .CP(wclk), .Q(ram[11540]) );
  DFF ram_reg_605__3_ ( .D(n15780), .CP(wclk), .Q(ram[11539]) );
  DFF ram_reg_605__2_ ( .D(n15779), .CP(wclk), .Q(ram[11538]) );
  DFF ram_reg_605__1_ ( .D(n15778), .CP(wclk), .Q(ram[11537]) );
  DFF ram_reg_605__0_ ( .D(n15777), .CP(wclk), .Q(ram[11536]) );
  DFF ram_reg_609__7_ ( .D(n15752), .CP(wclk), .Q(ram[11511]) );
  DFF ram_reg_609__6_ ( .D(n15751), .CP(wclk), .Q(ram[11510]) );
  DFF ram_reg_609__5_ ( .D(n15750), .CP(wclk), .Q(ram[11509]) );
  DFF ram_reg_609__4_ ( .D(n15749), .CP(wclk), .Q(ram[11508]) );
  DFF ram_reg_609__3_ ( .D(n15748), .CP(wclk), .Q(ram[11507]) );
  DFF ram_reg_609__2_ ( .D(n15747), .CP(wclk), .Q(ram[11506]) );
  DFF ram_reg_609__1_ ( .D(n15746), .CP(wclk), .Q(ram[11505]) );
  DFF ram_reg_609__0_ ( .D(n15745), .CP(wclk), .Q(ram[11504]) );
  DFF ram_reg_613__7_ ( .D(n15720), .CP(wclk), .Q(ram[11479]) );
  DFF ram_reg_613__6_ ( .D(n15719), .CP(wclk), .Q(ram[11478]) );
  DFF ram_reg_613__5_ ( .D(n15718), .CP(wclk), .Q(ram[11477]) );
  DFF ram_reg_613__4_ ( .D(n15717), .CP(wclk), .Q(ram[11476]) );
  DFF ram_reg_613__3_ ( .D(n15716), .CP(wclk), .Q(ram[11475]) );
  DFF ram_reg_613__2_ ( .D(n15715), .CP(wclk), .Q(ram[11474]) );
  DFF ram_reg_613__1_ ( .D(n15714), .CP(wclk), .Q(ram[11473]) );
  DFF ram_reg_613__0_ ( .D(n15713), .CP(wclk), .Q(ram[11472]) );
  DFF ram_reg_625__7_ ( .D(n15624), .CP(wclk), .Q(ram[11383]) );
  DFF ram_reg_625__6_ ( .D(n15623), .CP(wclk), .Q(ram[11382]) );
  DFF ram_reg_625__5_ ( .D(n15622), .CP(wclk), .Q(ram[11381]) );
  DFF ram_reg_625__4_ ( .D(n15621), .CP(wclk), .Q(ram[11380]) );
  DFF ram_reg_625__3_ ( .D(n15620), .CP(wclk), .Q(ram[11379]) );
  DFF ram_reg_625__2_ ( .D(n15619), .CP(wclk), .Q(ram[11378]) );
  DFF ram_reg_625__1_ ( .D(n15618), .CP(wclk), .Q(ram[11377]) );
  DFF ram_reg_625__0_ ( .D(n15617), .CP(wclk), .Q(ram[11376]) );
  DFF ram_reg_629__7_ ( .D(n15592), .CP(wclk), .Q(ram[11351]) );
  DFF ram_reg_629__6_ ( .D(n15591), .CP(wclk), .Q(ram[11350]) );
  DFF ram_reg_629__5_ ( .D(n15590), .CP(wclk), .Q(ram[11349]) );
  DFF ram_reg_629__4_ ( .D(n15589), .CP(wclk), .Q(ram[11348]) );
  DFF ram_reg_629__3_ ( .D(n15588), .CP(wclk), .Q(ram[11347]) );
  DFF ram_reg_629__2_ ( .D(n15587), .CP(wclk), .Q(ram[11346]) );
  DFF ram_reg_629__1_ ( .D(n15586), .CP(wclk), .Q(ram[11345]) );
  DFF ram_reg_629__0_ ( .D(n15585), .CP(wclk), .Q(ram[11344]) );
  DFF ram_reg_661__7_ ( .D(n15336), .CP(wclk), .Q(ram[11095]) );
  DFF ram_reg_661__6_ ( .D(n15335), .CP(wclk), .Q(ram[11094]) );
  DFF ram_reg_661__5_ ( .D(n15334), .CP(wclk), .Q(ram[11093]) );
  DFF ram_reg_661__4_ ( .D(n15333), .CP(wclk), .Q(ram[11092]) );
  DFF ram_reg_661__3_ ( .D(n15332), .CP(wclk), .Q(ram[11091]) );
  DFF ram_reg_661__2_ ( .D(n15331), .CP(wclk), .Q(ram[11090]) );
  DFF ram_reg_661__1_ ( .D(n15330), .CP(wclk), .Q(ram[11089]) );
  DFF ram_reg_661__0_ ( .D(n15329), .CP(wclk), .Q(ram[11088]) );
  DFF ram_reg_709__7_ ( .D(n14952), .CP(wclk), .Q(ram[10711]) );
  DFF ram_reg_709__6_ ( .D(n14951), .CP(wclk), .Q(ram[10710]) );
  DFF ram_reg_709__5_ ( .D(n14950), .CP(wclk), .Q(ram[10709]) );
  DFF ram_reg_709__4_ ( .D(n14949), .CP(wclk), .Q(ram[10708]) );
  DFF ram_reg_709__3_ ( .D(n14948), .CP(wclk), .Q(ram[10707]) );
  DFF ram_reg_709__2_ ( .D(n14947), .CP(wclk), .Q(ram[10706]) );
  DFF ram_reg_709__1_ ( .D(n14946), .CP(wclk), .Q(ram[10705]) );
  DFF ram_reg_709__0_ ( .D(n14945), .CP(wclk), .Q(ram[10704]) );
  DFF ram_reg_725__7_ ( .D(n14824), .CP(wclk), .Q(ram[10583]) );
  DFF ram_reg_725__6_ ( .D(n14823), .CP(wclk), .Q(ram[10582]) );
  DFF ram_reg_725__5_ ( .D(n14822), .CP(wclk), .Q(ram[10581]) );
  DFF ram_reg_725__4_ ( .D(n14821), .CP(wclk), .Q(ram[10580]) );
  DFF ram_reg_725__3_ ( .D(n14820), .CP(wclk), .Q(ram[10579]) );
  DFF ram_reg_725__2_ ( .D(n14819), .CP(wclk), .Q(ram[10578]) );
  DFF ram_reg_725__1_ ( .D(n14818), .CP(wclk), .Q(ram[10577]) );
  DFF ram_reg_725__0_ ( .D(n14817), .CP(wclk), .Q(ram[10576]) );
  DFF ram_reg_769__7_ ( .D(n14472), .CP(wclk), .Q(ram[10231]) );
  DFF ram_reg_769__6_ ( .D(n14471), .CP(wclk), .Q(ram[10230]) );
  DFF ram_reg_769__5_ ( .D(n14470), .CP(wclk), .Q(ram[10229]) );
  DFF ram_reg_769__4_ ( .D(n14469), .CP(wclk), .Q(ram[10228]) );
  DFF ram_reg_769__3_ ( .D(n14468), .CP(wclk), .Q(ram[10227]) );
  DFF ram_reg_769__2_ ( .D(n14467), .CP(wclk), .Q(ram[10226]) );
  DFF ram_reg_769__1_ ( .D(n14466), .CP(wclk), .Q(ram[10225]) );
  DFF ram_reg_769__0_ ( .D(n14465), .CP(wclk), .Q(ram[10224]) );
  DFF ram_reg_773__7_ ( .D(n14440), .CP(wclk), .Q(ram[10199]) );
  DFF ram_reg_773__6_ ( .D(n14439), .CP(wclk), .Q(ram[10198]) );
  DFF ram_reg_773__5_ ( .D(n14438), .CP(wclk), .Q(ram[10197]) );
  DFF ram_reg_773__4_ ( .D(n14437), .CP(wclk), .Q(ram[10196]) );
  DFF ram_reg_773__3_ ( .D(n14436), .CP(wclk), .Q(ram[10195]) );
  DFF ram_reg_773__2_ ( .D(n14435), .CP(wclk), .Q(ram[10194]) );
  DFF ram_reg_773__1_ ( .D(n14434), .CP(wclk), .Q(ram[10193]) );
  DFF ram_reg_773__0_ ( .D(n14433), .CP(wclk), .Q(ram[10192]) );
  DFF ram_reg_785__7_ ( .D(n14344), .CP(wclk), .Q(ram[10103]) );
  DFF ram_reg_785__6_ ( .D(n14343), .CP(wclk), .Q(ram[10102]) );
  DFF ram_reg_785__5_ ( .D(n14342), .CP(wclk), .Q(ram[10101]) );
  DFF ram_reg_785__4_ ( .D(n14341), .CP(wclk), .Q(ram[10100]) );
  DFF ram_reg_785__3_ ( .D(n14340), .CP(wclk), .Q(ram[10099]) );
  DFF ram_reg_785__2_ ( .D(n14339), .CP(wclk), .Q(ram[10098]) );
  DFF ram_reg_785__1_ ( .D(n14338), .CP(wclk), .Q(ram[10097]) );
  DFF ram_reg_785__0_ ( .D(n14337), .CP(wclk), .Q(ram[10096]) );
  DFF ram_reg_789__7_ ( .D(n14312), .CP(wclk), .Q(ram[10071]) );
  DFF ram_reg_789__6_ ( .D(n14311), .CP(wclk), .Q(ram[10070]) );
  DFF ram_reg_789__5_ ( .D(n14310), .CP(wclk), .Q(ram[10069]) );
  DFF ram_reg_789__4_ ( .D(n14309), .CP(wclk), .Q(ram[10068]) );
  DFF ram_reg_789__3_ ( .D(n14308), .CP(wclk), .Q(ram[10067]) );
  DFF ram_reg_789__2_ ( .D(n14307), .CP(wclk), .Q(ram[10066]) );
  DFF ram_reg_789__1_ ( .D(n14306), .CP(wclk), .Q(ram[10065]) );
  DFF ram_reg_789__0_ ( .D(n14305), .CP(wclk), .Q(ram[10064]) );
  DFF ram_reg_805__7_ ( .D(n14184), .CP(wclk), .Q(ram[9943]) );
  DFF ram_reg_805__6_ ( .D(n14183), .CP(wclk), .Q(ram[9942]) );
  DFF ram_reg_805__5_ ( .D(n14182), .CP(wclk), .Q(ram[9941]) );
  DFF ram_reg_805__4_ ( .D(n14181), .CP(wclk), .Q(ram[9940]) );
  DFF ram_reg_805__3_ ( .D(n14180), .CP(wclk), .Q(ram[9939]) );
  DFF ram_reg_805__2_ ( .D(n14179), .CP(wclk), .Q(ram[9938]) );
  DFF ram_reg_805__1_ ( .D(n14178), .CP(wclk), .Q(ram[9937]) );
  DFF ram_reg_805__0_ ( .D(n14177), .CP(wclk), .Q(ram[9936]) );
  DFF ram_reg_821__7_ ( .D(n14056), .CP(wclk), .Q(ram[9815]) );
  DFF ram_reg_821__6_ ( .D(n14055), .CP(wclk), .Q(ram[9814]) );
  DFF ram_reg_821__5_ ( .D(n14054), .CP(wclk), .Q(ram[9813]) );
  DFF ram_reg_821__4_ ( .D(n14053), .CP(wclk), .Q(ram[9812]) );
  DFF ram_reg_821__3_ ( .D(n14052), .CP(wclk), .Q(ram[9811]) );
  DFF ram_reg_821__2_ ( .D(n14051), .CP(wclk), .Q(ram[9810]) );
  DFF ram_reg_821__1_ ( .D(n14050), .CP(wclk), .Q(ram[9809]) );
  DFF ram_reg_821__0_ ( .D(n14049), .CP(wclk), .Q(ram[9808]) );
  DFF ram_reg_833__7_ ( .D(n13960), .CP(wclk), .Q(ram[9719]) );
  DFF ram_reg_833__6_ ( .D(n13959), .CP(wclk), .Q(ram[9718]) );
  DFF ram_reg_833__5_ ( .D(n13958), .CP(wclk), .Q(ram[9717]) );
  DFF ram_reg_833__4_ ( .D(n13957), .CP(wclk), .Q(ram[9716]) );
  DFF ram_reg_833__3_ ( .D(n13956), .CP(wclk), .Q(ram[9715]) );
  DFF ram_reg_833__2_ ( .D(n13955), .CP(wclk), .Q(ram[9714]) );
  DFF ram_reg_833__1_ ( .D(n13954), .CP(wclk), .Q(ram[9713]) );
  DFF ram_reg_833__0_ ( .D(n13953), .CP(wclk), .Q(ram[9712]) );
  DFF ram_reg_837__7_ ( .D(n13928), .CP(wclk), .Q(ram[9687]) );
  DFF ram_reg_837__6_ ( .D(n13927), .CP(wclk), .Q(ram[9686]) );
  DFF ram_reg_837__5_ ( .D(n13926), .CP(wclk), .Q(ram[9685]) );
  DFF ram_reg_837__4_ ( .D(n13925), .CP(wclk), .Q(ram[9684]) );
  DFF ram_reg_837__3_ ( .D(n13924), .CP(wclk), .Q(ram[9683]) );
  DFF ram_reg_837__2_ ( .D(n13923), .CP(wclk), .Q(ram[9682]) );
  DFF ram_reg_837__1_ ( .D(n13922), .CP(wclk), .Q(ram[9681]) );
  DFF ram_reg_837__0_ ( .D(n13921), .CP(wclk), .Q(ram[9680]) );
  DFF ram_reg_845__7_ ( .D(n13864), .CP(wclk), .Q(ram[9623]) );
  DFF ram_reg_845__6_ ( .D(n13863), .CP(wclk), .Q(ram[9622]) );
  DFF ram_reg_845__5_ ( .D(n13862), .CP(wclk), .Q(ram[9621]) );
  DFF ram_reg_845__4_ ( .D(n13861), .CP(wclk), .Q(ram[9620]) );
  DFF ram_reg_845__3_ ( .D(n13860), .CP(wclk), .Q(ram[9619]) );
  DFF ram_reg_845__2_ ( .D(n13859), .CP(wclk), .Q(ram[9618]) );
  DFF ram_reg_845__1_ ( .D(n13858), .CP(wclk), .Q(ram[9617]) );
  DFF ram_reg_845__0_ ( .D(n13857), .CP(wclk), .Q(ram[9616]) );
  DFF ram_reg_849__7_ ( .D(n13832), .CP(wclk), .Q(ram[9591]) );
  DFF ram_reg_849__6_ ( .D(n13831), .CP(wclk), .Q(ram[9590]) );
  DFF ram_reg_849__5_ ( .D(n13830), .CP(wclk), .Q(ram[9589]) );
  DFF ram_reg_849__4_ ( .D(n13829), .CP(wclk), .Q(ram[9588]) );
  DFF ram_reg_849__3_ ( .D(n13828), .CP(wclk), .Q(ram[9587]) );
  DFF ram_reg_849__2_ ( .D(n13827), .CP(wclk), .Q(ram[9586]) );
  DFF ram_reg_849__1_ ( .D(n13826), .CP(wclk), .Q(ram[9585]) );
  DFF ram_reg_849__0_ ( .D(n13825), .CP(wclk), .Q(ram[9584]) );
  DFF ram_reg_853__7_ ( .D(n13800), .CP(wclk), .Q(ram[9559]) );
  DFF ram_reg_853__6_ ( .D(n13799), .CP(wclk), .Q(ram[9558]) );
  DFF ram_reg_853__5_ ( .D(n13798), .CP(wclk), .Q(ram[9557]) );
  DFF ram_reg_853__4_ ( .D(n13797), .CP(wclk), .Q(ram[9556]) );
  DFF ram_reg_853__3_ ( .D(n13796), .CP(wclk), .Q(ram[9555]) );
  DFF ram_reg_853__2_ ( .D(n13795), .CP(wclk), .Q(ram[9554]) );
  DFF ram_reg_853__1_ ( .D(n13794), .CP(wclk), .Q(ram[9553]) );
  DFF ram_reg_853__0_ ( .D(n13793), .CP(wclk), .Q(ram[9552]) );
  DFF ram_reg_857__7_ ( .D(n13768), .CP(wclk), .Q(ram[9527]) );
  DFF ram_reg_857__6_ ( .D(n13767), .CP(wclk), .Q(ram[9526]) );
  DFF ram_reg_857__5_ ( .D(n13766), .CP(wclk), .Q(ram[9525]) );
  DFF ram_reg_857__4_ ( .D(n13765), .CP(wclk), .Q(ram[9524]) );
  DFF ram_reg_857__3_ ( .D(n13764), .CP(wclk), .Q(ram[9523]) );
  DFF ram_reg_857__2_ ( .D(n13763), .CP(wclk), .Q(ram[9522]) );
  DFF ram_reg_857__1_ ( .D(n13762), .CP(wclk), .Q(ram[9521]) );
  DFF ram_reg_857__0_ ( .D(n13761), .CP(wclk), .Q(ram[9520]) );
  DFF ram_reg_861__7_ ( .D(n13736), .CP(wclk), .Q(ram[9495]) );
  DFF ram_reg_861__6_ ( .D(n13735), .CP(wclk), .Q(ram[9494]) );
  DFF ram_reg_861__5_ ( .D(n13734), .CP(wclk), .Q(ram[9493]) );
  DFF ram_reg_861__4_ ( .D(n13733), .CP(wclk), .Q(ram[9492]) );
  DFF ram_reg_861__3_ ( .D(n13732), .CP(wclk), .Q(ram[9491]) );
  DFF ram_reg_861__2_ ( .D(n13731), .CP(wclk), .Q(ram[9490]) );
  DFF ram_reg_861__1_ ( .D(n13730), .CP(wclk), .Q(ram[9489]) );
  DFF ram_reg_861__0_ ( .D(n13729), .CP(wclk), .Q(ram[9488]) );
  DFF ram_reg_865__7_ ( .D(n13704), .CP(wclk), .Q(ram[9463]) );
  DFF ram_reg_865__6_ ( .D(n13703), .CP(wclk), .Q(ram[9462]) );
  DFF ram_reg_865__5_ ( .D(n13702), .CP(wclk), .Q(ram[9461]) );
  DFF ram_reg_865__4_ ( .D(n13701), .CP(wclk), .Q(ram[9460]) );
  DFF ram_reg_865__3_ ( .D(n13700), .CP(wclk), .Q(ram[9459]) );
  DFF ram_reg_865__2_ ( .D(n13699), .CP(wclk), .Q(ram[9458]) );
  DFF ram_reg_865__1_ ( .D(n13698), .CP(wclk), .Q(ram[9457]) );
  DFF ram_reg_865__0_ ( .D(n13697), .CP(wclk), .Q(ram[9456]) );
  DFF ram_reg_869__7_ ( .D(n13672), .CP(wclk), .Q(ram[9431]) );
  DFF ram_reg_869__6_ ( .D(n13671), .CP(wclk), .Q(ram[9430]) );
  DFF ram_reg_869__5_ ( .D(n13670), .CP(wclk), .Q(ram[9429]) );
  DFF ram_reg_869__4_ ( .D(n13669), .CP(wclk), .Q(ram[9428]) );
  DFF ram_reg_869__3_ ( .D(n13668), .CP(wclk), .Q(ram[9427]) );
  DFF ram_reg_869__2_ ( .D(n13667), .CP(wclk), .Q(ram[9426]) );
  DFF ram_reg_869__1_ ( .D(n13666), .CP(wclk), .Q(ram[9425]) );
  DFF ram_reg_869__0_ ( .D(n13665), .CP(wclk), .Q(ram[9424]) );
  DFF ram_reg_881__7_ ( .D(n13576), .CP(wclk), .Q(ram[9335]) );
  DFF ram_reg_881__6_ ( .D(n13575), .CP(wclk), .Q(ram[9334]) );
  DFF ram_reg_881__5_ ( .D(n13574), .CP(wclk), .Q(ram[9333]) );
  DFF ram_reg_881__4_ ( .D(n13573), .CP(wclk), .Q(ram[9332]) );
  DFF ram_reg_881__3_ ( .D(n13572), .CP(wclk), .Q(ram[9331]) );
  DFF ram_reg_881__2_ ( .D(n13571), .CP(wclk), .Q(ram[9330]) );
  DFF ram_reg_881__1_ ( .D(n13570), .CP(wclk), .Q(ram[9329]) );
  DFF ram_reg_881__0_ ( .D(n13569), .CP(wclk), .Q(ram[9328]) );
  DFF ram_reg_885__7_ ( .D(n13544), .CP(wclk), .Q(ram[9303]) );
  DFF ram_reg_885__6_ ( .D(n13543), .CP(wclk), .Q(ram[9302]) );
  DFF ram_reg_885__5_ ( .D(n13542), .CP(wclk), .Q(ram[9301]) );
  DFF ram_reg_885__4_ ( .D(n13541), .CP(wclk), .Q(ram[9300]) );
  DFF ram_reg_885__3_ ( .D(n13540), .CP(wclk), .Q(ram[9299]) );
  DFF ram_reg_885__2_ ( .D(n13539), .CP(wclk), .Q(ram[9298]) );
  DFF ram_reg_885__1_ ( .D(n13538), .CP(wclk), .Q(ram[9297]) );
  DFF ram_reg_885__0_ ( .D(n13537), .CP(wclk), .Q(ram[9296]) );
  DFF ram_reg_917__7_ ( .D(n13288), .CP(wclk), .Q(ram[9047]) );
  DFF ram_reg_917__6_ ( .D(n13287), .CP(wclk), .Q(ram[9046]) );
  DFF ram_reg_917__5_ ( .D(n13286), .CP(wclk), .Q(ram[9045]) );
  DFF ram_reg_917__4_ ( .D(n13285), .CP(wclk), .Q(ram[9044]) );
  DFF ram_reg_917__3_ ( .D(n13284), .CP(wclk), .Q(ram[9043]) );
  DFF ram_reg_917__2_ ( .D(n13283), .CP(wclk), .Q(ram[9042]) );
  DFF ram_reg_917__1_ ( .D(n13282), .CP(wclk), .Q(ram[9041]) );
  DFF ram_reg_917__0_ ( .D(n13281), .CP(wclk), .Q(ram[9040]) );
  DFF ram_reg_965__7_ ( .D(n12904), .CP(wclk), .Q(ram[8663]) );
  DFF ram_reg_965__6_ ( .D(n12903), .CP(wclk), .Q(ram[8662]) );
  DFF ram_reg_965__5_ ( .D(n12902), .CP(wclk), .Q(ram[8661]) );
  DFF ram_reg_965__4_ ( .D(n12901), .CP(wclk), .Q(ram[8660]) );
  DFF ram_reg_965__3_ ( .D(n12900), .CP(wclk), .Q(ram[8659]) );
  DFF ram_reg_965__2_ ( .D(n12899), .CP(wclk), .Q(ram[8658]) );
  DFF ram_reg_965__1_ ( .D(n12898), .CP(wclk), .Q(ram[8657]) );
  DFF ram_reg_965__0_ ( .D(n12897), .CP(wclk), .Q(ram[8656]) );
  DFF ram_reg_981__7_ ( .D(n12776), .CP(wclk), .Q(ram[8535]) );
  DFF ram_reg_981__6_ ( .D(n12775), .CP(wclk), .Q(ram[8534]) );
  DFF ram_reg_981__5_ ( .D(n12774), .CP(wclk), .Q(ram[8533]) );
  DFF ram_reg_981__4_ ( .D(n12773), .CP(wclk), .Q(ram[8532]) );
  DFF ram_reg_981__3_ ( .D(n12772), .CP(wclk), .Q(ram[8531]) );
  DFF ram_reg_981__2_ ( .D(n12771), .CP(wclk), .Q(ram[8530]) );
  DFF ram_reg_981__1_ ( .D(n12770), .CP(wclk), .Q(ram[8529]) );
  DFF ram_reg_981__0_ ( .D(n12769), .CP(wclk), .Q(ram[8528]) );
  DFF ram_reg_1025__7_ ( .D(n12424), .CP(wclk), .Q(ram[8183]) );
  DFF ram_reg_1025__6_ ( .D(n12423), .CP(wclk), .Q(ram[8182]) );
  DFF ram_reg_1025__5_ ( .D(n12422), .CP(wclk), .Q(ram[8181]) );
  DFF ram_reg_1025__4_ ( .D(n12421), .CP(wclk), .Q(ram[8180]) );
  DFF ram_reg_1025__3_ ( .D(n12420), .CP(wclk), .Q(ram[8179]) );
  DFF ram_reg_1025__2_ ( .D(n12419), .CP(wclk), .Q(ram[8178]) );
  DFF ram_reg_1025__1_ ( .D(n12418), .CP(wclk), .Q(ram[8177]) );
  DFF ram_reg_1025__0_ ( .D(n12417), .CP(wclk), .Q(ram[8176]) );
  DFF ram_reg_1029__7_ ( .D(n12392), .CP(wclk), .Q(ram[8151]) );
  DFF ram_reg_1029__6_ ( .D(n12391), .CP(wclk), .Q(ram[8150]) );
  DFF ram_reg_1029__5_ ( .D(n12390), .CP(wclk), .Q(ram[8149]) );
  DFF ram_reg_1029__4_ ( .D(n12389), .CP(wclk), .Q(ram[8148]) );
  DFF ram_reg_1029__3_ ( .D(n12388), .CP(wclk), .Q(ram[8147]) );
  DFF ram_reg_1029__2_ ( .D(n12387), .CP(wclk), .Q(ram[8146]) );
  DFF ram_reg_1029__1_ ( .D(n12386), .CP(wclk), .Q(ram[8145]) );
  DFF ram_reg_1029__0_ ( .D(n12385), .CP(wclk), .Q(ram[8144]) );
  DFF ram_reg_1041__7_ ( .D(n12296), .CP(wclk), .Q(ram[8055]) );
  DFF ram_reg_1041__6_ ( .D(n12295), .CP(wclk), .Q(ram[8054]) );
  DFF ram_reg_1041__5_ ( .D(n12294), .CP(wclk), .Q(ram[8053]) );
  DFF ram_reg_1041__4_ ( .D(n12293), .CP(wclk), .Q(ram[8052]) );
  DFF ram_reg_1041__3_ ( .D(n12292), .CP(wclk), .Q(ram[8051]) );
  DFF ram_reg_1041__2_ ( .D(n12291), .CP(wclk), .Q(ram[8050]) );
  DFF ram_reg_1041__1_ ( .D(n12290), .CP(wclk), .Q(ram[8049]) );
  DFF ram_reg_1041__0_ ( .D(n12289), .CP(wclk), .Q(ram[8048]) );
  DFF ram_reg_1045__7_ ( .D(n12264), .CP(wclk), .Q(ram[8023]) );
  DFF ram_reg_1045__6_ ( .D(n12263), .CP(wclk), .Q(ram[8022]) );
  DFF ram_reg_1045__5_ ( .D(n12262), .CP(wclk), .Q(ram[8021]) );
  DFF ram_reg_1045__4_ ( .D(n12261), .CP(wclk), .Q(ram[8020]) );
  DFF ram_reg_1045__3_ ( .D(n12260), .CP(wclk), .Q(ram[8019]) );
  DFF ram_reg_1045__2_ ( .D(n12259), .CP(wclk), .Q(ram[8018]) );
  DFF ram_reg_1045__1_ ( .D(n12258), .CP(wclk), .Q(ram[8017]) );
  DFF ram_reg_1045__0_ ( .D(n12257), .CP(wclk), .Q(ram[8016]) );
  DFF ram_reg_1053__7_ ( .D(n12200), .CP(wclk), .Q(ram[7959]) );
  DFF ram_reg_1053__6_ ( .D(n12199), .CP(wclk), .Q(ram[7958]) );
  DFF ram_reg_1053__5_ ( .D(n12198), .CP(wclk), .Q(ram[7957]) );
  DFF ram_reg_1053__4_ ( .D(n12197), .CP(wclk), .Q(ram[7956]) );
  DFF ram_reg_1053__3_ ( .D(n12196), .CP(wclk), .Q(ram[7955]) );
  DFF ram_reg_1053__2_ ( .D(n12195), .CP(wclk), .Q(ram[7954]) );
  DFF ram_reg_1053__1_ ( .D(n12194), .CP(wclk), .Q(ram[7953]) );
  DFF ram_reg_1053__0_ ( .D(n12193), .CP(wclk), .Q(ram[7952]) );
  DFF ram_reg_1057__7_ ( .D(n12168), .CP(wclk), .Q(ram[7927]) );
  DFF ram_reg_1057__6_ ( .D(n12167), .CP(wclk), .Q(ram[7926]) );
  DFF ram_reg_1057__5_ ( .D(n12166), .CP(wclk), .Q(ram[7925]) );
  DFF ram_reg_1057__4_ ( .D(n12165), .CP(wclk), .Q(ram[7924]) );
  DFF ram_reg_1057__3_ ( .D(n12164), .CP(wclk), .Q(ram[7923]) );
  DFF ram_reg_1057__2_ ( .D(n12163), .CP(wclk), .Q(ram[7922]) );
  DFF ram_reg_1057__1_ ( .D(n12162), .CP(wclk), .Q(ram[7921]) );
  DFF ram_reg_1057__0_ ( .D(n12161), .CP(wclk), .Q(ram[7920]) );
  DFF ram_reg_1061__7_ ( .D(n12136), .CP(wclk), .Q(ram[7895]) );
  DFF ram_reg_1061__6_ ( .D(n12135), .CP(wclk), .Q(ram[7894]) );
  DFF ram_reg_1061__5_ ( .D(n12134), .CP(wclk), .Q(ram[7893]) );
  DFF ram_reg_1061__4_ ( .D(n12133), .CP(wclk), .Q(ram[7892]) );
  DFF ram_reg_1061__3_ ( .D(n12132), .CP(wclk), .Q(ram[7891]) );
  DFF ram_reg_1061__2_ ( .D(n12131), .CP(wclk), .Q(ram[7890]) );
  DFF ram_reg_1061__1_ ( .D(n12130), .CP(wclk), .Q(ram[7889]) );
  DFF ram_reg_1061__0_ ( .D(n12129), .CP(wclk), .Q(ram[7888]) );
  DFF ram_reg_1077__7_ ( .D(n12008), .CP(wclk), .Q(ram[7767]) );
  DFF ram_reg_1077__6_ ( .D(n12007), .CP(wclk), .Q(ram[7766]) );
  DFF ram_reg_1077__5_ ( .D(n12006), .CP(wclk), .Q(ram[7765]) );
  DFF ram_reg_1077__4_ ( .D(n12005), .CP(wclk), .Q(ram[7764]) );
  DFF ram_reg_1077__3_ ( .D(n12004), .CP(wclk), .Q(ram[7763]) );
  DFF ram_reg_1077__2_ ( .D(n12003), .CP(wclk), .Q(ram[7762]) );
  DFF ram_reg_1077__1_ ( .D(n12002), .CP(wclk), .Q(ram[7761]) );
  DFF ram_reg_1077__0_ ( .D(n12001), .CP(wclk), .Q(ram[7760]) );
  DFF ram_reg_1089__7_ ( .D(n11912), .CP(wclk), .Q(ram[7671]) );
  DFF ram_reg_1089__6_ ( .D(n11911), .CP(wclk), .Q(ram[7670]) );
  DFF ram_reg_1089__5_ ( .D(n11910), .CP(wclk), .Q(ram[7669]) );
  DFF ram_reg_1089__4_ ( .D(n11909), .CP(wclk), .Q(ram[7668]) );
  DFF ram_reg_1089__3_ ( .D(n11908), .CP(wclk), .Q(ram[7667]) );
  DFF ram_reg_1089__2_ ( .D(n11907), .CP(wclk), .Q(ram[7666]) );
  DFF ram_reg_1089__1_ ( .D(n11906), .CP(wclk), .Q(ram[7665]) );
  DFF ram_reg_1089__0_ ( .D(n11905), .CP(wclk), .Q(ram[7664]) );
  DFF ram_reg_1093__7_ ( .D(n11880), .CP(wclk), .Q(ram[7639]) );
  DFF ram_reg_1093__6_ ( .D(n11879), .CP(wclk), .Q(ram[7638]) );
  DFF ram_reg_1093__5_ ( .D(n11878), .CP(wclk), .Q(ram[7637]) );
  DFF ram_reg_1093__4_ ( .D(n11877), .CP(wclk), .Q(ram[7636]) );
  DFF ram_reg_1093__3_ ( .D(n11876), .CP(wclk), .Q(ram[7635]) );
  DFF ram_reg_1093__2_ ( .D(n11875), .CP(wclk), .Q(ram[7634]) );
  DFF ram_reg_1093__1_ ( .D(n11874), .CP(wclk), .Q(ram[7633]) );
  DFF ram_reg_1093__0_ ( .D(n11873), .CP(wclk), .Q(ram[7632]) );
  DFF ram_reg_1097__7_ ( .D(n11848), .CP(wclk), .Q(ram[7607]) );
  DFF ram_reg_1097__6_ ( .D(n11847), .CP(wclk), .Q(ram[7606]) );
  DFF ram_reg_1097__5_ ( .D(n11846), .CP(wclk), .Q(ram[7605]) );
  DFF ram_reg_1097__4_ ( .D(n11845), .CP(wclk), .Q(ram[7604]) );
  DFF ram_reg_1097__3_ ( .D(n11844), .CP(wclk), .Q(ram[7603]) );
  DFF ram_reg_1097__2_ ( .D(n11843), .CP(wclk), .Q(ram[7602]) );
  DFF ram_reg_1097__1_ ( .D(n11842), .CP(wclk), .Q(ram[7601]) );
  DFF ram_reg_1097__0_ ( .D(n11841), .CP(wclk), .Q(ram[7600]) );
  DFF ram_reg_1101__7_ ( .D(n11816), .CP(wclk), .Q(ram[7575]) );
  DFF ram_reg_1101__6_ ( .D(n11815), .CP(wclk), .Q(ram[7574]) );
  DFF ram_reg_1101__5_ ( .D(n11814), .CP(wclk), .Q(ram[7573]) );
  DFF ram_reg_1101__4_ ( .D(n11813), .CP(wclk), .Q(ram[7572]) );
  DFF ram_reg_1101__3_ ( .D(n11812), .CP(wclk), .Q(ram[7571]) );
  DFF ram_reg_1101__2_ ( .D(n11811), .CP(wclk), .Q(ram[7570]) );
  DFF ram_reg_1101__1_ ( .D(n11810), .CP(wclk), .Q(ram[7569]) );
  DFF ram_reg_1101__0_ ( .D(n11809), .CP(wclk), .Q(ram[7568]) );
  DFF ram_reg_1105__7_ ( .D(n11784), .CP(wclk), .Q(ram[7543]) );
  DFF ram_reg_1105__6_ ( .D(n11783), .CP(wclk), .Q(ram[7542]) );
  DFF ram_reg_1105__5_ ( .D(n11782), .CP(wclk), .Q(ram[7541]) );
  DFF ram_reg_1105__4_ ( .D(n11781), .CP(wclk), .Q(ram[7540]) );
  DFF ram_reg_1105__3_ ( .D(n11780), .CP(wclk), .Q(ram[7539]) );
  DFF ram_reg_1105__2_ ( .D(n11779), .CP(wclk), .Q(ram[7538]) );
  DFF ram_reg_1105__1_ ( .D(n11778), .CP(wclk), .Q(ram[7537]) );
  DFF ram_reg_1105__0_ ( .D(n11777), .CP(wclk), .Q(ram[7536]) );
  DFF ram_reg_1109__7_ ( .D(n11752), .CP(wclk), .Q(ram[7511]) );
  DFF ram_reg_1109__6_ ( .D(n11751), .CP(wclk), .Q(ram[7510]) );
  DFF ram_reg_1109__5_ ( .D(n11750), .CP(wclk), .Q(ram[7509]) );
  DFF ram_reg_1109__4_ ( .D(n11749), .CP(wclk), .Q(ram[7508]) );
  DFF ram_reg_1109__3_ ( .D(n11748), .CP(wclk), .Q(ram[7507]) );
  DFF ram_reg_1109__2_ ( .D(n11747), .CP(wclk), .Q(ram[7506]) );
  DFF ram_reg_1109__1_ ( .D(n11746), .CP(wclk), .Q(ram[7505]) );
  DFF ram_reg_1109__0_ ( .D(n11745), .CP(wclk), .Q(ram[7504]) );
  DFF ram_reg_1113__7_ ( .D(n11720), .CP(wclk), .Q(ram[7479]) );
  DFF ram_reg_1113__6_ ( .D(n11719), .CP(wclk), .Q(ram[7478]) );
  DFF ram_reg_1113__5_ ( .D(n11718), .CP(wclk), .Q(ram[7477]) );
  DFF ram_reg_1113__4_ ( .D(n11717), .CP(wclk), .Q(ram[7476]) );
  DFF ram_reg_1113__3_ ( .D(n11716), .CP(wclk), .Q(ram[7475]) );
  DFF ram_reg_1113__2_ ( .D(n11715), .CP(wclk), .Q(ram[7474]) );
  DFF ram_reg_1113__1_ ( .D(n11714), .CP(wclk), .Q(ram[7473]) );
  DFF ram_reg_1113__0_ ( .D(n11713), .CP(wclk), .Q(ram[7472]) );
  DFF ram_reg_1117__7_ ( .D(n11688), .CP(wclk), .Q(ram[7447]) );
  DFF ram_reg_1117__6_ ( .D(n11687), .CP(wclk), .Q(ram[7446]) );
  DFF ram_reg_1117__5_ ( .D(n11686), .CP(wclk), .Q(ram[7445]) );
  DFF ram_reg_1117__4_ ( .D(n11685), .CP(wclk), .Q(ram[7444]) );
  DFF ram_reg_1117__3_ ( .D(n11684), .CP(wclk), .Q(ram[7443]) );
  DFF ram_reg_1117__2_ ( .D(n11683), .CP(wclk), .Q(ram[7442]) );
  DFF ram_reg_1117__1_ ( .D(n11682), .CP(wclk), .Q(ram[7441]) );
  DFF ram_reg_1117__0_ ( .D(n11681), .CP(wclk), .Q(ram[7440]) );
  DFF ram_reg_1121__7_ ( .D(n11656), .CP(wclk), .Q(ram[7415]) );
  DFF ram_reg_1121__6_ ( .D(n11655), .CP(wclk), .Q(ram[7414]) );
  DFF ram_reg_1121__5_ ( .D(n11654), .CP(wclk), .Q(ram[7413]) );
  DFF ram_reg_1121__4_ ( .D(n11653), .CP(wclk), .Q(ram[7412]) );
  DFF ram_reg_1121__3_ ( .D(n11652), .CP(wclk), .Q(ram[7411]) );
  DFF ram_reg_1121__2_ ( .D(n11651), .CP(wclk), .Q(ram[7410]) );
  DFF ram_reg_1121__1_ ( .D(n11650), .CP(wclk), .Q(ram[7409]) );
  DFF ram_reg_1121__0_ ( .D(n11649), .CP(wclk), .Q(ram[7408]) );
  DFF ram_reg_1125__7_ ( .D(n11624), .CP(wclk), .Q(ram[7383]) );
  DFF ram_reg_1125__6_ ( .D(n11623), .CP(wclk), .Q(ram[7382]) );
  DFF ram_reg_1125__5_ ( .D(n11622), .CP(wclk), .Q(ram[7381]) );
  DFF ram_reg_1125__4_ ( .D(n11621), .CP(wclk), .Q(ram[7380]) );
  DFF ram_reg_1125__3_ ( .D(n11620), .CP(wclk), .Q(ram[7379]) );
  DFF ram_reg_1125__2_ ( .D(n11619), .CP(wclk), .Q(ram[7378]) );
  DFF ram_reg_1125__1_ ( .D(n11618), .CP(wclk), .Q(ram[7377]) );
  DFF ram_reg_1125__0_ ( .D(n11617), .CP(wclk), .Q(ram[7376]) );
  DFF ram_reg_1133__7_ ( .D(n11560), .CP(wclk), .Q(ram[7319]) );
  DFF ram_reg_1133__6_ ( .D(n11559), .CP(wclk), .Q(ram[7318]) );
  DFF ram_reg_1133__5_ ( .D(n11558), .CP(wclk), .Q(ram[7317]) );
  DFF ram_reg_1133__4_ ( .D(n11557), .CP(wclk), .Q(ram[7316]) );
  DFF ram_reg_1133__3_ ( .D(n11556), .CP(wclk), .Q(ram[7315]) );
  DFF ram_reg_1133__2_ ( .D(n11555), .CP(wclk), .Q(ram[7314]) );
  DFF ram_reg_1133__1_ ( .D(n11554), .CP(wclk), .Q(ram[7313]) );
  DFF ram_reg_1133__0_ ( .D(n11553), .CP(wclk), .Q(ram[7312]) );
  DFF ram_reg_1137__7_ ( .D(n11528), .CP(wclk), .Q(ram[7287]) );
  DFF ram_reg_1137__6_ ( .D(n11527), .CP(wclk), .Q(ram[7286]) );
  DFF ram_reg_1137__5_ ( .D(n11526), .CP(wclk), .Q(ram[7285]) );
  DFF ram_reg_1137__4_ ( .D(n11525), .CP(wclk), .Q(ram[7284]) );
  DFF ram_reg_1137__3_ ( .D(n11524), .CP(wclk), .Q(ram[7283]) );
  DFF ram_reg_1137__2_ ( .D(n11523), .CP(wclk), .Q(ram[7282]) );
  DFF ram_reg_1137__1_ ( .D(n11522), .CP(wclk), .Q(ram[7281]) );
  DFF ram_reg_1137__0_ ( .D(n11521), .CP(wclk), .Q(ram[7280]) );
  DFF ram_reg_1141__7_ ( .D(n11496), .CP(wclk), .Q(ram[7255]) );
  DFF ram_reg_1141__6_ ( .D(n11495), .CP(wclk), .Q(ram[7254]) );
  DFF ram_reg_1141__5_ ( .D(n11494), .CP(wclk), .Q(ram[7253]) );
  DFF ram_reg_1141__4_ ( .D(n11493), .CP(wclk), .Q(ram[7252]) );
  DFF ram_reg_1141__3_ ( .D(n11492), .CP(wclk), .Q(ram[7251]) );
  DFF ram_reg_1141__2_ ( .D(n11491), .CP(wclk), .Q(ram[7250]) );
  DFF ram_reg_1141__1_ ( .D(n11490), .CP(wclk), .Q(ram[7249]) );
  DFF ram_reg_1141__0_ ( .D(n11489), .CP(wclk), .Q(ram[7248]) );
  DFF ram_reg_1149__7_ ( .D(n11432), .CP(wclk), .Q(ram[7191]) );
  DFF ram_reg_1149__6_ ( .D(n11431), .CP(wclk), .Q(ram[7190]) );
  DFF ram_reg_1149__5_ ( .D(n11430), .CP(wclk), .Q(ram[7189]) );
  DFF ram_reg_1149__4_ ( .D(n11429), .CP(wclk), .Q(ram[7188]) );
  DFF ram_reg_1149__3_ ( .D(n11428), .CP(wclk), .Q(ram[7187]) );
  DFF ram_reg_1149__2_ ( .D(n11427), .CP(wclk), .Q(ram[7186]) );
  DFF ram_reg_1149__1_ ( .D(n11426), .CP(wclk), .Q(ram[7185]) );
  DFF ram_reg_1149__0_ ( .D(n11425), .CP(wclk), .Q(ram[7184]) );
  DFF ram_reg_1157__7_ ( .D(n11368), .CP(wclk), .Q(ram[7127]) );
  DFF ram_reg_1157__6_ ( .D(n11367), .CP(wclk), .Q(ram[7126]) );
  DFF ram_reg_1157__5_ ( .D(n11366), .CP(wclk), .Q(ram[7125]) );
  DFF ram_reg_1157__4_ ( .D(n11365), .CP(wclk), .Q(ram[7124]) );
  DFF ram_reg_1157__3_ ( .D(n11364), .CP(wclk), .Q(ram[7123]) );
  DFF ram_reg_1157__2_ ( .D(n11363), .CP(wclk), .Q(ram[7122]) );
  DFF ram_reg_1157__1_ ( .D(n11362), .CP(wclk), .Q(ram[7121]) );
  DFF ram_reg_1157__0_ ( .D(n11361), .CP(wclk), .Q(ram[7120]) );
  DFF ram_reg_1173__7_ ( .D(n11240), .CP(wclk), .Q(ram[6999]) );
  DFF ram_reg_1173__6_ ( .D(n11239), .CP(wclk), .Q(ram[6998]) );
  DFF ram_reg_1173__5_ ( .D(n11238), .CP(wclk), .Q(ram[6997]) );
  DFF ram_reg_1173__4_ ( .D(n11237), .CP(wclk), .Q(ram[6996]) );
  DFF ram_reg_1173__3_ ( .D(n11236), .CP(wclk), .Q(ram[6995]) );
  DFF ram_reg_1173__2_ ( .D(n11235), .CP(wclk), .Q(ram[6994]) );
  DFF ram_reg_1173__1_ ( .D(n11234), .CP(wclk), .Q(ram[6993]) );
  DFF ram_reg_1173__0_ ( .D(n11233), .CP(wclk), .Q(ram[6992]) );
  DFF ram_reg_1221__7_ ( .D(n10856), .CP(wclk), .Q(ram[6615]) );
  DFF ram_reg_1221__6_ ( .D(n10855), .CP(wclk), .Q(ram[6614]) );
  DFF ram_reg_1221__5_ ( .D(n10854), .CP(wclk), .Q(ram[6613]) );
  DFF ram_reg_1221__4_ ( .D(n10853), .CP(wclk), .Q(ram[6612]) );
  DFF ram_reg_1221__3_ ( .D(n10852), .CP(wclk), .Q(ram[6611]) );
  DFF ram_reg_1221__2_ ( .D(n10851), .CP(wclk), .Q(ram[6610]) );
  DFF ram_reg_1221__1_ ( .D(n10850), .CP(wclk), .Q(ram[6609]) );
  DFF ram_reg_1221__0_ ( .D(n10849), .CP(wclk), .Q(ram[6608]) );
  DFF ram_reg_1233__7_ ( .D(n10760), .CP(wclk), .Q(ram[6519]) );
  DFF ram_reg_1233__6_ ( .D(n10759), .CP(wclk), .Q(ram[6518]) );
  DFF ram_reg_1233__5_ ( .D(n10758), .CP(wclk), .Q(ram[6517]) );
  DFF ram_reg_1233__4_ ( .D(n10757), .CP(wclk), .Q(ram[6516]) );
  DFF ram_reg_1233__3_ ( .D(n10756), .CP(wclk), .Q(ram[6515]) );
  DFF ram_reg_1233__2_ ( .D(n10755), .CP(wclk), .Q(ram[6514]) );
  DFF ram_reg_1233__1_ ( .D(n10754), .CP(wclk), .Q(ram[6513]) );
  DFF ram_reg_1233__0_ ( .D(n10753), .CP(wclk), .Q(ram[6512]) );
  DFF ram_reg_1237__7_ ( .D(n10728), .CP(wclk), .Q(ram[6487]) );
  DFF ram_reg_1237__6_ ( .D(n10727), .CP(wclk), .Q(ram[6486]) );
  DFF ram_reg_1237__5_ ( .D(n10726), .CP(wclk), .Q(ram[6485]) );
  DFF ram_reg_1237__4_ ( .D(n10725), .CP(wclk), .Q(ram[6484]) );
  DFF ram_reg_1237__3_ ( .D(n10724), .CP(wclk), .Q(ram[6483]) );
  DFF ram_reg_1237__2_ ( .D(n10723), .CP(wclk), .Q(ram[6482]) );
  DFF ram_reg_1237__1_ ( .D(n10722), .CP(wclk), .Q(ram[6481]) );
  DFF ram_reg_1237__0_ ( .D(n10721), .CP(wclk), .Q(ram[6480]) );
  DFF ram_reg_1253__7_ ( .D(n10600), .CP(wclk), .Q(ram[6359]) );
  DFF ram_reg_1253__6_ ( .D(n10599), .CP(wclk), .Q(ram[6358]) );
  DFF ram_reg_1253__5_ ( .D(n10598), .CP(wclk), .Q(ram[6357]) );
  DFF ram_reg_1253__4_ ( .D(n10597), .CP(wclk), .Q(ram[6356]) );
  DFF ram_reg_1253__3_ ( .D(n10596), .CP(wclk), .Q(ram[6355]) );
  DFF ram_reg_1253__2_ ( .D(n10595), .CP(wclk), .Q(ram[6354]) );
  DFF ram_reg_1253__1_ ( .D(n10594), .CP(wclk), .Q(ram[6353]) );
  DFF ram_reg_1253__0_ ( .D(n10593), .CP(wclk), .Q(ram[6352]) );
  DFF ram_reg_1269__7_ ( .D(n10472), .CP(wclk), .Q(ram[6231]) );
  DFF ram_reg_1269__6_ ( .D(n10471), .CP(wclk), .Q(ram[6230]) );
  DFF ram_reg_1269__5_ ( .D(n10470), .CP(wclk), .Q(ram[6229]) );
  DFF ram_reg_1269__4_ ( .D(n10469), .CP(wclk), .Q(ram[6228]) );
  DFF ram_reg_1269__3_ ( .D(n10468), .CP(wclk), .Q(ram[6227]) );
  DFF ram_reg_1269__2_ ( .D(n10467), .CP(wclk), .Q(ram[6226]) );
  DFF ram_reg_1269__1_ ( .D(n10466), .CP(wclk), .Q(ram[6225]) );
  DFF ram_reg_1269__0_ ( .D(n10465), .CP(wclk), .Q(ram[6224]) );
  DFF ram_reg_1285__7_ ( .D(n10344), .CP(wclk), .Q(ram[6103]) );
  DFF ram_reg_1285__6_ ( .D(n10343), .CP(wclk), .Q(ram[6102]) );
  DFF ram_reg_1285__5_ ( .D(n10342), .CP(wclk), .Q(ram[6101]) );
  DFF ram_reg_1285__4_ ( .D(n10341), .CP(wclk), .Q(ram[6100]) );
  DFF ram_reg_1285__3_ ( .D(n10340), .CP(wclk), .Q(ram[6099]) );
  DFF ram_reg_1285__2_ ( .D(n10339), .CP(wclk), .Q(ram[6098]) );
  DFF ram_reg_1285__1_ ( .D(n10338), .CP(wclk), .Q(ram[6097]) );
  DFF ram_reg_1285__0_ ( .D(n10337), .CP(wclk), .Q(ram[6096]) );
  DFF ram_reg_1297__7_ ( .D(n10248), .CP(wclk), .Q(ram[6007]) );
  DFF ram_reg_1297__6_ ( .D(n10247), .CP(wclk), .Q(ram[6006]) );
  DFF ram_reg_1297__5_ ( .D(n10246), .CP(wclk), .Q(ram[6005]) );
  DFF ram_reg_1297__4_ ( .D(n10245), .CP(wclk), .Q(ram[6004]) );
  DFF ram_reg_1297__3_ ( .D(n10244), .CP(wclk), .Q(ram[6003]) );
  DFF ram_reg_1297__2_ ( .D(n10243), .CP(wclk), .Q(ram[6002]) );
  DFF ram_reg_1297__1_ ( .D(n10242), .CP(wclk), .Q(ram[6001]) );
  DFF ram_reg_1297__0_ ( .D(n10241), .CP(wclk), .Q(ram[6000]) );
  DFF ram_reg_1301__7_ ( .D(n10216), .CP(wclk), .Q(ram[5975]) );
  DFF ram_reg_1301__6_ ( .D(n10215), .CP(wclk), .Q(ram[5974]) );
  DFF ram_reg_1301__5_ ( .D(n10214), .CP(wclk), .Q(ram[5973]) );
  DFF ram_reg_1301__4_ ( .D(n10213), .CP(wclk), .Q(ram[5972]) );
  DFF ram_reg_1301__3_ ( .D(n10212), .CP(wclk), .Q(ram[5971]) );
  DFF ram_reg_1301__2_ ( .D(n10211), .CP(wclk), .Q(ram[5970]) );
  DFF ram_reg_1301__1_ ( .D(n10210), .CP(wclk), .Q(ram[5969]) );
  DFF ram_reg_1301__0_ ( .D(n10209), .CP(wclk), .Q(ram[5968]) );
  DFF ram_reg_1317__7_ ( .D(n10088), .CP(wclk), .Q(ram[5847]) );
  DFF ram_reg_1317__6_ ( .D(n10087), .CP(wclk), .Q(ram[5846]) );
  DFF ram_reg_1317__5_ ( .D(n10086), .CP(wclk), .Q(ram[5845]) );
  DFF ram_reg_1317__4_ ( .D(n10085), .CP(wclk), .Q(ram[5844]) );
  DFF ram_reg_1317__3_ ( .D(n10084), .CP(wclk), .Q(ram[5843]) );
  DFF ram_reg_1317__2_ ( .D(n10083), .CP(wclk), .Q(ram[5842]) );
  DFF ram_reg_1317__1_ ( .D(n10082), .CP(wclk), .Q(ram[5841]) );
  DFF ram_reg_1317__0_ ( .D(n10081), .CP(wclk), .Q(ram[5840]) );
  DFF ram_reg_1333__7_ ( .D(n9960), .CP(wclk), .Q(ram[5719]) );
  DFF ram_reg_1333__6_ ( .D(n9959), .CP(wclk), .Q(ram[5718]) );
  DFF ram_reg_1333__5_ ( .D(n9958), .CP(wclk), .Q(ram[5717]) );
  DFF ram_reg_1333__4_ ( .D(n9957), .CP(wclk), .Q(ram[5716]) );
  DFF ram_reg_1333__3_ ( .D(n9956), .CP(wclk), .Q(ram[5715]) );
  DFF ram_reg_1333__2_ ( .D(n9955), .CP(wclk), .Q(ram[5714]) );
  DFF ram_reg_1333__1_ ( .D(n9954), .CP(wclk), .Q(ram[5713]) );
  DFF ram_reg_1333__0_ ( .D(n9953), .CP(wclk), .Q(ram[5712]) );
  DFF ram_reg_1345__7_ ( .D(n9864), .CP(wclk), .Q(ram[5623]) );
  DFF ram_reg_1345__6_ ( .D(n9863), .CP(wclk), .Q(ram[5622]) );
  DFF ram_reg_1345__5_ ( .D(n9862), .CP(wclk), .Q(ram[5621]) );
  DFF ram_reg_1345__4_ ( .D(n9861), .CP(wclk), .Q(ram[5620]) );
  DFF ram_reg_1345__3_ ( .D(n9860), .CP(wclk), .Q(ram[5619]) );
  DFF ram_reg_1345__2_ ( .D(n9859), .CP(wclk), .Q(ram[5618]) );
  DFF ram_reg_1345__1_ ( .D(n9858), .CP(wclk), .Q(ram[5617]) );
  DFF ram_reg_1345__0_ ( .D(n9857), .CP(wclk), .Q(ram[5616]) );
  DFF ram_reg_1349__7_ ( .D(n9832), .CP(wclk), .Q(ram[5591]) );
  DFF ram_reg_1349__6_ ( .D(n9831), .CP(wclk), .Q(ram[5590]) );
  DFF ram_reg_1349__5_ ( .D(n9830), .CP(wclk), .Q(ram[5589]) );
  DFF ram_reg_1349__4_ ( .D(n9829), .CP(wclk), .Q(ram[5588]) );
  DFF ram_reg_1349__3_ ( .D(n9828), .CP(wclk), .Q(ram[5587]) );
  DFF ram_reg_1349__2_ ( .D(n9827), .CP(wclk), .Q(ram[5586]) );
  DFF ram_reg_1349__1_ ( .D(n9826), .CP(wclk), .Q(ram[5585]) );
  DFF ram_reg_1349__0_ ( .D(n9825), .CP(wclk), .Q(ram[5584]) );
  DFF ram_reg_1361__7_ ( .D(n9736), .CP(wclk), .Q(ram[5495]) );
  DFF ram_reg_1361__6_ ( .D(n9735), .CP(wclk), .Q(ram[5494]) );
  DFF ram_reg_1361__5_ ( .D(n9734), .CP(wclk), .Q(ram[5493]) );
  DFF ram_reg_1361__4_ ( .D(n9733), .CP(wclk), .Q(ram[5492]) );
  DFF ram_reg_1361__3_ ( .D(n9732), .CP(wclk), .Q(ram[5491]) );
  DFF ram_reg_1361__2_ ( .D(n9731), .CP(wclk), .Q(ram[5490]) );
  DFF ram_reg_1361__1_ ( .D(n9730), .CP(wclk), .Q(ram[5489]) );
  DFF ram_reg_1361__0_ ( .D(n9729), .CP(wclk), .Q(ram[5488]) );
  DFF ram_reg_1365__7_ ( .D(n9704), .CP(wclk), .Q(ram[5463]) );
  DFF ram_reg_1365__6_ ( .D(n9703), .CP(wclk), .Q(ram[5462]) );
  DFF ram_reg_1365__5_ ( .D(n9702), .CP(wclk), .Q(ram[5461]) );
  DFF ram_reg_1365__4_ ( .D(n9701), .CP(wclk), .Q(ram[5460]) );
  DFF ram_reg_1365__3_ ( .D(n9700), .CP(wclk), .Q(ram[5459]) );
  DFF ram_reg_1365__2_ ( .D(n9699), .CP(wclk), .Q(ram[5458]) );
  DFF ram_reg_1365__1_ ( .D(n9698), .CP(wclk), .Q(ram[5457]) );
  DFF ram_reg_1365__0_ ( .D(n9697), .CP(wclk), .Q(ram[5456]) );
  DFF ram_reg_1373__7_ ( .D(n9640), .CP(wclk), .Q(ram[5399]) );
  DFF ram_reg_1373__6_ ( .D(n9639), .CP(wclk), .Q(ram[5398]) );
  DFF ram_reg_1373__5_ ( .D(n9638), .CP(wclk), .Q(ram[5397]) );
  DFF ram_reg_1373__4_ ( .D(n9637), .CP(wclk), .Q(ram[5396]) );
  DFF ram_reg_1373__3_ ( .D(n9636), .CP(wclk), .Q(ram[5395]) );
  DFF ram_reg_1373__2_ ( .D(n9635), .CP(wclk), .Q(ram[5394]) );
  DFF ram_reg_1373__1_ ( .D(n9634), .CP(wclk), .Q(ram[5393]) );
  DFF ram_reg_1373__0_ ( .D(n9633), .CP(wclk), .Q(ram[5392]) );
  DFF ram_reg_1377__7_ ( .D(n9608), .CP(wclk), .Q(ram[5367]) );
  DFF ram_reg_1377__6_ ( .D(n9607), .CP(wclk), .Q(ram[5366]) );
  DFF ram_reg_1377__5_ ( .D(n9606), .CP(wclk), .Q(ram[5365]) );
  DFF ram_reg_1377__4_ ( .D(n9605), .CP(wclk), .Q(ram[5364]) );
  DFF ram_reg_1377__3_ ( .D(n9604), .CP(wclk), .Q(ram[5363]) );
  DFF ram_reg_1377__2_ ( .D(n9603), .CP(wclk), .Q(ram[5362]) );
  DFF ram_reg_1377__1_ ( .D(n9602), .CP(wclk), .Q(ram[5361]) );
  DFF ram_reg_1377__0_ ( .D(n9601), .CP(wclk), .Q(ram[5360]) );
  DFF ram_reg_1381__7_ ( .D(n9576), .CP(wclk), .Q(ram[5335]) );
  DFF ram_reg_1381__6_ ( .D(n9575), .CP(wclk), .Q(ram[5334]) );
  DFF ram_reg_1381__5_ ( .D(n9574), .CP(wclk), .Q(ram[5333]) );
  DFF ram_reg_1381__4_ ( .D(n9573), .CP(wclk), .Q(ram[5332]) );
  DFF ram_reg_1381__3_ ( .D(n9572), .CP(wclk), .Q(ram[5331]) );
  DFF ram_reg_1381__2_ ( .D(n9571), .CP(wclk), .Q(ram[5330]) );
  DFF ram_reg_1381__1_ ( .D(n9570), .CP(wclk), .Q(ram[5329]) );
  DFF ram_reg_1381__0_ ( .D(n9569), .CP(wclk), .Q(ram[5328]) );
  DFF ram_reg_1393__7_ ( .D(n9480), .CP(wclk), .Q(ram[5239]) );
  DFF ram_reg_1393__6_ ( .D(n9479), .CP(wclk), .Q(ram[5238]) );
  DFF ram_reg_1393__5_ ( .D(n9478), .CP(wclk), .Q(ram[5237]) );
  DFF ram_reg_1393__4_ ( .D(n9477), .CP(wclk), .Q(ram[5236]) );
  DFF ram_reg_1393__3_ ( .D(n9476), .CP(wclk), .Q(ram[5235]) );
  DFF ram_reg_1393__2_ ( .D(n9475), .CP(wclk), .Q(ram[5234]) );
  DFF ram_reg_1393__1_ ( .D(n9474), .CP(wclk), .Q(ram[5233]) );
  DFF ram_reg_1393__0_ ( .D(n9473), .CP(wclk), .Q(ram[5232]) );
  DFF ram_reg_1397__7_ ( .D(n9448), .CP(wclk), .Q(ram[5207]) );
  DFF ram_reg_1397__6_ ( .D(n9447), .CP(wclk), .Q(ram[5206]) );
  DFF ram_reg_1397__5_ ( .D(n9446), .CP(wclk), .Q(ram[5205]) );
  DFF ram_reg_1397__4_ ( .D(n9445), .CP(wclk), .Q(ram[5204]) );
  DFF ram_reg_1397__3_ ( .D(n9444), .CP(wclk), .Q(ram[5203]) );
  DFF ram_reg_1397__2_ ( .D(n9443), .CP(wclk), .Q(ram[5202]) );
  DFF ram_reg_1397__1_ ( .D(n9442), .CP(wclk), .Q(ram[5201]) );
  DFF ram_reg_1397__0_ ( .D(n9441), .CP(wclk), .Q(ram[5200]) );
  DFF ram_reg_1493__7_ ( .D(n8680), .CP(wclk), .Q(ram[4439]) );
  DFF ram_reg_1493__6_ ( .D(n8679), .CP(wclk), .Q(ram[4438]) );
  DFF ram_reg_1493__5_ ( .D(n8678), .CP(wclk), .Q(ram[4437]) );
  DFF ram_reg_1493__4_ ( .D(n8677), .CP(wclk), .Q(ram[4436]) );
  DFF ram_reg_1493__3_ ( .D(n8676), .CP(wclk), .Q(ram[4435]) );
  DFF ram_reg_1493__2_ ( .D(n8675), .CP(wclk), .Q(ram[4434]) );
  DFF ram_reg_1493__1_ ( .D(n8674), .CP(wclk), .Q(ram[4433]) );
  DFF ram_reg_1493__0_ ( .D(n8673), .CP(wclk), .Q(ram[4432]) );
  DFF ram_reg_1537__7_ ( .D(n8328), .CP(wclk), .Q(ram[4087]) );
  DFF ram_reg_1537__6_ ( .D(n8327), .CP(wclk), .Q(ram[4086]) );
  DFF ram_reg_1537__5_ ( .D(n8326), .CP(wclk), .Q(ram[4085]) );
  DFF ram_reg_1537__4_ ( .D(n8325), .CP(wclk), .Q(ram[4084]) );
  DFF ram_reg_1537__3_ ( .D(n8324), .CP(wclk), .Q(ram[4083]) );
  DFF ram_reg_1537__2_ ( .D(n8323), .CP(wclk), .Q(ram[4082]) );
  DFF ram_reg_1537__1_ ( .D(n8322), .CP(wclk), .Q(ram[4081]) );
  DFF ram_reg_1537__0_ ( .D(n8321), .CP(wclk), .Q(ram[4080]) );
  DFF ram_reg_1541__7_ ( .D(n8296), .CP(wclk), .Q(ram[4055]) );
  DFF ram_reg_1541__6_ ( .D(n8295), .CP(wclk), .Q(ram[4054]) );
  DFF ram_reg_1541__5_ ( .D(n8294), .CP(wclk), .Q(ram[4053]) );
  DFF ram_reg_1541__4_ ( .D(n8293), .CP(wclk), .Q(ram[4052]) );
  DFF ram_reg_1541__3_ ( .D(n8292), .CP(wclk), .Q(ram[4051]) );
  DFF ram_reg_1541__2_ ( .D(n8291), .CP(wclk), .Q(ram[4050]) );
  DFF ram_reg_1541__1_ ( .D(n8290), .CP(wclk), .Q(ram[4049]) );
  DFF ram_reg_1541__0_ ( .D(n8289), .CP(wclk), .Q(ram[4048]) );
  DFF ram_reg_1553__7_ ( .D(n8200), .CP(wclk), .Q(ram[3959]) );
  DFF ram_reg_1553__6_ ( .D(n8199), .CP(wclk), .Q(ram[3958]) );
  DFF ram_reg_1553__5_ ( .D(n8198), .CP(wclk), .Q(ram[3957]) );
  DFF ram_reg_1553__4_ ( .D(n8197), .CP(wclk), .Q(ram[3956]) );
  DFF ram_reg_1553__3_ ( .D(n8196), .CP(wclk), .Q(ram[3955]) );
  DFF ram_reg_1553__2_ ( .D(n8195), .CP(wclk), .Q(ram[3954]) );
  DFF ram_reg_1553__1_ ( .D(n8194), .CP(wclk), .Q(ram[3953]) );
  DFF ram_reg_1553__0_ ( .D(n8193), .CP(wclk), .Q(ram[3952]) );
  DFF ram_reg_1557__7_ ( .D(n8168), .CP(wclk), .Q(ram[3927]) );
  DFF ram_reg_1557__6_ ( .D(n8167), .CP(wclk), .Q(ram[3926]) );
  DFF ram_reg_1557__5_ ( .D(n8166), .CP(wclk), .Q(ram[3925]) );
  DFF ram_reg_1557__4_ ( .D(n8165), .CP(wclk), .Q(ram[3924]) );
  DFF ram_reg_1557__3_ ( .D(n8164), .CP(wclk), .Q(ram[3923]) );
  DFF ram_reg_1557__2_ ( .D(n8163), .CP(wclk), .Q(ram[3922]) );
  DFF ram_reg_1557__1_ ( .D(n8162), .CP(wclk), .Q(ram[3921]) );
  DFF ram_reg_1557__0_ ( .D(n8161), .CP(wclk), .Q(ram[3920]) );
  DFF ram_reg_1565__7_ ( .D(n8104), .CP(wclk), .Q(ram[3863]) );
  DFF ram_reg_1565__6_ ( .D(n8103), .CP(wclk), .Q(ram[3862]) );
  DFF ram_reg_1565__5_ ( .D(n8102), .CP(wclk), .Q(ram[3861]) );
  DFF ram_reg_1565__4_ ( .D(n8101), .CP(wclk), .Q(ram[3860]) );
  DFF ram_reg_1565__3_ ( .D(n8100), .CP(wclk), .Q(ram[3859]) );
  DFF ram_reg_1565__2_ ( .D(n8099), .CP(wclk), .Q(ram[3858]) );
  DFF ram_reg_1565__1_ ( .D(n8098), .CP(wclk), .Q(ram[3857]) );
  DFF ram_reg_1565__0_ ( .D(n8097), .CP(wclk), .Q(ram[3856]) );
  DFF ram_reg_1569__7_ ( .D(n8072), .CP(wclk), .Q(ram[3831]) );
  DFF ram_reg_1569__6_ ( .D(n8071), .CP(wclk), .Q(ram[3830]) );
  DFF ram_reg_1569__5_ ( .D(n8070), .CP(wclk), .Q(ram[3829]) );
  DFF ram_reg_1569__4_ ( .D(n8069), .CP(wclk), .Q(ram[3828]) );
  DFF ram_reg_1569__3_ ( .D(n8068), .CP(wclk), .Q(ram[3827]) );
  DFF ram_reg_1569__2_ ( .D(n8067), .CP(wclk), .Q(ram[3826]) );
  DFF ram_reg_1569__1_ ( .D(n8066), .CP(wclk), .Q(ram[3825]) );
  DFF ram_reg_1569__0_ ( .D(n8065), .CP(wclk), .Q(ram[3824]) );
  DFF ram_reg_1573__7_ ( .D(n8040), .CP(wclk), .Q(ram[3799]) );
  DFF ram_reg_1573__6_ ( .D(n8039), .CP(wclk), .Q(ram[3798]) );
  DFF ram_reg_1573__5_ ( .D(n8038), .CP(wclk), .Q(ram[3797]) );
  DFF ram_reg_1573__4_ ( .D(n8037), .CP(wclk), .Q(ram[3796]) );
  DFF ram_reg_1573__3_ ( .D(n8036), .CP(wclk), .Q(ram[3795]) );
  DFF ram_reg_1573__2_ ( .D(n8035), .CP(wclk), .Q(ram[3794]) );
  DFF ram_reg_1573__1_ ( .D(n8034), .CP(wclk), .Q(ram[3793]) );
  DFF ram_reg_1573__0_ ( .D(n8033), .CP(wclk), .Q(ram[3792]) );
  DFF ram_reg_1589__7_ ( .D(n7912), .CP(wclk), .Q(ram[3671]) );
  DFF ram_reg_1589__6_ ( .D(n7911), .CP(wclk), .Q(ram[3670]) );
  DFF ram_reg_1589__5_ ( .D(n7910), .CP(wclk), .Q(ram[3669]) );
  DFF ram_reg_1589__4_ ( .D(n7909), .CP(wclk), .Q(ram[3668]) );
  DFF ram_reg_1589__3_ ( .D(n7908), .CP(wclk), .Q(ram[3667]) );
  DFF ram_reg_1589__2_ ( .D(n7907), .CP(wclk), .Q(ram[3666]) );
  DFF ram_reg_1589__1_ ( .D(n7906), .CP(wclk), .Q(ram[3665]) );
  DFF ram_reg_1589__0_ ( .D(n7905), .CP(wclk), .Q(ram[3664]) );
  DFF ram_reg_1601__7_ ( .D(n7816), .CP(wclk), .Q(ram[3575]) );
  DFF ram_reg_1601__6_ ( .D(n7815), .CP(wclk), .Q(ram[3574]) );
  DFF ram_reg_1601__5_ ( .D(n7814), .CP(wclk), .Q(ram[3573]) );
  DFF ram_reg_1601__4_ ( .D(n7813), .CP(wclk), .Q(ram[3572]) );
  DFF ram_reg_1601__3_ ( .D(n7812), .CP(wclk), .Q(ram[3571]) );
  DFF ram_reg_1601__2_ ( .D(n7811), .CP(wclk), .Q(ram[3570]) );
  DFF ram_reg_1601__1_ ( .D(n7810), .CP(wclk), .Q(ram[3569]) );
  DFF ram_reg_1601__0_ ( .D(n7809), .CP(wclk), .Q(ram[3568]) );
  DFF ram_reg_1605__7_ ( .D(n7784), .CP(wclk), .Q(ram[3543]) );
  DFF ram_reg_1605__6_ ( .D(n7783), .CP(wclk), .Q(ram[3542]) );
  DFF ram_reg_1605__5_ ( .D(n7782), .CP(wclk), .Q(ram[3541]) );
  DFF ram_reg_1605__4_ ( .D(n7781), .CP(wclk), .Q(ram[3540]) );
  DFF ram_reg_1605__3_ ( .D(n7780), .CP(wclk), .Q(ram[3539]) );
  DFF ram_reg_1605__2_ ( .D(n7779), .CP(wclk), .Q(ram[3538]) );
  DFF ram_reg_1605__1_ ( .D(n7778), .CP(wclk), .Q(ram[3537]) );
  DFF ram_reg_1605__0_ ( .D(n7777), .CP(wclk), .Q(ram[3536]) );
  DFF ram_reg_1609__7_ ( .D(n7752), .CP(wclk), .Q(ram[3511]) );
  DFF ram_reg_1609__6_ ( .D(n7751), .CP(wclk), .Q(ram[3510]) );
  DFF ram_reg_1609__5_ ( .D(n7750), .CP(wclk), .Q(ram[3509]) );
  DFF ram_reg_1609__4_ ( .D(n7749), .CP(wclk), .Q(ram[3508]) );
  DFF ram_reg_1609__3_ ( .D(n7748), .CP(wclk), .Q(ram[3507]) );
  DFF ram_reg_1609__2_ ( .D(n7747), .CP(wclk), .Q(ram[3506]) );
  DFF ram_reg_1609__1_ ( .D(n7746), .CP(wclk), .Q(ram[3505]) );
  DFF ram_reg_1609__0_ ( .D(n7745), .CP(wclk), .Q(ram[3504]) );
  DFF ram_reg_1613__7_ ( .D(n7720), .CP(wclk), .Q(ram[3479]) );
  DFF ram_reg_1613__6_ ( .D(n7719), .CP(wclk), .Q(ram[3478]) );
  DFF ram_reg_1613__5_ ( .D(n7718), .CP(wclk), .Q(ram[3477]) );
  DFF ram_reg_1613__4_ ( .D(n7717), .CP(wclk), .Q(ram[3476]) );
  DFF ram_reg_1613__3_ ( .D(n7716), .CP(wclk), .Q(ram[3475]) );
  DFF ram_reg_1613__2_ ( .D(n7715), .CP(wclk), .Q(ram[3474]) );
  DFF ram_reg_1613__1_ ( .D(n7714), .CP(wclk), .Q(ram[3473]) );
  DFF ram_reg_1613__0_ ( .D(n7713), .CP(wclk), .Q(ram[3472]) );
  DFF ram_reg_1617__7_ ( .D(n7688), .CP(wclk), .Q(ram[3447]) );
  DFF ram_reg_1617__6_ ( .D(n7687), .CP(wclk), .Q(ram[3446]) );
  DFF ram_reg_1617__5_ ( .D(n7686), .CP(wclk), .Q(ram[3445]) );
  DFF ram_reg_1617__4_ ( .D(n7685), .CP(wclk), .Q(ram[3444]) );
  DFF ram_reg_1617__3_ ( .D(n7684), .CP(wclk), .Q(ram[3443]) );
  DFF ram_reg_1617__2_ ( .D(n7683), .CP(wclk), .Q(ram[3442]) );
  DFF ram_reg_1617__1_ ( .D(n7682), .CP(wclk), .Q(ram[3441]) );
  DFF ram_reg_1617__0_ ( .D(n7681), .CP(wclk), .Q(ram[3440]) );
  DFF ram_reg_1621__7_ ( .D(n7656), .CP(wclk), .Q(ram[3415]) );
  DFF ram_reg_1621__6_ ( .D(n7655), .CP(wclk), .Q(ram[3414]) );
  DFF ram_reg_1621__5_ ( .D(n7654), .CP(wclk), .Q(ram[3413]) );
  DFF ram_reg_1621__4_ ( .D(n7653), .CP(wclk), .Q(ram[3412]) );
  DFF ram_reg_1621__3_ ( .D(n7652), .CP(wclk), .Q(ram[3411]) );
  DFF ram_reg_1621__2_ ( .D(n7651), .CP(wclk), .Q(ram[3410]) );
  DFF ram_reg_1621__1_ ( .D(n7650), .CP(wclk), .Q(ram[3409]) );
  DFF ram_reg_1621__0_ ( .D(n7649), .CP(wclk), .Q(ram[3408]) );
  DFF ram_reg_1625__7_ ( .D(n7624), .CP(wclk), .Q(ram[3383]) );
  DFF ram_reg_1625__6_ ( .D(n7623), .CP(wclk), .Q(ram[3382]) );
  DFF ram_reg_1625__5_ ( .D(n7622), .CP(wclk), .Q(ram[3381]) );
  DFF ram_reg_1625__4_ ( .D(n7621), .CP(wclk), .Q(ram[3380]) );
  DFF ram_reg_1625__3_ ( .D(n7620), .CP(wclk), .Q(ram[3379]) );
  DFF ram_reg_1625__2_ ( .D(n7619), .CP(wclk), .Q(ram[3378]) );
  DFF ram_reg_1625__1_ ( .D(n7618), .CP(wclk), .Q(ram[3377]) );
  DFF ram_reg_1625__0_ ( .D(n7617), .CP(wclk), .Q(ram[3376]) );
  DFF ram_reg_1629__7_ ( .D(n7592), .CP(wclk), .Q(ram[3351]) );
  DFF ram_reg_1629__6_ ( .D(n7591), .CP(wclk), .Q(ram[3350]) );
  DFF ram_reg_1629__5_ ( .D(n7590), .CP(wclk), .Q(ram[3349]) );
  DFF ram_reg_1629__4_ ( .D(n7589), .CP(wclk), .Q(ram[3348]) );
  DFF ram_reg_1629__3_ ( .D(n7588), .CP(wclk), .Q(ram[3347]) );
  DFF ram_reg_1629__2_ ( .D(n7587), .CP(wclk), .Q(ram[3346]) );
  DFF ram_reg_1629__1_ ( .D(n7586), .CP(wclk), .Q(ram[3345]) );
  DFF ram_reg_1629__0_ ( .D(n7585), .CP(wclk), .Q(ram[3344]) );
  DFF ram_reg_1633__7_ ( .D(n7560), .CP(wclk), .Q(ram[3319]) );
  DFF ram_reg_1633__6_ ( .D(n7559), .CP(wclk), .Q(ram[3318]) );
  DFF ram_reg_1633__5_ ( .D(n7558), .CP(wclk), .Q(ram[3317]) );
  DFF ram_reg_1633__4_ ( .D(n7557), .CP(wclk), .Q(ram[3316]) );
  DFF ram_reg_1633__3_ ( .D(n7556), .CP(wclk), .Q(ram[3315]) );
  DFF ram_reg_1633__2_ ( .D(n7555), .CP(wclk), .Q(ram[3314]) );
  DFF ram_reg_1633__1_ ( .D(n7554), .CP(wclk), .Q(ram[3313]) );
  DFF ram_reg_1633__0_ ( .D(n7553), .CP(wclk), .Q(ram[3312]) );
  DFF ram_reg_1637__7_ ( .D(n7528), .CP(wclk), .Q(ram[3287]) );
  DFF ram_reg_1637__6_ ( .D(n7527), .CP(wclk), .Q(ram[3286]) );
  DFF ram_reg_1637__5_ ( .D(n7526), .CP(wclk), .Q(ram[3285]) );
  DFF ram_reg_1637__4_ ( .D(n7525), .CP(wclk), .Q(ram[3284]) );
  DFF ram_reg_1637__3_ ( .D(n7524), .CP(wclk), .Q(ram[3283]) );
  DFF ram_reg_1637__2_ ( .D(n7523), .CP(wclk), .Q(ram[3282]) );
  DFF ram_reg_1637__1_ ( .D(n7522), .CP(wclk), .Q(ram[3281]) );
  DFF ram_reg_1637__0_ ( .D(n7521), .CP(wclk), .Q(ram[3280]) );
  DFF ram_reg_1645__7_ ( .D(n7464), .CP(wclk), .Q(ram[3223]) );
  DFF ram_reg_1645__6_ ( .D(n7463), .CP(wclk), .Q(ram[3222]) );
  DFF ram_reg_1645__5_ ( .D(n7462), .CP(wclk), .Q(ram[3221]) );
  DFF ram_reg_1645__4_ ( .D(n7461), .CP(wclk), .Q(ram[3220]) );
  DFF ram_reg_1645__3_ ( .D(n7460), .CP(wclk), .Q(ram[3219]) );
  DFF ram_reg_1645__2_ ( .D(n7459), .CP(wclk), .Q(ram[3218]) );
  DFF ram_reg_1645__1_ ( .D(n7458), .CP(wclk), .Q(ram[3217]) );
  DFF ram_reg_1645__0_ ( .D(n7457), .CP(wclk), .Q(ram[3216]) );
  DFF ram_reg_1649__7_ ( .D(n7432), .CP(wclk), .Q(ram[3191]) );
  DFF ram_reg_1649__6_ ( .D(n7431), .CP(wclk), .Q(ram[3190]) );
  DFF ram_reg_1649__5_ ( .D(n7430), .CP(wclk), .Q(ram[3189]) );
  DFF ram_reg_1649__4_ ( .D(n7429), .CP(wclk), .Q(ram[3188]) );
  DFF ram_reg_1649__3_ ( .D(n7428), .CP(wclk), .Q(ram[3187]) );
  DFF ram_reg_1649__2_ ( .D(n7427), .CP(wclk), .Q(ram[3186]) );
  DFF ram_reg_1649__1_ ( .D(n7426), .CP(wclk), .Q(ram[3185]) );
  DFF ram_reg_1649__0_ ( .D(n7425), .CP(wclk), .Q(ram[3184]) );
  DFF ram_reg_1653__7_ ( .D(n7400), .CP(wclk), .Q(ram[3159]) );
  DFF ram_reg_1653__6_ ( .D(n7399), .CP(wclk), .Q(ram[3158]) );
  DFF ram_reg_1653__5_ ( .D(n7398), .CP(wclk), .Q(ram[3157]) );
  DFF ram_reg_1653__4_ ( .D(n7397), .CP(wclk), .Q(ram[3156]) );
  DFF ram_reg_1653__3_ ( .D(n7396), .CP(wclk), .Q(ram[3155]) );
  DFF ram_reg_1653__2_ ( .D(n7395), .CP(wclk), .Q(ram[3154]) );
  DFF ram_reg_1653__1_ ( .D(n7394), .CP(wclk), .Q(ram[3153]) );
  DFF ram_reg_1653__0_ ( .D(n7393), .CP(wclk), .Q(ram[3152]) );
  DFF ram_reg_1661__7_ ( .D(n7336), .CP(wclk), .Q(ram[3095]) );
  DFF ram_reg_1661__6_ ( .D(n7335), .CP(wclk), .Q(ram[3094]) );
  DFF ram_reg_1661__5_ ( .D(n7334), .CP(wclk), .Q(ram[3093]) );
  DFF ram_reg_1661__4_ ( .D(n7333), .CP(wclk), .Q(ram[3092]) );
  DFF ram_reg_1661__3_ ( .D(n7332), .CP(wclk), .Q(ram[3091]) );
  DFF ram_reg_1661__2_ ( .D(n7331), .CP(wclk), .Q(ram[3090]) );
  DFF ram_reg_1661__1_ ( .D(n7330), .CP(wclk), .Q(ram[3089]) );
  DFF ram_reg_1661__0_ ( .D(n7329), .CP(wclk), .Q(ram[3088]) );
  DFF ram_reg_1669__7_ ( .D(n7272), .CP(wclk), .Q(ram[3031]) );
  DFF ram_reg_1669__6_ ( .D(n7271), .CP(wclk), .Q(ram[3030]) );
  DFF ram_reg_1669__5_ ( .D(n7270), .CP(wclk), .Q(ram[3029]) );
  DFF ram_reg_1669__4_ ( .D(n7269), .CP(wclk), .Q(ram[3028]) );
  DFF ram_reg_1669__3_ ( .D(n7268), .CP(wclk), .Q(ram[3027]) );
  DFF ram_reg_1669__2_ ( .D(n7267), .CP(wclk), .Q(ram[3026]) );
  DFF ram_reg_1669__1_ ( .D(n7266), .CP(wclk), .Q(ram[3025]) );
  DFF ram_reg_1669__0_ ( .D(n7265), .CP(wclk), .Q(ram[3024]) );
  DFF ram_reg_1685__7_ ( .D(n7144), .CP(wclk), .Q(ram[2903]) );
  DFF ram_reg_1685__6_ ( .D(n7143), .CP(wclk), .Q(ram[2902]) );
  DFF ram_reg_1685__5_ ( .D(n7142), .CP(wclk), .Q(ram[2901]) );
  DFF ram_reg_1685__4_ ( .D(n7141), .CP(wclk), .Q(ram[2900]) );
  DFF ram_reg_1685__3_ ( .D(n7140), .CP(wclk), .Q(ram[2899]) );
  DFF ram_reg_1685__2_ ( .D(n7139), .CP(wclk), .Q(ram[2898]) );
  DFF ram_reg_1685__1_ ( .D(n7138), .CP(wclk), .Q(ram[2897]) );
  DFF ram_reg_1685__0_ ( .D(n7137), .CP(wclk), .Q(ram[2896]) );
  DFF ram_reg_1733__7_ ( .D(n6760), .CP(wclk), .Q(ram[2519]) );
  DFF ram_reg_1733__6_ ( .D(n6759), .CP(wclk), .Q(ram[2518]) );
  DFF ram_reg_1733__5_ ( .D(n6758), .CP(wclk), .Q(ram[2517]) );
  DFF ram_reg_1733__4_ ( .D(n6757), .CP(wclk), .Q(ram[2516]) );
  DFF ram_reg_1733__3_ ( .D(n6756), .CP(wclk), .Q(ram[2515]) );
  DFF ram_reg_1733__2_ ( .D(n6755), .CP(wclk), .Q(ram[2514]) );
  DFF ram_reg_1733__1_ ( .D(n6754), .CP(wclk), .Q(ram[2513]) );
  DFF ram_reg_1733__0_ ( .D(n6753), .CP(wclk), .Q(ram[2512]) );
  DFF ram_reg_1745__7_ ( .D(n6664), .CP(wclk), .Q(ram[2423]) );
  DFF ram_reg_1745__6_ ( .D(n6663), .CP(wclk), .Q(ram[2422]) );
  DFF ram_reg_1745__5_ ( .D(n6662), .CP(wclk), .Q(ram[2421]) );
  DFF ram_reg_1745__4_ ( .D(n6661), .CP(wclk), .Q(ram[2420]) );
  DFF ram_reg_1745__3_ ( .D(n6660), .CP(wclk), .Q(ram[2419]) );
  DFF ram_reg_1745__2_ ( .D(n6659), .CP(wclk), .Q(ram[2418]) );
  DFF ram_reg_1745__1_ ( .D(n6658), .CP(wclk), .Q(ram[2417]) );
  DFF ram_reg_1745__0_ ( .D(n6657), .CP(wclk), .Q(ram[2416]) );
  DFF ram_reg_1749__7_ ( .D(n6632), .CP(wclk), .Q(ram[2391]) );
  DFF ram_reg_1749__6_ ( .D(n6631), .CP(wclk), .Q(ram[2390]) );
  DFF ram_reg_1749__5_ ( .D(n6630), .CP(wclk), .Q(ram[2389]) );
  DFF ram_reg_1749__4_ ( .D(n6629), .CP(wclk), .Q(ram[2388]) );
  DFF ram_reg_1749__3_ ( .D(n6628), .CP(wclk), .Q(ram[2387]) );
  DFF ram_reg_1749__2_ ( .D(n6627), .CP(wclk), .Q(ram[2386]) );
  DFF ram_reg_1749__1_ ( .D(n6626), .CP(wclk), .Q(ram[2385]) );
  DFF ram_reg_1749__0_ ( .D(n6625), .CP(wclk), .Q(ram[2384]) );
  DFF ram_reg_1765__7_ ( .D(n6504), .CP(wclk), .Q(ram[2263]) );
  DFF ram_reg_1765__6_ ( .D(n6503), .CP(wclk), .Q(ram[2262]) );
  DFF ram_reg_1765__5_ ( .D(n6502), .CP(wclk), .Q(ram[2261]) );
  DFF ram_reg_1765__4_ ( .D(n6501), .CP(wclk), .Q(ram[2260]) );
  DFF ram_reg_1765__3_ ( .D(n6500), .CP(wclk), .Q(ram[2259]) );
  DFF ram_reg_1765__2_ ( .D(n6499), .CP(wclk), .Q(ram[2258]) );
  DFF ram_reg_1765__1_ ( .D(n6498), .CP(wclk), .Q(ram[2257]) );
  DFF ram_reg_1765__0_ ( .D(n6497), .CP(wclk), .Q(ram[2256]) );
  DFF ram_reg_1781__7_ ( .D(n6376), .CP(wclk), .Q(ram[2135]) );
  DFF ram_reg_1781__6_ ( .D(n6375), .CP(wclk), .Q(ram[2134]) );
  DFF ram_reg_1781__5_ ( .D(n6374), .CP(wclk), .Q(ram[2133]) );
  DFF ram_reg_1781__4_ ( .D(n6373), .CP(wclk), .Q(ram[2132]) );
  DFF ram_reg_1781__3_ ( .D(n6372), .CP(wclk), .Q(ram[2131]) );
  DFF ram_reg_1781__2_ ( .D(n6371), .CP(wclk), .Q(ram[2130]) );
  DFF ram_reg_1781__1_ ( .D(n6370), .CP(wclk), .Q(ram[2129]) );
  DFF ram_reg_1781__0_ ( .D(n6369), .CP(wclk), .Q(ram[2128]) );
  DFF ram_reg_1793__7_ ( .D(n6280), .CP(wclk), .Q(ram[2039]) );
  DFF ram_reg_1793__6_ ( .D(n6279), .CP(wclk), .Q(ram[2038]) );
  DFF ram_reg_1793__5_ ( .D(n6278), .CP(wclk), .Q(ram[2037]) );
  DFF ram_reg_1793__4_ ( .D(n6277), .CP(wclk), .Q(ram[2036]) );
  DFF ram_reg_1793__3_ ( .D(n6276), .CP(wclk), .Q(ram[2035]) );
  DFF ram_reg_1793__2_ ( .D(n6275), .CP(wclk), .Q(ram[2034]) );
  DFF ram_reg_1793__1_ ( .D(n6274), .CP(wclk), .Q(ram[2033]) );
  DFF ram_reg_1793__0_ ( .D(n6273), .CP(wclk), .Q(ram[2032]) );
  DFF ram_reg_1797__7_ ( .D(n6248), .CP(wclk), .Q(ram[2007]) );
  DFF ram_reg_1797__6_ ( .D(n6247), .CP(wclk), .Q(ram[2006]) );
  DFF ram_reg_1797__5_ ( .D(n6246), .CP(wclk), .Q(ram[2005]) );
  DFF ram_reg_1797__4_ ( .D(n6245), .CP(wclk), .Q(ram[2004]) );
  DFF ram_reg_1797__3_ ( .D(n6244), .CP(wclk), .Q(ram[2003]) );
  DFF ram_reg_1797__2_ ( .D(n6243), .CP(wclk), .Q(ram[2002]) );
  DFF ram_reg_1797__1_ ( .D(n6242), .CP(wclk), .Q(ram[2001]) );
  DFF ram_reg_1797__0_ ( .D(n6241), .CP(wclk), .Q(ram[2000]) );
  DFF ram_reg_1809__7_ ( .D(n6152), .CP(wclk), .Q(ram[1911]) );
  DFF ram_reg_1809__6_ ( .D(n6151), .CP(wclk), .Q(ram[1910]) );
  DFF ram_reg_1809__5_ ( .D(n6150), .CP(wclk), .Q(ram[1909]) );
  DFF ram_reg_1809__4_ ( .D(n6149), .CP(wclk), .Q(ram[1908]) );
  DFF ram_reg_1809__3_ ( .D(n6148), .CP(wclk), .Q(ram[1907]) );
  DFF ram_reg_1809__2_ ( .D(n6147), .CP(wclk), .Q(ram[1906]) );
  DFF ram_reg_1809__1_ ( .D(n6146), .CP(wclk), .Q(ram[1905]) );
  DFF ram_reg_1809__0_ ( .D(n6145), .CP(wclk), .Q(ram[1904]) );
  DFF ram_reg_1813__7_ ( .D(n6120), .CP(wclk), .Q(ram[1879]) );
  DFF ram_reg_1813__6_ ( .D(n6119), .CP(wclk), .Q(ram[1878]) );
  DFF ram_reg_1813__5_ ( .D(n6118), .CP(wclk), .Q(ram[1877]) );
  DFF ram_reg_1813__4_ ( .D(n6117), .CP(wclk), .Q(ram[1876]) );
  DFF ram_reg_1813__3_ ( .D(n6116), .CP(wclk), .Q(ram[1875]) );
  DFF ram_reg_1813__2_ ( .D(n6115), .CP(wclk), .Q(ram[1874]) );
  DFF ram_reg_1813__1_ ( .D(n6114), .CP(wclk), .Q(ram[1873]) );
  DFF ram_reg_1813__0_ ( .D(n6113), .CP(wclk), .Q(ram[1872]) );
  DFF ram_reg_1821__7_ ( .D(n6056), .CP(wclk), .Q(ram[1815]) );
  DFF ram_reg_1821__6_ ( .D(n6055), .CP(wclk), .Q(ram[1814]) );
  DFF ram_reg_1821__5_ ( .D(n6054), .CP(wclk), .Q(ram[1813]) );
  DFF ram_reg_1821__4_ ( .D(n6053), .CP(wclk), .Q(ram[1812]) );
  DFF ram_reg_1821__3_ ( .D(n6052), .CP(wclk), .Q(ram[1811]) );
  DFF ram_reg_1821__2_ ( .D(n6051), .CP(wclk), .Q(ram[1810]) );
  DFF ram_reg_1821__1_ ( .D(n6050), .CP(wclk), .Q(ram[1809]) );
  DFF ram_reg_1821__0_ ( .D(n6049), .CP(wclk), .Q(ram[1808]) );
  DFF ram_reg_1829__7_ ( .D(n5992), .CP(wclk), .Q(ram[1751]) );
  DFF ram_reg_1829__6_ ( .D(n5991), .CP(wclk), .Q(ram[1750]) );
  DFF ram_reg_1829__5_ ( .D(n5990), .CP(wclk), .Q(ram[1749]) );
  DFF ram_reg_1829__4_ ( .D(n5989), .CP(wclk), .Q(ram[1748]) );
  DFF ram_reg_1829__3_ ( .D(n5988), .CP(wclk), .Q(ram[1747]) );
  DFF ram_reg_1829__2_ ( .D(n5987), .CP(wclk), .Q(ram[1746]) );
  DFF ram_reg_1829__1_ ( .D(n5986), .CP(wclk), .Q(ram[1745]) );
  DFF ram_reg_1829__0_ ( .D(n5985), .CP(wclk), .Q(ram[1744]) );
  DFF ram_reg_1845__7_ ( .D(n5864), .CP(wclk), .Q(ram[1623]) );
  DFF ram_reg_1845__6_ ( .D(n5863), .CP(wclk), .Q(ram[1622]) );
  DFF ram_reg_1845__5_ ( .D(n5862), .CP(wclk), .Q(ram[1621]) );
  DFF ram_reg_1845__4_ ( .D(n5861), .CP(wclk), .Q(ram[1620]) );
  DFF ram_reg_1845__3_ ( .D(n5860), .CP(wclk), .Q(ram[1619]) );
  DFF ram_reg_1845__2_ ( .D(n5859), .CP(wclk), .Q(ram[1618]) );
  DFF ram_reg_1845__1_ ( .D(n5858), .CP(wclk), .Q(ram[1617]) );
  DFF ram_reg_1845__0_ ( .D(n5857), .CP(wclk), .Q(ram[1616]) );
  DFF ram_reg_1857__7_ ( .D(n5768), .CP(wclk), .Q(ram[1527]) );
  DFF ram_reg_1857__6_ ( .D(n5767), .CP(wclk), .Q(ram[1526]) );
  DFF ram_reg_1857__5_ ( .D(n5766), .CP(wclk), .Q(ram[1525]) );
  DFF ram_reg_1857__4_ ( .D(n5765), .CP(wclk), .Q(ram[1524]) );
  DFF ram_reg_1857__3_ ( .D(n5764), .CP(wclk), .Q(ram[1523]) );
  DFF ram_reg_1857__2_ ( .D(n5763), .CP(wclk), .Q(ram[1522]) );
  DFF ram_reg_1857__1_ ( .D(n5762), .CP(wclk), .Q(ram[1521]) );
  DFF ram_reg_1857__0_ ( .D(n5761), .CP(wclk), .Q(ram[1520]) );
  DFF ram_reg_1861__7_ ( .D(n5736), .CP(wclk), .Q(ram[1495]) );
  DFF ram_reg_1861__6_ ( .D(n5735), .CP(wclk), .Q(ram[1494]) );
  DFF ram_reg_1861__5_ ( .D(n5734), .CP(wclk), .Q(ram[1493]) );
  DFF ram_reg_1861__4_ ( .D(n5733), .CP(wclk), .Q(ram[1492]) );
  DFF ram_reg_1861__3_ ( .D(n5732), .CP(wclk), .Q(ram[1491]) );
  DFF ram_reg_1861__2_ ( .D(n5731), .CP(wclk), .Q(ram[1490]) );
  DFF ram_reg_1861__1_ ( .D(n5730), .CP(wclk), .Q(ram[1489]) );
  DFF ram_reg_1861__0_ ( .D(n5729), .CP(wclk), .Q(ram[1488]) );
  DFF ram_reg_1865__7_ ( .D(n5704), .CP(wclk), .Q(ram[1463]) );
  DFF ram_reg_1865__6_ ( .D(n5703), .CP(wclk), .Q(ram[1462]) );
  DFF ram_reg_1865__5_ ( .D(n5702), .CP(wclk), .Q(ram[1461]) );
  DFF ram_reg_1865__4_ ( .D(n5701), .CP(wclk), .Q(ram[1460]) );
  DFF ram_reg_1865__3_ ( .D(n5700), .CP(wclk), .Q(ram[1459]) );
  DFF ram_reg_1865__2_ ( .D(n5699), .CP(wclk), .Q(ram[1458]) );
  DFF ram_reg_1865__1_ ( .D(n5698), .CP(wclk), .Q(ram[1457]) );
  DFF ram_reg_1865__0_ ( .D(n5697), .CP(wclk), .Q(ram[1456]) );
  DFF ram_reg_1869__7_ ( .D(n5672), .CP(wclk), .Q(ram[1431]) );
  DFF ram_reg_1869__6_ ( .D(n5671), .CP(wclk), .Q(ram[1430]) );
  DFF ram_reg_1869__5_ ( .D(n5670), .CP(wclk), .Q(ram[1429]) );
  DFF ram_reg_1869__4_ ( .D(n5669), .CP(wclk), .Q(ram[1428]) );
  DFF ram_reg_1869__3_ ( .D(n5668), .CP(wclk), .Q(ram[1427]) );
  DFF ram_reg_1869__2_ ( .D(n5667), .CP(wclk), .Q(ram[1426]) );
  DFF ram_reg_1869__1_ ( .D(n5666), .CP(wclk), .Q(ram[1425]) );
  DFF ram_reg_1869__0_ ( .D(n5665), .CP(wclk), .Q(ram[1424]) );
  DFF ram_reg_1873__7_ ( .D(n5640), .CP(wclk), .Q(ram[1399]) );
  DFF ram_reg_1873__6_ ( .D(n5639), .CP(wclk), .Q(ram[1398]) );
  DFF ram_reg_1873__5_ ( .D(n5638), .CP(wclk), .Q(ram[1397]) );
  DFF ram_reg_1873__4_ ( .D(n5637), .CP(wclk), .Q(ram[1396]) );
  DFF ram_reg_1873__3_ ( .D(n5636), .CP(wclk), .Q(ram[1395]) );
  DFF ram_reg_1873__2_ ( .D(n5635), .CP(wclk), .Q(ram[1394]) );
  DFF ram_reg_1873__1_ ( .D(n5634), .CP(wclk), .Q(ram[1393]) );
  DFF ram_reg_1873__0_ ( .D(n5633), .CP(wclk), .Q(ram[1392]) );
  DFF ram_reg_1877__7_ ( .D(n5608), .CP(wclk), .Q(ram[1367]) );
  DFF ram_reg_1877__6_ ( .D(n5607), .CP(wclk), .Q(ram[1366]) );
  DFF ram_reg_1877__5_ ( .D(n5606), .CP(wclk), .Q(ram[1365]) );
  DFF ram_reg_1877__4_ ( .D(n5605), .CP(wclk), .Q(ram[1364]) );
  DFF ram_reg_1877__3_ ( .D(n5604), .CP(wclk), .Q(ram[1363]) );
  DFF ram_reg_1877__2_ ( .D(n5603), .CP(wclk), .Q(ram[1362]) );
  DFF ram_reg_1877__1_ ( .D(n5602), .CP(wclk), .Q(ram[1361]) );
  DFF ram_reg_1877__0_ ( .D(n5601), .CP(wclk), .Q(ram[1360]) );
  DFF ram_reg_1881__7_ ( .D(n5576), .CP(wclk), .Q(ram[1335]) );
  DFF ram_reg_1881__6_ ( .D(n5575), .CP(wclk), .Q(ram[1334]) );
  DFF ram_reg_1881__5_ ( .D(n5574), .CP(wclk), .Q(ram[1333]) );
  DFF ram_reg_1881__4_ ( .D(n5573), .CP(wclk), .Q(ram[1332]) );
  DFF ram_reg_1881__3_ ( .D(n5572), .CP(wclk), .Q(ram[1331]) );
  DFF ram_reg_1881__2_ ( .D(n5571), .CP(wclk), .Q(ram[1330]) );
  DFF ram_reg_1881__1_ ( .D(n5570), .CP(wclk), .Q(ram[1329]) );
  DFF ram_reg_1881__0_ ( .D(n5569), .CP(wclk), .Q(ram[1328]) );
  DFF ram_reg_1885__7_ ( .D(n5544), .CP(wclk), .Q(ram[1303]) );
  DFF ram_reg_1885__6_ ( .D(n5543), .CP(wclk), .Q(ram[1302]) );
  DFF ram_reg_1885__5_ ( .D(n5542), .CP(wclk), .Q(ram[1301]) );
  DFF ram_reg_1885__4_ ( .D(n5541), .CP(wclk), .Q(ram[1300]) );
  DFF ram_reg_1885__3_ ( .D(n5540), .CP(wclk), .Q(ram[1299]) );
  DFF ram_reg_1885__2_ ( .D(n5539), .CP(wclk), .Q(ram[1298]) );
  DFF ram_reg_1885__1_ ( .D(n5538), .CP(wclk), .Q(ram[1297]) );
  DFF ram_reg_1885__0_ ( .D(n5537), .CP(wclk), .Q(ram[1296]) );
  DFF ram_reg_1889__7_ ( .D(n5512), .CP(wclk), .Q(ram[1271]) );
  DFF ram_reg_1889__6_ ( .D(n5511), .CP(wclk), .Q(ram[1270]) );
  DFF ram_reg_1889__5_ ( .D(n5510), .CP(wclk), .Q(ram[1269]) );
  DFF ram_reg_1889__4_ ( .D(n5509), .CP(wclk), .Q(ram[1268]) );
  DFF ram_reg_1889__3_ ( .D(n5508), .CP(wclk), .Q(ram[1267]) );
  DFF ram_reg_1889__2_ ( .D(n5507), .CP(wclk), .Q(ram[1266]) );
  DFF ram_reg_1889__1_ ( .D(n5506), .CP(wclk), .Q(ram[1265]) );
  DFF ram_reg_1889__0_ ( .D(n5505), .CP(wclk), .Q(ram[1264]) );
  DFF ram_reg_1893__7_ ( .D(n5480), .CP(wclk), .Q(ram[1239]) );
  DFF ram_reg_1893__6_ ( .D(n5479), .CP(wclk), .Q(ram[1238]) );
  DFF ram_reg_1893__5_ ( .D(n5478), .CP(wclk), .Q(ram[1237]) );
  DFF ram_reg_1893__4_ ( .D(n5477), .CP(wclk), .Q(ram[1236]) );
  DFF ram_reg_1893__3_ ( .D(n5476), .CP(wclk), .Q(ram[1235]) );
  DFF ram_reg_1893__2_ ( .D(n5475), .CP(wclk), .Q(ram[1234]) );
  DFF ram_reg_1893__1_ ( .D(n5474), .CP(wclk), .Q(ram[1233]) );
  DFF ram_reg_1893__0_ ( .D(n5473), .CP(wclk), .Q(ram[1232]) );
  DFF ram_reg_1901__7_ ( .D(n5416), .CP(wclk), .Q(ram[1175]) );
  DFF ram_reg_1901__6_ ( .D(n5415), .CP(wclk), .Q(ram[1174]) );
  DFF ram_reg_1901__5_ ( .D(n5414), .CP(wclk), .Q(ram[1173]) );
  DFF ram_reg_1901__4_ ( .D(n5413), .CP(wclk), .Q(ram[1172]) );
  DFF ram_reg_1901__3_ ( .D(n5412), .CP(wclk), .Q(ram[1171]) );
  DFF ram_reg_1901__2_ ( .D(n5411), .CP(wclk), .Q(ram[1170]) );
  DFF ram_reg_1901__1_ ( .D(n5410), .CP(wclk), .Q(ram[1169]) );
  DFF ram_reg_1901__0_ ( .D(n5409), .CP(wclk), .Q(ram[1168]) );
  DFF ram_reg_1905__7_ ( .D(n5384), .CP(wclk), .Q(ram[1143]) );
  DFF ram_reg_1905__6_ ( .D(n5383), .CP(wclk), .Q(ram[1142]) );
  DFF ram_reg_1905__5_ ( .D(n5382), .CP(wclk), .Q(ram[1141]) );
  DFF ram_reg_1905__4_ ( .D(n5381), .CP(wclk), .Q(ram[1140]) );
  DFF ram_reg_1905__3_ ( .D(n5380), .CP(wclk), .Q(ram[1139]) );
  DFF ram_reg_1905__2_ ( .D(n5379), .CP(wclk), .Q(ram[1138]) );
  DFF ram_reg_1905__1_ ( .D(n5378), .CP(wclk), .Q(ram[1137]) );
  DFF ram_reg_1905__0_ ( .D(n5377), .CP(wclk), .Q(ram[1136]) );
  DFF ram_reg_1909__7_ ( .D(n5352), .CP(wclk), .Q(ram[1111]) );
  DFF ram_reg_1909__6_ ( .D(n5351), .CP(wclk), .Q(ram[1110]) );
  DFF ram_reg_1909__5_ ( .D(n5350), .CP(wclk), .Q(ram[1109]) );
  DFF ram_reg_1909__4_ ( .D(n5349), .CP(wclk), .Q(ram[1108]) );
  DFF ram_reg_1909__3_ ( .D(n5348), .CP(wclk), .Q(ram[1107]) );
  DFF ram_reg_1909__2_ ( .D(n5347), .CP(wclk), .Q(ram[1106]) );
  DFF ram_reg_1909__1_ ( .D(n5346), .CP(wclk), .Q(ram[1105]) );
  DFF ram_reg_1909__0_ ( .D(n5345), .CP(wclk), .Q(ram[1104]) );
  DFF ram_reg_1925__7_ ( .D(n5224), .CP(wclk), .Q(ram[983]) );
  DFF ram_reg_1925__6_ ( .D(n5223), .CP(wclk), .Q(ram[982]) );
  DFF ram_reg_1925__5_ ( .D(n5222), .CP(wclk), .Q(ram[981]) );
  DFF ram_reg_1925__4_ ( .D(n5221), .CP(wclk), .Q(ram[980]) );
  DFF ram_reg_1925__3_ ( .D(n5220), .CP(wclk), .Q(ram[979]) );
  DFF ram_reg_1925__2_ ( .D(n5219), .CP(wclk), .Q(ram[978]) );
  DFF ram_reg_1925__1_ ( .D(n5218), .CP(wclk), .Q(ram[977]) );
  DFF ram_reg_1925__0_ ( .D(n5217), .CP(wclk), .Q(ram[976]) );
  DFF ram_reg_1941__7_ ( .D(n5096), .CP(wclk), .Q(ram[855]) );
  DFF ram_reg_1941__6_ ( .D(n5095), .CP(wclk), .Q(ram[854]) );
  DFF ram_reg_1941__5_ ( .D(n5094), .CP(wclk), .Q(ram[853]) );
  DFF ram_reg_1941__4_ ( .D(n5093), .CP(wclk), .Q(ram[852]) );
  DFF ram_reg_1941__3_ ( .D(n5092), .CP(wclk), .Q(ram[851]) );
  DFF ram_reg_1941__2_ ( .D(n5091), .CP(wclk), .Q(ram[850]) );
  DFF ram_reg_1941__1_ ( .D(n5090), .CP(wclk), .Q(ram[849]) );
  DFF ram_reg_1941__0_ ( .D(n5089), .CP(wclk), .Q(ram[848]) );
  DFF ram_reg_1989__7_ ( .D(n4712), .CP(wclk), .Q(ram[471]) );
  DFF ram_reg_1989__6_ ( .D(n4711), .CP(wclk), .Q(ram[470]) );
  DFF ram_reg_1989__5_ ( .D(n4710), .CP(wclk), .Q(ram[469]) );
  DFF ram_reg_1989__4_ ( .D(n4709), .CP(wclk), .Q(ram[468]) );
  DFF ram_reg_1989__3_ ( .D(n4708), .CP(wclk), .Q(ram[467]) );
  DFF ram_reg_1989__2_ ( .D(n4707), .CP(wclk), .Q(ram[466]) );
  DFF ram_reg_1989__1_ ( .D(n4706), .CP(wclk), .Q(ram[465]) );
  DFF ram_reg_1989__0_ ( .D(n4705), .CP(wclk), .Q(ram[464]) );
  DFF ram_reg_2001__7_ ( .D(n4616), .CP(wclk), .Q(ram[375]) );
  DFF ram_reg_2001__6_ ( .D(n4615), .CP(wclk), .Q(ram[374]) );
  DFF ram_reg_2001__5_ ( .D(n4614), .CP(wclk), .Q(ram[373]) );
  DFF ram_reg_2001__4_ ( .D(n4613), .CP(wclk), .Q(ram[372]) );
  DFF ram_reg_2001__3_ ( .D(n4612), .CP(wclk), .Q(ram[371]) );
  DFF ram_reg_2001__2_ ( .D(n4611), .CP(wclk), .Q(ram[370]) );
  DFF ram_reg_2001__1_ ( .D(n4610), .CP(wclk), .Q(ram[369]) );
  DFF ram_reg_2001__0_ ( .D(n4609), .CP(wclk), .Q(ram[368]) );
  DFF ram_reg_2005__7_ ( .D(n4584), .CP(wclk), .Q(ram[343]) );
  DFF ram_reg_2005__6_ ( .D(n4583), .CP(wclk), .Q(ram[342]) );
  DFF ram_reg_2005__5_ ( .D(n4582), .CP(wclk), .Q(ram[341]) );
  DFF ram_reg_2005__4_ ( .D(n4581), .CP(wclk), .Q(ram[340]) );
  DFF ram_reg_2005__3_ ( .D(n4580), .CP(wclk), .Q(ram[339]) );
  DFF ram_reg_2005__2_ ( .D(n4579), .CP(wclk), .Q(ram[338]) );
  DFF ram_reg_2005__1_ ( .D(n4578), .CP(wclk), .Q(ram[337]) );
  DFF ram_reg_2005__0_ ( .D(n4577), .CP(wclk), .Q(ram[336]) );
  DFF ram_reg_2021__7_ ( .D(n4456), .CP(wclk), .Q(ram[215]) );
  DFF ram_reg_2021__6_ ( .D(n4455), .CP(wclk), .Q(ram[214]) );
  DFF ram_reg_2021__5_ ( .D(n4454), .CP(wclk), .Q(ram[213]) );
  DFF ram_reg_2021__4_ ( .D(n4453), .CP(wclk), .Q(ram[212]) );
  DFF ram_reg_2021__3_ ( .D(n4452), .CP(wclk), .Q(ram[211]) );
  DFF ram_reg_2021__2_ ( .D(n4451), .CP(wclk), .Q(ram[210]) );
  DFF ram_reg_2021__1_ ( .D(n4450), .CP(wclk), .Q(ram[209]) );
  DFF ram_reg_2021__0_ ( .D(n4449), .CP(wclk), .Q(ram[208]) );
  DFF ram_reg_3__7_ ( .D(n20600), .CP(wclk), .Q(ram[16359]) );
  DFF ram_reg_3__6_ ( .D(n20599), .CP(wclk), .Q(ram[16358]) );
  DFF ram_reg_3__5_ ( .D(n20598), .CP(wclk), .Q(ram[16357]) );
  DFF ram_reg_3__4_ ( .D(n20597), .CP(wclk), .Q(ram[16356]) );
  DFF ram_reg_3__3_ ( .D(n20596), .CP(wclk), .Q(ram[16355]) );
  DFF ram_reg_3__2_ ( .D(n20595), .CP(wclk), .Q(ram[16354]) );
  DFF ram_reg_3__1_ ( .D(n20594), .CP(wclk), .Q(ram[16353]) );
  DFF ram_reg_3__0_ ( .D(n20593), .CP(wclk), .Q(ram[16352]) );
  DFF ram_reg_7__7_ ( .D(n20568), .CP(wclk), .Q(ram[16327]) );
  DFF ram_reg_7__6_ ( .D(n20567), .CP(wclk), .Q(ram[16326]) );
  DFF ram_reg_7__5_ ( .D(n20566), .CP(wclk), .Q(ram[16325]) );
  DFF ram_reg_7__4_ ( .D(n20565), .CP(wclk), .Q(ram[16324]) );
  DFF ram_reg_7__3_ ( .D(n20564), .CP(wclk), .Q(ram[16323]) );
  DFF ram_reg_7__2_ ( .D(n20563), .CP(wclk), .Q(ram[16322]) );
  DFF ram_reg_7__1_ ( .D(n20562), .CP(wclk), .Q(ram[16321]) );
  DFF ram_reg_7__0_ ( .D(n20561), .CP(wclk), .Q(ram[16320]) );
  DFF ram_reg_15__7_ ( .D(n20504), .CP(wclk), .Q(ram[16263]) );
  DFF ram_reg_15__6_ ( .D(n20503), .CP(wclk), .Q(ram[16262]) );
  DFF ram_reg_15__5_ ( .D(n20502), .CP(wclk), .Q(ram[16261]) );
  DFF ram_reg_15__4_ ( .D(n20501), .CP(wclk), .Q(ram[16260]) );
  DFF ram_reg_15__3_ ( .D(n20500), .CP(wclk), .Q(ram[16259]) );
  DFF ram_reg_15__2_ ( .D(n20499), .CP(wclk), .Q(ram[16258]) );
  DFF ram_reg_15__1_ ( .D(n20498), .CP(wclk), .Q(ram[16257]) );
  DFF ram_reg_15__0_ ( .D(n20497), .CP(wclk), .Q(ram[16256]) );
  DFF ram_reg_19__7_ ( .D(n20472), .CP(wclk), .Q(ram[16231]) );
  DFF ram_reg_19__6_ ( .D(n20471), .CP(wclk), .Q(ram[16230]) );
  DFF ram_reg_19__5_ ( .D(n20470), .CP(wclk), .Q(ram[16229]) );
  DFF ram_reg_19__4_ ( .D(n20469), .CP(wclk), .Q(ram[16228]) );
  DFF ram_reg_19__3_ ( .D(n20468), .CP(wclk), .Q(ram[16227]) );
  DFF ram_reg_19__2_ ( .D(n20467), .CP(wclk), .Q(ram[16226]) );
  DFF ram_reg_19__1_ ( .D(n20466), .CP(wclk), .Q(ram[16225]) );
  DFF ram_reg_19__0_ ( .D(n20465), .CP(wclk), .Q(ram[16224]) );
  DFF ram_reg_23__7_ ( .D(n20440), .CP(wclk), .Q(ram[16199]) );
  DFF ram_reg_23__6_ ( .D(n20439), .CP(wclk), .Q(ram[16198]) );
  DFF ram_reg_23__5_ ( .D(n20438), .CP(wclk), .Q(ram[16197]) );
  DFF ram_reg_23__4_ ( .D(n20437), .CP(wclk), .Q(ram[16196]) );
  DFF ram_reg_23__3_ ( .D(n20436), .CP(wclk), .Q(ram[16195]) );
  DFF ram_reg_23__2_ ( .D(n20435), .CP(wclk), .Q(ram[16194]) );
  DFF ram_reg_23__1_ ( .D(n20434), .CP(wclk), .Q(ram[16193]) );
  DFF ram_reg_23__0_ ( .D(n20433), .CP(wclk), .Q(ram[16192]) );
  DFF ram_reg_27__7_ ( .D(n20408), .CP(wclk), .Q(ram[16167]) );
  DFF ram_reg_27__6_ ( .D(n20407), .CP(wclk), .Q(ram[16166]) );
  DFF ram_reg_27__5_ ( .D(n20406), .CP(wclk), .Q(ram[16165]) );
  DFF ram_reg_27__4_ ( .D(n20405), .CP(wclk), .Q(ram[16164]) );
  DFF ram_reg_27__3_ ( .D(n20404), .CP(wclk), .Q(ram[16163]) );
  DFF ram_reg_27__2_ ( .D(n20403), .CP(wclk), .Q(ram[16162]) );
  DFF ram_reg_27__1_ ( .D(n20402), .CP(wclk), .Q(ram[16161]) );
  DFF ram_reg_27__0_ ( .D(n20401), .CP(wclk), .Q(ram[16160]) );
  DFF ram_reg_31__7_ ( .D(n20376), .CP(wclk), .Q(ram[16135]) );
  DFF ram_reg_31__6_ ( .D(n20375), .CP(wclk), .Q(ram[16134]) );
  DFF ram_reg_31__5_ ( .D(n20374), .CP(wclk), .Q(ram[16133]) );
  DFF ram_reg_31__4_ ( .D(n20373), .CP(wclk), .Q(ram[16132]) );
  DFF ram_reg_31__3_ ( .D(n20372), .CP(wclk), .Q(ram[16131]) );
  DFF ram_reg_31__2_ ( .D(n20371), .CP(wclk), .Q(ram[16130]) );
  DFF ram_reg_31__1_ ( .D(n20370), .CP(wclk), .Q(ram[16129]) );
  DFF ram_reg_31__0_ ( .D(n20369), .CP(wclk), .Q(ram[16128]) );
  DFF ram_reg_35__7_ ( .D(n20344), .CP(wclk), .Q(ram[16103]) );
  DFF ram_reg_35__6_ ( .D(n20343), .CP(wclk), .Q(ram[16102]) );
  DFF ram_reg_35__5_ ( .D(n20342), .CP(wclk), .Q(ram[16101]) );
  DFF ram_reg_35__4_ ( .D(n20341), .CP(wclk), .Q(ram[16100]) );
  DFF ram_reg_35__3_ ( .D(n20340), .CP(wclk), .Q(ram[16099]) );
  DFF ram_reg_35__2_ ( .D(n20339), .CP(wclk), .Q(ram[16098]) );
  DFF ram_reg_35__1_ ( .D(n20338), .CP(wclk), .Q(ram[16097]) );
  DFF ram_reg_35__0_ ( .D(n20337), .CP(wclk), .Q(ram[16096]) );
  DFF ram_reg_39__7_ ( .D(n20312), .CP(wclk), .Q(ram[16071]) );
  DFF ram_reg_39__6_ ( .D(n20311), .CP(wclk), .Q(ram[16070]) );
  DFF ram_reg_39__5_ ( .D(n20310), .CP(wclk), .Q(ram[16069]) );
  DFF ram_reg_39__4_ ( .D(n20309), .CP(wclk), .Q(ram[16068]) );
  DFF ram_reg_39__3_ ( .D(n20308), .CP(wclk), .Q(ram[16067]) );
  DFF ram_reg_39__2_ ( .D(n20307), .CP(wclk), .Q(ram[16066]) );
  DFF ram_reg_39__1_ ( .D(n20306), .CP(wclk), .Q(ram[16065]) );
  DFF ram_reg_39__0_ ( .D(n20305), .CP(wclk), .Q(ram[16064]) );
  DFF ram_reg_51__7_ ( .D(n20216), .CP(wclk), .Q(ram[15975]) );
  DFF ram_reg_51__6_ ( .D(n20215), .CP(wclk), .Q(ram[15974]) );
  DFF ram_reg_51__5_ ( .D(n20214), .CP(wclk), .Q(ram[15973]) );
  DFF ram_reg_51__4_ ( .D(n20213), .CP(wclk), .Q(ram[15972]) );
  DFF ram_reg_51__3_ ( .D(n20212), .CP(wclk), .Q(ram[15971]) );
  DFF ram_reg_51__2_ ( .D(n20211), .CP(wclk), .Q(ram[15970]) );
  DFF ram_reg_51__1_ ( .D(n20210), .CP(wclk), .Q(ram[15969]) );
  DFF ram_reg_51__0_ ( .D(n20209), .CP(wclk), .Q(ram[15968]) );
  DFF ram_reg_55__7_ ( .D(n20184), .CP(wclk), .Q(ram[15943]) );
  DFF ram_reg_55__6_ ( .D(n20183), .CP(wclk), .Q(ram[15942]) );
  DFF ram_reg_55__5_ ( .D(n20182), .CP(wclk), .Q(ram[15941]) );
  DFF ram_reg_55__4_ ( .D(n20181), .CP(wclk), .Q(ram[15940]) );
  DFF ram_reg_55__3_ ( .D(n20180), .CP(wclk), .Q(ram[15939]) );
  DFF ram_reg_55__2_ ( .D(n20179), .CP(wclk), .Q(ram[15938]) );
  DFF ram_reg_55__1_ ( .D(n20178), .CP(wclk), .Q(ram[15937]) );
  DFF ram_reg_55__0_ ( .D(n20177), .CP(wclk), .Q(ram[15936]) );
  DFF ram_reg_67__7_ ( .D(n20088), .CP(wclk), .Q(ram[15847]) );
  DFF ram_reg_67__6_ ( .D(n20087), .CP(wclk), .Q(ram[15846]) );
  DFF ram_reg_67__5_ ( .D(n20086), .CP(wclk), .Q(ram[15845]) );
  DFF ram_reg_67__4_ ( .D(n20085), .CP(wclk), .Q(ram[15844]) );
  DFF ram_reg_67__3_ ( .D(n20084), .CP(wclk), .Q(ram[15843]) );
  DFF ram_reg_67__2_ ( .D(n20083), .CP(wclk), .Q(ram[15842]) );
  DFF ram_reg_67__1_ ( .D(n20082), .CP(wclk), .Q(ram[15841]) );
  DFF ram_reg_67__0_ ( .D(n20081), .CP(wclk), .Q(ram[15840]) );
  DFF ram_reg_71__7_ ( .D(n20056), .CP(wclk), .Q(ram[15815]) );
  DFF ram_reg_71__6_ ( .D(n20055), .CP(wclk), .Q(ram[15814]) );
  DFF ram_reg_71__5_ ( .D(n20054), .CP(wclk), .Q(ram[15813]) );
  DFF ram_reg_71__4_ ( .D(n20053), .CP(wclk), .Q(ram[15812]) );
  DFF ram_reg_71__3_ ( .D(n20052), .CP(wclk), .Q(ram[15811]) );
  DFF ram_reg_71__2_ ( .D(n20051), .CP(wclk), .Q(ram[15810]) );
  DFF ram_reg_71__1_ ( .D(n20050), .CP(wclk), .Q(ram[15809]) );
  DFF ram_reg_71__0_ ( .D(n20049), .CP(wclk), .Q(ram[15808]) );
  DFF ram_reg_75__7_ ( .D(n20024), .CP(wclk), .Q(ram[15783]) );
  DFF ram_reg_75__6_ ( .D(n20023), .CP(wclk), .Q(ram[15782]) );
  DFF ram_reg_75__5_ ( .D(n20022), .CP(wclk), .Q(ram[15781]) );
  DFF ram_reg_75__4_ ( .D(n20021), .CP(wclk), .Q(ram[15780]) );
  DFF ram_reg_75__3_ ( .D(n20020), .CP(wclk), .Q(ram[15779]) );
  DFF ram_reg_75__2_ ( .D(n20019), .CP(wclk), .Q(ram[15778]) );
  DFF ram_reg_75__1_ ( .D(n20018), .CP(wclk), .Q(ram[15777]) );
  DFF ram_reg_75__0_ ( .D(n20017), .CP(wclk), .Q(ram[15776]) );
  DFF ram_reg_79__7_ ( .D(n19992), .CP(wclk), .Q(ram[15751]) );
  DFF ram_reg_79__6_ ( .D(n19991), .CP(wclk), .Q(ram[15750]) );
  DFF ram_reg_79__5_ ( .D(n19990), .CP(wclk), .Q(ram[15749]) );
  DFF ram_reg_79__4_ ( .D(n19989), .CP(wclk), .Q(ram[15748]) );
  DFF ram_reg_79__3_ ( .D(n19988), .CP(wclk), .Q(ram[15747]) );
  DFF ram_reg_79__2_ ( .D(n19987), .CP(wclk), .Q(ram[15746]) );
  DFF ram_reg_79__1_ ( .D(n19986), .CP(wclk), .Q(ram[15745]) );
  DFF ram_reg_79__0_ ( .D(n19985), .CP(wclk), .Q(ram[15744]) );
  DFF ram_reg_83__7_ ( .D(n19960), .CP(wclk), .Q(ram[15719]) );
  DFF ram_reg_83__6_ ( .D(n19959), .CP(wclk), .Q(ram[15718]) );
  DFF ram_reg_83__5_ ( .D(n19958), .CP(wclk), .Q(ram[15717]) );
  DFF ram_reg_83__4_ ( .D(n19957), .CP(wclk), .Q(ram[15716]) );
  DFF ram_reg_83__3_ ( .D(n19956), .CP(wclk), .Q(ram[15715]) );
  DFF ram_reg_83__2_ ( .D(n19955), .CP(wclk), .Q(ram[15714]) );
  DFF ram_reg_83__1_ ( .D(n19954), .CP(wclk), .Q(ram[15713]) );
  DFF ram_reg_83__0_ ( .D(n19953), .CP(wclk), .Q(ram[15712]) );
  DFF ram_reg_87__7_ ( .D(n19928), .CP(wclk), .Q(ram[15687]) );
  DFF ram_reg_87__6_ ( .D(n19927), .CP(wclk), .Q(ram[15686]) );
  DFF ram_reg_87__5_ ( .D(n19926), .CP(wclk), .Q(ram[15685]) );
  DFF ram_reg_87__4_ ( .D(n19925), .CP(wclk), .Q(ram[15684]) );
  DFF ram_reg_87__3_ ( .D(n19924), .CP(wclk), .Q(ram[15683]) );
  DFF ram_reg_87__2_ ( .D(n19923), .CP(wclk), .Q(ram[15682]) );
  DFF ram_reg_87__1_ ( .D(n19922), .CP(wclk), .Q(ram[15681]) );
  DFF ram_reg_87__0_ ( .D(n19921), .CP(wclk), .Q(ram[15680]) );
  DFF ram_reg_91__7_ ( .D(n19896), .CP(wclk), .Q(ram[15655]) );
  DFF ram_reg_91__6_ ( .D(n19895), .CP(wclk), .Q(ram[15654]) );
  DFF ram_reg_91__5_ ( .D(n19894), .CP(wclk), .Q(ram[15653]) );
  DFF ram_reg_91__4_ ( .D(n19893), .CP(wclk), .Q(ram[15652]) );
  DFF ram_reg_91__3_ ( .D(n19892), .CP(wclk), .Q(ram[15651]) );
  DFF ram_reg_91__2_ ( .D(n19891), .CP(wclk), .Q(ram[15650]) );
  DFF ram_reg_91__1_ ( .D(n19890), .CP(wclk), .Q(ram[15649]) );
  DFF ram_reg_91__0_ ( .D(n19889), .CP(wclk), .Q(ram[15648]) );
  DFF ram_reg_95__7_ ( .D(n19864), .CP(wclk), .Q(ram[15623]) );
  DFF ram_reg_95__6_ ( .D(n19863), .CP(wclk), .Q(ram[15622]) );
  DFF ram_reg_95__5_ ( .D(n19862), .CP(wclk), .Q(ram[15621]) );
  DFF ram_reg_95__4_ ( .D(n19861), .CP(wclk), .Q(ram[15620]) );
  DFF ram_reg_95__3_ ( .D(n19860), .CP(wclk), .Q(ram[15619]) );
  DFF ram_reg_95__2_ ( .D(n19859), .CP(wclk), .Q(ram[15618]) );
  DFF ram_reg_95__1_ ( .D(n19858), .CP(wclk), .Q(ram[15617]) );
  DFF ram_reg_95__0_ ( .D(n19857), .CP(wclk), .Q(ram[15616]) );
  DFF ram_reg_99__7_ ( .D(n19832), .CP(wclk), .Q(ram[15591]) );
  DFF ram_reg_99__6_ ( .D(n19831), .CP(wclk), .Q(ram[15590]) );
  DFF ram_reg_99__5_ ( .D(n19830), .CP(wclk), .Q(ram[15589]) );
  DFF ram_reg_99__4_ ( .D(n19829), .CP(wclk), .Q(ram[15588]) );
  DFF ram_reg_99__3_ ( .D(n19828), .CP(wclk), .Q(ram[15587]) );
  DFF ram_reg_99__2_ ( .D(n19827), .CP(wclk), .Q(ram[15586]) );
  DFF ram_reg_99__1_ ( .D(n19826), .CP(wclk), .Q(ram[15585]) );
  DFF ram_reg_99__0_ ( .D(n19825), .CP(wclk), .Q(ram[15584]) );
  DFF ram_reg_103__7_ ( .D(n19800), .CP(wclk), .Q(ram[15559]) );
  DFF ram_reg_103__6_ ( .D(n19799), .CP(wclk), .Q(ram[15558]) );
  DFF ram_reg_103__5_ ( .D(n19798), .CP(wclk), .Q(ram[15557]) );
  DFF ram_reg_103__4_ ( .D(n19797), .CP(wclk), .Q(ram[15556]) );
  DFF ram_reg_103__3_ ( .D(n19796), .CP(wclk), .Q(ram[15555]) );
  DFF ram_reg_103__2_ ( .D(n19795), .CP(wclk), .Q(ram[15554]) );
  DFF ram_reg_103__1_ ( .D(n19794), .CP(wclk), .Q(ram[15553]) );
  DFF ram_reg_103__0_ ( .D(n19793), .CP(wclk), .Q(ram[15552]) );
  DFF ram_reg_107__7_ ( .D(n19768), .CP(wclk), .Q(ram[15527]) );
  DFF ram_reg_107__6_ ( .D(n19767), .CP(wclk), .Q(ram[15526]) );
  DFF ram_reg_107__5_ ( .D(n19766), .CP(wclk), .Q(ram[15525]) );
  DFF ram_reg_107__4_ ( .D(n19765), .CP(wclk), .Q(ram[15524]) );
  DFF ram_reg_107__3_ ( .D(n19764), .CP(wclk), .Q(ram[15523]) );
  DFF ram_reg_107__2_ ( .D(n19763), .CP(wclk), .Q(ram[15522]) );
  DFF ram_reg_107__1_ ( .D(n19762), .CP(wclk), .Q(ram[15521]) );
  DFF ram_reg_107__0_ ( .D(n19761), .CP(wclk), .Q(ram[15520]) );
  DFF ram_reg_111__7_ ( .D(n19736), .CP(wclk), .Q(ram[15495]) );
  DFF ram_reg_111__6_ ( .D(n19735), .CP(wclk), .Q(ram[15494]) );
  DFF ram_reg_111__5_ ( .D(n19734), .CP(wclk), .Q(ram[15493]) );
  DFF ram_reg_111__4_ ( .D(n19733), .CP(wclk), .Q(ram[15492]) );
  DFF ram_reg_111__3_ ( .D(n19732), .CP(wclk), .Q(ram[15491]) );
  DFF ram_reg_111__2_ ( .D(n19731), .CP(wclk), .Q(ram[15490]) );
  DFF ram_reg_111__1_ ( .D(n19730), .CP(wclk), .Q(ram[15489]) );
  DFF ram_reg_111__0_ ( .D(n19729), .CP(wclk), .Q(ram[15488]) );
  DFF ram_reg_115__7_ ( .D(n19704), .CP(wclk), .Q(ram[15463]) );
  DFF ram_reg_115__6_ ( .D(n19703), .CP(wclk), .Q(ram[15462]) );
  DFF ram_reg_115__5_ ( .D(n19702), .CP(wclk), .Q(ram[15461]) );
  DFF ram_reg_115__4_ ( .D(n19701), .CP(wclk), .Q(ram[15460]) );
  DFF ram_reg_115__3_ ( .D(n19700), .CP(wclk), .Q(ram[15459]) );
  DFF ram_reg_115__2_ ( .D(n19699), .CP(wclk), .Q(ram[15458]) );
  DFF ram_reg_115__1_ ( .D(n19698), .CP(wclk), .Q(ram[15457]) );
  DFF ram_reg_115__0_ ( .D(n19697), .CP(wclk), .Q(ram[15456]) );
  DFF ram_reg_119__7_ ( .D(n19672), .CP(wclk), .Q(ram[15431]) );
  DFF ram_reg_119__6_ ( .D(n19671), .CP(wclk), .Q(ram[15430]) );
  DFF ram_reg_119__5_ ( .D(n19670), .CP(wclk), .Q(ram[15429]) );
  DFF ram_reg_119__4_ ( .D(n19669), .CP(wclk), .Q(ram[15428]) );
  DFF ram_reg_119__3_ ( .D(n19668), .CP(wclk), .Q(ram[15427]) );
  DFF ram_reg_119__2_ ( .D(n19667), .CP(wclk), .Q(ram[15426]) );
  DFF ram_reg_119__1_ ( .D(n19666), .CP(wclk), .Q(ram[15425]) );
  DFF ram_reg_119__0_ ( .D(n19665), .CP(wclk), .Q(ram[15424]) );
  DFF ram_reg_127__7_ ( .D(n19608), .CP(wclk), .Q(ram[15367]) );
  DFF ram_reg_127__6_ ( .D(n19607), .CP(wclk), .Q(ram[15366]) );
  DFF ram_reg_127__5_ ( .D(n19606), .CP(wclk), .Q(ram[15365]) );
  DFF ram_reg_127__4_ ( .D(n19605), .CP(wclk), .Q(ram[15364]) );
  DFF ram_reg_127__3_ ( .D(n19604), .CP(wclk), .Q(ram[15363]) );
  DFF ram_reg_127__2_ ( .D(n19603), .CP(wclk), .Q(ram[15362]) );
  DFF ram_reg_127__1_ ( .D(n19602), .CP(wclk), .Q(ram[15361]) );
  DFF ram_reg_127__0_ ( .D(n19601), .CP(wclk), .Q(ram[15360]) );
  DFF ram_reg_135__7_ ( .D(n19544), .CP(wclk), .Q(ram[15303]) );
  DFF ram_reg_135__6_ ( .D(n19543), .CP(wclk), .Q(ram[15302]) );
  DFF ram_reg_135__5_ ( .D(n19542), .CP(wclk), .Q(ram[15301]) );
  DFF ram_reg_135__4_ ( .D(n19541), .CP(wclk), .Q(ram[15300]) );
  DFF ram_reg_135__3_ ( .D(n19540), .CP(wclk), .Q(ram[15299]) );
  DFF ram_reg_135__2_ ( .D(n19539), .CP(wclk), .Q(ram[15298]) );
  DFF ram_reg_135__1_ ( .D(n19538), .CP(wclk), .Q(ram[15297]) );
  DFF ram_reg_135__0_ ( .D(n19537), .CP(wclk), .Q(ram[15296]) );
  DFF ram_reg_147__7_ ( .D(n19448), .CP(wclk), .Q(ram[15207]) );
  DFF ram_reg_147__6_ ( .D(n19447), .CP(wclk), .Q(ram[15206]) );
  DFF ram_reg_147__5_ ( .D(n19446), .CP(wclk), .Q(ram[15205]) );
  DFF ram_reg_147__4_ ( .D(n19445), .CP(wclk), .Q(ram[15204]) );
  DFF ram_reg_147__3_ ( .D(n19444), .CP(wclk), .Q(ram[15203]) );
  DFF ram_reg_147__2_ ( .D(n19443), .CP(wclk), .Q(ram[15202]) );
  DFF ram_reg_147__1_ ( .D(n19442), .CP(wclk), .Q(ram[15201]) );
  DFF ram_reg_147__0_ ( .D(n19441), .CP(wclk), .Q(ram[15200]) );
  DFF ram_reg_151__7_ ( .D(n19416), .CP(wclk), .Q(ram[15175]) );
  DFF ram_reg_151__6_ ( .D(n19415), .CP(wclk), .Q(ram[15174]) );
  DFF ram_reg_151__5_ ( .D(n19414), .CP(wclk), .Q(ram[15173]) );
  DFF ram_reg_151__4_ ( .D(n19413), .CP(wclk), .Q(ram[15172]) );
  DFF ram_reg_151__3_ ( .D(n19412), .CP(wclk), .Q(ram[15171]) );
  DFF ram_reg_151__2_ ( .D(n19411), .CP(wclk), .Q(ram[15170]) );
  DFF ram_reg_151__1_ ( .D(n19410), .CP(wclk), .Q(ram[15169]) );
  DFF ram_reg_151__0_ ( .D(n19409), .CP(wclk), .Q(ram[15168]) );
  DFF ram_reg_167__7_ ( .D(n19288), .CP(wclk), .Q(ram[15047]) );
  DFF ram_reg_167__6_ ( .D(n19287), .CP(wclk), .Q(ram[15046]) );
  DFF ram_reg_167__5_ ( .D(n19286), .CP(wclk), .Q(ram[15045]) );
  DFF ram_reg_167__4_ ( .D(n19285), .CP(wclk), .Q(ram[15044]) );
  DFF ram_reg_167__3_ ( .D(n19284), .CP(wclk), .Q(ram[15043]) );
  DFF ram_reg_167__2_ ( .D(n19283), .CP(wclk), .Q(ram[15042]) );
  DFF ram_reg_167__1_ ( .D(n19282), .CP(wclk), .Q(ram[15041]) );
  DFF ram_reg_167__0_ ( .D(n19281), .CP(wclk), .Q(ram[15040]) );
  DFF ram_reg_195__7_ ( .D(n19064), .CP(wclk), .Q(ram[14823]) );
  DFF ram_reg_195__6_ ( .D(n19063), .CP(wclk), .Q(ram[14822]) );
  DFF ram_reg_195__5_ ( .D(n19062), .CP(wclk), .Q(ram[14821]) );
  DFF ram_reg_195__4_ ( .D(n19061), .CP(wclk), .Q(ram[14820]) );
  DFF ram_reg_195__3_ ( .D(n19060), .CP(wclk), .Q(ram[14819]) );
  DFF ram_reg_195__2_ ( .D(n19059), .CP(wclk), .Q(ram[14818]) );
  DFF ram_reg_195__1_ ( .D(n19058), .CP(wclk), .Q(ram[14817]) );
  DFF ram_reg_195__0_ ( .D(n19057), .CP(wclk), .Q(ram[14816]) );
  DFF ram_reg_199__7_ ( .D(n19032), .CP(wclk), .Q(ram[14791]) );
  DFF ram_reg_199__6_ ( .D(n19031), .CP(wclk), .Q(ram[14790]) );
  DFF ram_reg_199__5_ ( .D(n19030), .CP(wclk), .Q(ram[14789]) );
  DFF ram_reg_199__4_ ( .D(n19029), .CP(wclk), .Q(ram[14788]) );
  DFF ram_reg_199__3_ ( .D(n19028), .CP(wclk), .Q(ram[14787]) );
  DFF ram_reg_199__2_ ( .D(n19027), .CP(wclk), .Q(ram[14786]) );
  DFF ram_reg_199__1_ ( .D(n19026), .CP(wclk), .Q(ram[14785]) );
  DFF ram_reg_199__0_ ( .D(n19025), .CP(wclk), .Q(ram[14784]) );
  DFF ram_reg_211__7_ ( .D(n18936), .CP(wclk), .Q(ram[14695]) );
  DFF ram_reg_211__6_ ( .D(n18935), .CP(wclk), .Q(ram[14694]) );
  DFF ram_reg_211__5_ ( .D(n18934), .CP(wclk), .Q(ram[14693]) );
  DFF ram_reg_211__4_ ( .D(n18933), .CP(wclk), .Q(ram[14692]) );
  DFF ram_reg_211__3_ ( .D(n18932), .CP(wclk), .Q(ram[14691]) );
  DFF ram_reg_211__2_ ( .D(n18931), .CP(wclk), .Q(ram[14690]) );
  DFF ram_reg_211__1_ ( .D(n18930), .CP(wclk), .Q(ram[14689]) );
  DFF ram_reg_211__0_ ( .D(n18929), .CP(wclk), .Q(ram[14688]) );
  DFF ram_reg_215__7_ ( .D(n18904), .CP(wclk), .Q(ram[14663]) );
  DFF ram_reg_215__6_ ( .D(n18903), .CP(wclk), .Q(ram[14662]) );
  DFF ram_reg_215__5_ ( .D(n18902), .CP(wclk), .Q(ram[14661]) );
  DFF ram_reg_215__4_ ( .D(n18901), .CP(wclk), .Q(ram[14660]) );
  DFF ram_reg_215__3_ ( .D(n18900), .CP(wclk), .Q(ram[14659]) );
  DFF ram_reg_215__2_ ( .D(n18899), .CP(wclk), .Q(ram[14658]) );
  DFF ram_reg_215__1_ ( .D(n18898), .CP(wclk), .Q(ram[14657]) );
  DFF ram_reg_215__0_ ( .D(n18897), .CP(wclk), .Q(ram[14656]) );
  DFF ram_reg_231__7_ ( .D(n18776), .CP(wclk), .Q(ram[14535]) );
  DFF ram_reg_231__6_ ( .D(n18775), .CP(wclk), .Q(ram[14534]) );
  DFF ram_reg_231__5_ ( .D(n18774), .CP(wclk), .Q(ram[14533]) );
  DFF ram_reg_231__4_ ( .D(n18773), .CP(wclk), .Q(ram[14532]) );
  DFF ram_reg_231__3_ ( .D(n18772), .CP(wclk), .Q(ram[14531]) );
  DFF ram_reg_231__2_ ( .D(n18771), .CP(wclk), .Q(ram[14530]) );
  DFF ram_reg_231__1_ ( .D(n18770), .CP(wclk), .Q(ram[14529]) );
  DFF ram_reg_231__0_ ( .D(n18769), .CP(wclk), .Q(ram[14528]) );
  DFF ram_reg_247__7_ ( .D(n18648), .CP(wclk), .Q(ram[14407]) );
  DFF ram_reg_247__6_ ( .D(n18647), .CP(wclk), .Q(ram[14406]) );
  DFF ram_reg_247__5_ ( .D(n18646), .CP(wclk), .Q(ram[14405]) );
  DFF ram_reg_247__4_ ( .D(n18645), .CP(wclk), .Q(ram[14404]) );
  DFF ram_reg_247__3_ ( .D(n18644), .CP(wclk), .Q(ram[14403]) );
  DFF ram_reg_247__2_ ( .D(n18643), .CP(wclk), .Q(ram[14402]) );
  DFF ram_reg_247__1_ ( .D(n18642), .CP(wclk), .Q(ram[14401]) );
  DFF ram_reg_247__0_ ( .D(n18641), .CP(wclk), .Q(ram[14400]) );
  DFF ram_reg_259__7_ ( .D(n18552), .CP(wclk), .Q(ram[14311]) );
  DFF ram_reg_259__6_ ( .D(n18551), .CP(wclk), .Q(ram[14310]) );
  DFF ram_reg_259__5_ ( .D(n18550), .CP(wclk), .Q(ram[14309]) );
  DFF ram_reg_259__4_ ( .D(n18549), .CP(wclk), .Q(ram[14308]) );
  DFF ram_reg_259__3_ ( .D(n18548), .CP(wclk), .Q(ram[14307]) );
  DFF ram_reg_259__2_ ( .D(n18547), .CP(wclk), .Q(ram[14306]) );
  DFF ram_reg_259__1_ ( .D(n18546), .CP(wclk), .Q(ram[14305]) );
  DFF ram_reg_259__0_ ( .D(n18545), .CP(wclk), .Q(ram[14304]) );
  DFF ram_reg_263__7_ ( .D(n18520), .CP(wclk), .Q(ram[14279]) );
  DFF ram_reg_263__6_ ( .D(n18519), .CP(wclk), .Q(ram[14278]) );
  DFF ram_reg_263__5_ ( .D(n18518), .CP(wclk), .Q(ram[14277]) );
  DFF ram_reg_263__4_ ( .D(n18517), .CP(wclk), .Q(ram[14276]) );
  DFF ram_reg_263__3_ ( .D(n18516), .CP(wclk), .Q(ram[14275]) );
  DFF ram_reg_263__2_ ( .D(n18515), .CP(wclk), .Q(ram[14274]) );
  DFF ram_reg_263__1_ ( .D(n18514), .CP(wclk), .Q(ram[14273]) );
  DFF ram_reg_263__0_ ( .D(n18513), .CP(wclk), .Q(ram[14272]) );
  DFF ram_reg_275__7_ ( .D(n18424), .CP(wclk), .Q(ram[14183]) );
  DFF ram_reg_275__6_ ( .D(n18423), .CP(wclk), .Q(ram[14182]) );
  DFF ram_reg_275__5_ ( .D(n18422), .CP(wclk), .Q(ram[14181]) );
  DFF ram_reg_275__4_ ( .D(n18421), .CP(wclk), .Q(ram[14180]) );
  DFF ram_reg_275__3_ ( .D(n18420), .CP(wclk), .Q(ram[14179]) );
  DFF ram_reg_275__2_ ( .D(n18419), .CP(wclk), .Q(ram[14178]) );
  DFF ram_reg_275__1_ ( .D(n18418), .CP(wclk), .Q(ram[14177]) );
  DFF ram_reg_275__0_ ( .D(n18417), .CP(wclk), .Q(ram[14176]) );
  DFF ram_reg_279__7_ ( .D(n18392), .CP(wclk), .Q(ram[14151]) );
  DFF ram_reg_279__6_ ( .D(n18391), .CP(wclk), .Q(ram[14150]) );
  DFF ram_reg_279__5_ ( .D(n18390), .CP(wclk), .Q(ram[14149]) );
  DFF ram_reg_279__4_ ( .D(n18389), .CP(wclk), .Q(ram[14148]) );
  DFF ram_reg_279__3_ ( .D(n18388), .CP(wclk), .Q(ram[14147]) );
  DFF ram_reg_279__2_ ( .D(n18387), .CP(wclk), .Q(ram[14146]) );
  DFF ram_reg_279__1_ ( .D(n18386), .CP(wclk), .Q(ram[14145]) );
  DFF ram_reg_279__0_ ( .D(n18385), .CP(wclk), .Q(ram[14144]) );
  DFF ram_reg_287__7_ ( .D(n18328), .CP(wclk), .Q(ram[14087]) );
  DFF ram_reg_287__6_ ( .D(n18327), .CP(wclk), .Q(ram[14086]) );
  DFF ram_reg_287__5_ ( .D(n18326), .CP(wclk), .Q(ram[14085]) );
  DFF ram_reg_287__4_ ( .D(n18325), .CP(wclk), .Q(ram[14084]) );
  DFF ram_reg_287__3_ ( .D(n18324), .CP(wclk), .Q(ram[14083]) );
  DFF ram_reg_287__2_ ( .D(n18323), .CP(wclk), .Q(ram[14082]) );
  DFF ram_reg_287__1_ ( .D(n18322), .CP(wclk), .Q(ram[14081]) );
  DFF ram_reg_287__0_ ( .D(n18321), .CP(wclk), .Q(ram[14080]) );
  DFF ram_reg_291__7_ ( .D(n18296), .CP(wclk), .Q(ram[14055]) );
  DFF ram_reg_291__6_ ( .D(n18295), .CP(wclk), .Q(ram[14054]) );
  DFF ram_reg_291__5_ ( .D(n18294), .CP(wclk), .Q(ram[14053]) );
  DFF ram_reg_291__4_ ( .D(n18293), .CP(wclk), .Q(ram[14052]) );
  DFF ram_reg_291__3_ ( .D(n18292), .CP(wclk), .Q(ram[14051]) );
  DFF ram_reg_291__2_ ( .D(n18291), .CP(wclk), .Q(ram[14050]) );
  DFF ram_reg_291__1_ ( .D(n18290), .CP(wclk), .Q(ram[14049]) );
  DFF ram_reg_291__0_ ( .D(n18289), .CP(wclk), .Q(ram[14048]) );
  DFF ram_reg_295__7_ ( .D(n18264), .CP(wclk), .Q(ram[14023]) );
  DFF ram_reg_295__6_ ( .D(n18263), .CP(wclk), .Q(ram[14022]) );
  DFF ram_reg_295__5_ ( .D(n18262), .CP(wclk), .Q(ram[14021]) );
  DFF ram_reg_295__4_ ( .D(n18261), .CP(wclk), .Q(ram[14020]) );
  DFF ram_reg_295__3_ ( .D(n18260), .CP(wclk), .Q(ram[14019]) );
  DFF ram_reg_295__2_ ( .D(n18259), .CP(wclk), .Q(ram[14018]) );
  DFF ram_reg_295__1_ ( .D(n18258), .CP(wclk), .Q(ram[14017]) );
  DFF ram_reg_295__0_ ( .D(n18257), .CP(wclk), .Q(ram[14016]) );
  DFF ram_reg_307__7_ ( .D(n18168), .CP(wclk), .Q(ram[13927]) );
  DFF ram_reg_307__6_ ( .D(n18167), .CP(wclk), .Q(ram[13926]) );
  DFF ram_reg_307__5_ ( .D(n18166), .CP(wclk), .Q(ram[13925]) );
  DFF ram_reg_307__4_ ( .D(n18165), .CP(wclk), .Q(ram[13924]) );
  DFF ram_reg_307__3_ ( .D(n18164), .CP(wclk), .Q(ram[13923]) );
  DFF ram_reg_307__2_ ( .D(n18163), .CP(wclk), .Q(ram[13922]) );
  DFF ram_reg_307__1_ ( .D(n18162), .CP(wclk), .Q(ram[13921]) );
  DFF ram_reg_307__0_ ( .D(n18161), .CP(wclk), .Q(ram[13920]) );
  DFF ram_reg_311__7_ ( .D(n18136), .CP(wclk), .Q(ram[13895]) );
  DFF ram_reg_311__6_ ( .D(n18135), .CP(wclk), .Q(ram[13894]) );
  DFF ram_reg_311__5_ ( .D(n18134), .CP(wclk), .Q(ram[13893]) );
  DFF ram_reg_311__4_ ( .D(n18133), .CP(wclk), .Q(ram[13892]) );
  DFF ram_reg_311__3_ ( .D(n18132), .CP(wclk), .Q(ram[13891]) );
  DFF ram_reg_311__2_ ( .D(n18131), .CP(wclk), .Q(ram[13890]) );
  DFF ram_reg_311__1_ ( .D(n18130), .CP(wclk), .Q(ram[13889]) );
  DFF ram_reg_311__0_ ( .D(n18129), .CP(wclk), .Q(ram[13888]) );
  DFF ram_reg_323__7_ ( .D(n18040), .CP(wclk), .Q(ram[13799]) );
  DFF ram_reg_323__6_ ( .D(n18039), .CP(wclk), .Q(ram[13798]) );
  DFF ram_reg_323__5_ ( .D(n18038), .CP(wclk), .Q(ram[13797]) );
  DFF ram_reg_323__4_ ( .D(n18037), .CP(wclk), .Q(ram[13796]) );
  DFF ram_reg_323__3_ ( .D(n18036), .CP(wclk), .Q(ram[13795]) );
  DFF ram_reg_323__2_ ( .D(n18035), .CP(wclk), .Q(ram[13794]) );
  DFF ram_reg_323__1_ ( .D(n18034), .CP(wclk), .Q(ram[13793]) );
  DFF ram_reg_323__0_ ( .D(n18033), .CP(wclk), .Q(ram[13792]) );
  DFF ram_reg_327__7_ ( .D(n18008), .CP(wclk), .Q(ram[13767]) );
  DFF ram_reg_327__6_ ( .D(n18007), .CP(wclk), .Q(ram[13766]) );
  DFF ram_reg_327__5_ ( .D(n18006), .CP(wclk), .Q(ram[13765]) );
  DFF ram_reg_327__4_ ( .D(n18005), .CP(wclk), .Q(ram[13764]) );
  DFF ram_reg_327__3_ ( .D(n18004), .CP(wclk), .Q(ram[13763]) );
  DFF ram_reg_327__2_ ( .D(n18003), .CP(wclk), .Q(ram[13762]) );
  DFF ram_reg_327__1_ ( .D(n18002), .CP(wclk), .Q(ram[13761]) );
  DFF ram_reg_327__0_ ( .D(n18001), .CP(wclk), .Q(ram[13760]) );
  DFF ram_reg_331__7_ ( .D(n17976), .CP(wclk), .Q(ram[13735]) );
  DFF ram_reg_331__6_ ( .D(n17975), .CP(wclk), .Q(ram[13734]) );
  DFF ram_reg_331__5_ ( .D(n17974), .CP(wclk), .Q(ram[13733]) );
  DFF ram_reg_331__4_ ( .D(n17973), .CP(wclk), .Q(ram[13732]) );
  DFF ram_reg_331__3_ ( .D(n17972), .CP(wclk), .Q(ram[13731]) );
  DFF ram_reg_331__2_ ( .D(n17971), .CP(wclk), .Q(ram[13730]) );
  DFF ram_reg_331__1_ ( .D(n17970), .CP(wclk), .Q(ram[13729]) );
  DFF ram_reg_331__0_ ( .D(n17969), .CP(wclk), .Q(ram[13728]) );
  DFF ram_reg_335__7_ ( .D(n17944), .CP(wclk), .Q(ram[13703]) );
  DFF ram_reg_335__6_ ( .D(n17943), .CP(wclk), .Q(ram[13702]) );
  DFF ram_reg_335__5_ ( .D(n17942), .CP(wclk), .Q(ram[13701]) );
  DFF ram_reg_335__4_ ( .D(n17941), .CP(wclk), .Q(ram[13700]) );
  DFF ram_reg_335__3_ ( .D(n17940), .CP(wclk), .Q(ram[13699]) );
  DFF ram_reg_335__2_ ( .D(n17939), .CP(wclk), .Q(ram[13698]) );
  DFF ram_reg_335__1_ ( .D(n17938), .CP(wclk), .Q(ram[13697]) );
  DFF ram_reg_335__0_ ( .D(n17937), .CP(wclk), .Q(ram[13696]) );
  DFF ram_reg_339__7_ ( .D(n17912), .CP(wclk), .Q(ram[13671]) );
  DFF ram_reg_339__6_ ( .D(n17911), .CP(wclk), .Q(ram[13670]) );
  DFF ram_reg_339__5_ ( .D(n17910), .CP(wclk), .Q(ram[13669]) );
  DFF ram_reg_339__4_ ( .D(n17909), .CP(wclk), .Q(ram[13668]) );
  DFF ram_reg_339__3_ ( .D(n17908), .CP(wclk), .Q(ram[13667]) );
  DFF ram_reg_339__2_ ( .D(n17907), .CP(wclk), .Q(ram[13666]) );
  DFF ram_reg_339__1_ ( .D(n17906), .CP(wclk), .Q(ram[13665]) );
  DFF ram_reg_339__0_ ( .D(n17905), .CP(wclk), .Q(ram[13664]) );
  DFF ram_reg_343__7_ ( .D(n17880), .CP(wclk), .Q(ram[13639]) );
  DFF ram_reg_343__6_ ( .D(n17879), .CP(wclk), .Q(ram[13638]) );
  DFF ram_reg_343__5_ ( .D(n17878), .CP(wclk), .Q(ram[13637]) );
  DFF ram_reg_343__4_ ( .D(n17877), .CP(wclk), .Q(ram[13636]) );
  DFF ram_reg_343__3_ ( .D(n17876), .CP(wclk), .Q(ram[13635]) );
  DFF ram_reg_343__2_ ( .D(n17875), .CP(wclk), .Q(ram[13634]) );
  DFF ram_reg_343__1_ ( .D(n17874), .CP(wclk), .Q(ram[13633]) );
  DFF ram_reg_343__0_ ( .D(n17873), .CP(wclk), .Q(ram[13632]) );
  DFF ram_reg_347__7_ ( .D(n17848), .CP(wclk), .Q(ram[13607]) );
  DFF ram_reg_347__6_ ( .D(n17847), .CP(wclk), .Q(ram[13606]) );
  DFF ram_reg_347__5_ ( .D(n17846), .CP(wclk), .Q(ram[13605]) );
  DFF ram_reg_347__4_ ( .D(n17845), .CP(wclk), .Q(ram[13604]) );
  DFF ram_reg_347__3_ ( .D(n17844), .CP(wclk), .Q(ram[13603]) );
  DFF ram_reg_347__2_ ( .D(n17843), .CP(wclk), .Q(ram[13602]) );
  DFF ram_reg_347__1_ ( .D(n17842), .CP(wclk), .Q(ram[13601]) );
  DFF ram_reg_347__0_ ( .D(n17841), .CP(wclk), .Q(ram[13600]) );
  DFF ram_reg_351__7_ ( .D(n17816), .CP(wclk), .Q(ram[13575]) );
  DFF ram_reg_351__6_ ( .D(n17815), .CP(wclk), .Q(ram[13574]) );
  DFF ram_reg_351__5_ ( .D(n17814), .CP(wclk), .Q(ram[13573]) );
  DFF ram_reg_351__4_ ( .D(n17813), .CP(wclk), .Q(ram[13572]) );
  DFF ram_reg_351__3_ ( .D(n17812), .CP(wclk), .Q(ram[13571]) );
  DFF ram_reg_351__2_ ( .D(n17811), .CP(wclk), .Q(ram[13570]) );
  DFF ram_reg_351__1_ ( .D(n17810), .CP(wclk), .Q(ram[13569]) );
  DFF ram_reg_351__0_ ( .D(n17809), .CP(wclk), .Q(ram[13568]) );
  DFF ram_reg_355__7_ ( .D(n17784), .CP(wclk), .Q(ram[13543]) );
  DFF ram_reg_355__6_ ( .D(n17783), .CP(wclk), .Q(ram[13542]) );
  DFF ram_reg_355__5_ ( .D(n17782), .CP(wclk), .Q(ram[13541]) );
  DFF ram_reg_355__4_ ( .D(n17781), .CP(wclk), .Q(ram[13540]) );
  DFF ram_reg_355__3_ ( .D(n17780), .CP(wclk), .Q(ram[13539]) );
  DFF ram_reg_355__2_ ( .D(n17779), .CP(wclk), .Q(ram[13538]) );
  DFF ram_reg_355__1_ ( .D(n17778), .CP(wclk), .Q(ram[13537]) );
  DFF ram_reg_355__0_ ( .D(n17777), .CP(wclk), .Q(ram[13536]) );
  DFF ram_reg_359__7_ ( .D(n17752), .CP(wclk), .Q(ram[13511]) );
  DFF ram_reg_359__6_ ( .D(n17751), .CP(wclk), .Q(ram[13510]) );
  DFF ram_reg_359__5_ ( .D(n17750), .CP(wclk), .Q(ram[13509]) );
  DFF ram_reg_359__4_ ( .D(n17749), .CP(wclk), .Q(ram[13508]) );
  DFF ram_reg_359__3_ ( .D(n17748), .CP(wclk), .Q(ram[13507]) );
  DFF ram_reg_359__2_ ( .D(n17747), .CP(wclk), .Q(ram[13506]) );
  DFF ram_reg_359__1_ ( .D(n17746), .CP(wclk), .Q(ram[13505]) );
  DFF ram_reg_359__0_ ( .D(n17745), .CP(wclk), .Q(ram[13504]) );
  DFF ram_reg_367__7_ ( .D(n17688), .CP(wclk), .Q(ram[13447]) );
  DFF ram_reg_367__6_ ( .D(n17687), .CP(wclk), .Q(ram[13446]) );
  DFF ram_reg_367__5_ ( .D(n17686), .CP(wclk), .Q(ram[13445]) );
  DFF ram_reg_367__4_ ( .D(n17685), .CP(wclk), .Q(ram[13444]) );
  DFF ram_reg_367__3_ ( .D(n17684), .CP(wclk), .Q(ram[13443]) );
  DFF ram_reg_367__2_ ( .D(n17683), .CP(wclk), .Q(ram[13442]) );
  DFF ram_reg_367__1_ ( .D(n17682), .CP(wclk), .Q(ram[13441]) );
  DFF ram_reg_367__0_ ( .D(n17681), .CP(wclk), .Q(ram[13440]) );
  DFF ram_reg_371__7_ ( .D(n17656), .CP(wclk), .Q(ram[13415]) );
  DFF ram_reg_371__6_ ( .D(n17655), .CP(wclk), .Q(ram[13414]) );
  DFF ram_reg_371__5_ ( .D(n17654), .CP(wclk), .Q(ram[13413]) );
  DFF ram_reg_371__4_ ( .D(n17653), .CP(wclk), .Q(ram[13412]) );
  DFF ram_reg_371__3_ ( .D(n17652), .CP(wclk), .Q(ram[13411]) );
  DFF ram_reg_371__2_ ( .D(n17651), .CP(wclk), .Q(ram[13410]) );
  DFF ram_reg_371__1_ ( .D(n17650), .CP(wclk), .Q(ram[13409]) );
  DFF ram_reg_371__0_ ( .D(n17649), .CP(wclk), .Q(ram[13408]) );
  DFF ram_reg_375__7_ ( .D(n17624), .CP(wclk), .Q(ram[13383]) );
  DFF ram_reg_375__6_ ( .D(n17623), .CP(wclk), .Q(ram[13382]) );
  DFF ram_reg_375__5_ ( .D(n17622), .CP(wclk), .Q(ram[13381]) );
  DFF ram_reg_375__4_ ( .D(n17621), .CP(wclk), .Q(ram[13380]) );
  DFF ram_reg_375__3_ ( .D(n17620), .CP(wclk), .Q(ram[13379]) );
  DFF ram_reg_375__2_ ( .D(n17619), .CP(wclk), .Q(ram[13378]) );
  DFF ram_reg_375__1_ ( .D(n17618), .CP(wclk), .Q(ram[13377]) );
  DFF ram_reg_375__0_ ( .D(n17617), .CP(wclk), .Q(ram[13376]) );
  DFF ram_reg_383__7_ ( .D(n17560), .CP(wclk), .Q(ram[13319]) );
  DFF ram_reg_383__6_ ( .D(n17559), .CP(wclk), .Q(ram[13318]) );
  DFF ram_reg_383__5_ ( .D(n17558), .CP(wclk), .Q(ram[13317]) );
  DFF ram_reg_383__4_ ( .D(n17557), .CP(wclk), .Q(ram[13316]) );
  DFF ram_reg_383__3_ ( .D(n17556), .CP(wclk), .Q(ram[13315]) );
  DFF ram_reg_383__2_ ( .D(n17555), .CP(wclk), .Q(ram[13314]) );
  DFF ram_reg_383__1_ ( .D(n17554), .CP(wclk), .Q(ram[13313]) );
  DFF ram_reg_383__0_ ( .D(n17553), .CP(wclk), .Q(ram[13312]) );
  DFF ram_reg_391__7_ ( .D(n17496), .CP(wclk), .Q(ram[13255]) );
  DFF ram_reg_391__6_ ( .D(n17495), .CP(wclk), .Q(ram[13254]) );
  DFF ram_reg_391__5_ ( .D(n17494), .CP(wclk), .Q(ram[13253]) );
  DFF ram_reg_391__4_ ( .D(n17493), .CP(wclk), .Q(ram[13252]) );
  DFF ram_reg_391__3_ ( .D(n17492), .CP(wclk), .Q(ram[13251]) );
  DFF ram_reg_391__2_ ( .D(n17491), .CP(wclk), .Q(ram[13250]) );
  DFF ram_reg_391__1_ ( .D(n17490), .CP(wclk), .Q(ram[13249]) );
  DFF ram_reg_391__0_ ( .D(n17489), .CP(wclk), .Q(ram[13248]) );
  DFF ram_reg_407__7_ ( .D(n17368), .CP(wclk), .Q(ram[13127]) );
  DFF ram_reg_407__6_ ( .D(n17367), .CP(wclk), .Q(ram[13126]) );
  DFF ram_reg_407__5_ ( .D(n17366), .CP(wclk), .Q(ram[13125]) );
  DFF ram_reg_407__4_ ( .D(n17365), .CP(wclk), .Q(ram[13124]) );
  DFF ram_reg_407__3_ ( .D(n17364), .CP(wclk), .Q(ram[13123]) );
  DFF ram_reg_407__2_ ( .D(n17363), .CP(wclk), .Q(ram[13122]) );
  DFF ram_reg_407__1_ ( .D(n17362), .CP(wclk), .Q(ram[13121]) );
  DFF ram_reg_407__0_ ( .D(n17361), .CP(wclk), .Q(ram[13120]) );
  DFF ram_reg_455__7_ ( .D(n16984), .CP(wclk), .Q(ram[12743]) );
  DFF ram_reg_455__6_ ( .D(n16983), .CP(wclk), .Q(ram[12742]) );
  DFF ram_reg_455__5_ ( .D(n16982), .CP(wclk), .Q(ram[12741]) );
  DFF ram_reg_455__4_ ( .D(n16981), .CP(wclk), .Q(ram[12740]) );
  DFF ram_reg_455__3_ ( .D(n16980), .CP(wclk), .Q(ram[12739]) );
  DFF ram_reg_455__2_ ( .D(n16979), .CP(wclk), .Q(ram[12738]) );
  DFF ram_reg_455__1_ ( .D(n16978), .CP(wclk), .Q(ram[12737]) );
  DFF ram_reg_455__0_ ( .D(n16977), .CP(wclk), .Q(ram[12736]) );
  DFF ram_reg_467__7_ ( .D(n16888), .CP(wclk), .Q(ram[12647]) );
  DFF ram_reg_467__6_ ( .D(n16887), .CP(wclk), .Q(ram[12646]) );
  DFF ram_reg_467__5_ ( .D(n16886), .CP(wclk), .Q(ram[12645]) );
  DFF ram_reg_467__4_ ( .D(n16885), .CP(wclk), .Q(ram[12644]) );
  DFF ram_reg_467__3_ ( .D(n16884), .CP(wclk), .Q(ram[12643]) );
  DFF ram_reg_467__2_ ( .D(n16883), .CP(wclk), .Q(ram[12642]) );
  DFF ram_reg_467__1_ ( .D(n16882), .CP(wclk), .Q(ram[12641]) );
  DFF ram_reg_467__0_ ( .D(n16881), .CP(wclk), .Q(ram[12640]) );
  DFF ram_reg_471__7_ ( .D(n16856), .CP(wclk), .Q(ram[12615]) );
  DFF ram_reg_471__6_ ( .D(n16855), .CP(wclk), .Q(ram[12614]) );
  DFF ram_reg_471__5_ ( .D(n16854), .CP(wclk), .Q(ram[12613]) );
  DFF ram_reg_471__4_ ( .D(n16853), .CP(wclk), .Q(ram[12612]) );
  DFF ram_reg_471__3_ ( .D(n16852), .CP(wclk), .Q(ram[12611]) );
  DFF ram_reg_471__2_ ( .D(n16851), .CP(wclk), .Q(ram[12610]) );
  DFF ram_reg_471__1_ ( .D(n16850), .CP(wclk), .Q(ram[12609]) );
  DFF ram_reg_471__0_ ( .D(n16849), .CP(wclk), .Q(ram[12608]) );
  DFF ram_reg_487__7_ ( .D(n16728), .CP(wclk), .Q(ram[12487]) );
  DFF ram_reg_487__6_ ( .D(n16727), .CP(wclk), .Q(ram[12486]) );
  DFF ram_reg_487__5_ ( .D(n16726), .CP(wclk), .Q(ram[12485]) );
  DFF ram_reg_487__4_ ( .D(n16725), .CP(wclk), .Q(ram[12484]) );
  DFF ram_reg_487__3_ ( .D(n16724), .CP(wclk), .Q(ram[12483]) );
  DFF ram_reg_487__2_ ( .D(n16723), .CP(wclk), .Q(ram[12482]) );
  DFF ram_reg_487__1_ ( .D(n16722), .CP(wclk), .Q(ram[12481]) );
  DFF ram_reg_487__0_ ( .D(n16721), .CP(wclk), .Q(ram[12480]) );
  DFF ram_reg_503__7_ ( .D(n16600), .CP(wclk), .Q(ram[12359]) );
  DFF ram_reg_503__6_ ( .D(n16599), .CP(wclk), .Q(ram[12358]) );
  DFF ram_reg_503__5_ ( .D(n16598), .CP(wclk), .Q(ram[12357]) );
  DFF ram_reg_503__4_ ( .D(n16597), .CP(wclk), .Q(ram[12356]) );
  DFF ram_reg_503__3_ ( .D(n16596), .CP(wclk), .Q(ram[12355]) );
  DFF ram_reg_503__2_ ( .D(n16595), .CP(wclk), .Q(ram[12354]) );
  DFF ram_reg_503__1_ ( .D(n16594), .CP(wclk), .Q(ram[12353]) );
  DFF ram_reg_503__0_ ( .D(n16593), .CP(wclk), .Q(ram[12352]) );
  DFF ram_reg_515__7_ ( .D(n16504), .CP(wclk), .Q(ram[12263]) );
  DFF ram_reg_515__6_ ( .D(n16503), .CP(wclk), .Q(ram[12262]) );
  DFF ram_reg_515__5_ ( .D(n16502), .CP(wclk), .Q(ram[12261]) );
  DFF ram_reg_515__4_ ( .D(n16501), .CP(wclk), .Q(ram[12260]) );
  DFF ram_reg_515__3_ ( .D(n16500), .CP(wclk), .Q(ram[12259]) );
  DFF ram_reg_515__2_ ( .D(n16499), .CP(wclk), .Q(ram[12258]) );
  DFF ram_reg_515__1_ ( .D(n16498), .CP(wclk), .Q(ram[12257]) );
  DFF ram_reg_515__0_ ( .D(n16497), .CP(wclk), .Q(ram[12256]) );
  DFF ram_reg_519__7_ ( .D(n16472), .CP(wclk), .Q(ram[12231]) );
  DFF ram_reg_519__6_ ( .D(n16471), .CP(wclk), .Q(ram[12230]) );
  DFF ram_reg_519__5_ ( .D(n16470), .CP(wclk), .Q(ram[12229]) );
  DFF ram_reg_519__4_ ( .D(n16469), .CP(wclk), .Q(ram[12228]) );
  DFF ram_reg_519__3_ ( .D(n16468), .CP(wclk), .Q(ram[12227]) );
  DFF ram_reg_519__2_ ( .D(n16467), .CP(wclk), .Q(ram[12226]) );
  DFF ram_reg_519__1_ ( .D(n16466), .CP(wclk), .Q(ram[12225]) );
  DFF ram_reg_519__0_ ( .D(n16465), .CP(wclk), .Q(ram[12224]) );
  DFF ram_reg_531__7_ ( .D(n16376), .CP(wclk), .Q(ram[12135]) );
  DFF ram_reg_531__6_ ( .D(n16375), .CP(wclk), .Q(ram[12134]) );
  DFF ram_reg_531__5_ ( .D(n16374), .CP(wclk), .Q(ram[12133]) );
  DFF ram_reg_531__4_ ( .D(n16373), .CP(wclk), .Q(ram[12132]) );
  DFF ram_reg_531__3_ ( .D(n16372), .CP(wclk), .Q(ram[12131]) );
  DFF ram_reg_531__2_ ( .D(n16371), .CP(wclk), .Q(ram[12130]) );
  DFF ram_reg_531__1_ ( .D(n16370), .CP(wclk), .Q(ram[12129]) );
  DFF ram_reg_531__0_ ( .D(n16369), .CP(wclk), .Q(ram[12128]) );
  DFF ram_reg_535__7_ ( .D(n16344), .CP(wclk), .Q(ram[12103]) );
  DFF ram_reg_535__6_ ( .D(n16343), .CP(wclk), .Q(ram[12102]) );
  DFF ram_reg_535__5_ ( .D(n16342), .CP(wclk), .Q(ram[12101]) );
  DFF ram_reg_535__4_ ( .D(n16341), .CP(wclk), .Q(ram[12100]) );
  DFF ram_reg_535__3_ ( .D(n16340), .CP(wclk), .Q(ram[12099]) );
  DFF ram_reg_535__2_ ( .D(n16339), .CP(wclk), .Q(ram[12098]) );
  DFF ram_reg_535__1_ ( .D(n16338), .CP(wclk), .Q(ram[12097]) );
  DFF ram_reg_535__0_ ( .D(n16337), .CP(wclk), .Q(ram[12096]) );
  DFF ram_reg_551__7_ ( .D(n16216), .CP(wclk), .Q(ram[11975]) );
  DFF ram_reg_551__6_ ( .D(n16215), .CP(wclk), .Q(ram[11974]) );
  DFF ram_reg_551__5_ ( .D(n16214), .CP(wclk), .Q(ram[11973]) );
  DFF ram_reg_551__4_ ( .D(n16213), .CP(wclk), .Q(ram[11972]) );
  DFF ram_reg_551__3_ ( .D(n16212), .CP(wclk), .Q(ram[11971]) );
  DFF ram_reg_551__2_ ( .D(n16211), .CP(wclk), .Q(ram[11970]) );
  DFF ram_reg_551__1_ ( .D(n16210), .CP(wclk), .Q(ram[11969]) );
  DFF ram_reg_551__0_ ( .D(n16209), .CP(wclk), .Q(ram[11968]) );
  DFF ram_reg_567__7_ ( .D(n16088), .CP(wclk), .Q(ram[11847]) );
  DFF ram_reg_567__6_ ( .D(n16087), .CP(wclk), .Q(ram[11846]) );
  DFF ram_reg_567__5_ ( .D(n16086), .CP(wclk), .Q(ram[11845]) );
  DFF ram_reg_567__4_ ( .D(n16085), .CP(wclk), .Q(ram[11844]) );
  DFF ram_reg_567__3_ ( .D(n16084), .CP(wclk), .Q(ram[11843]) );
  DFF ram_reg_567__2_ ( .D(n16083), .CP(wclk), .Q(ram[11842]) );
  DFF ram_reg_567__1_ ( .D(n16082), .CP(wclk), .Q(ram[11841]) );
  DFF ram_reg_567__0_ ( .D(n16081), .CP(wclk), .Q(ram[11840]) );
  DFF ram_reg_579__7_ ( .D(n15992), .CP(wclk), .Q(ram[11751]) );
  DFF ram_reg_579__6_ ( .D(n15991), .CP(wclk), .Q(ram[11750]) );
  DFF ram_reg_579__5_ ( .D(n15990), .CP(wclk), .Q(ram[11749]) );
  DFF ram_reg_579__4_ ( .D(n15989), .CP(wclk), .Q(ram[11748]) );
  DFF ram_reg_579__3_ ( .D(n15988), .CP(wclk), .Q(ram[11747]) );
  DFF ram_reg_579__2_ ( .D(n15987), .CP(wclk), .Q(ram[11746]) );
  DFF ram_reg_579__1_ ( .D(n15986), .CP(wclk), .Q(ram[11745]) );
  DFF ram_reg_579__0_ ( .D(n15985), .CP(wclk), .Q(ram[11744]) );
  DFF ram_reg_583__7_ ( .D(n15960), .CP(wclk), .Q(ram[11719]) );
  DFF ram_reg_583__6_ ( .D(n15959), .CP(wclk), .Q(ram[11718]) );
  DFF ram_reg_583__5_ ( .D(n15958), .CP(wclk), .Q(ram[11717]) );
  DFF ram_reg_583__4_ ( .D(n15957), .CP(wclk), .Q(ram[11716]) );
  DFF ram_reg_583__3_ ( .D(n15956), .CP(wclk), .Q(ram[11715]) );
  DFF ram_reg_583__2_ ( .D(n15955), .CP(wclk), .Q(ram[11714]) );
  DFF ram_reg_583__1_ ( .D(n15954), .CP(wclk), .Q(ram[11713]) );
  DFF ram_reg_583__0_ ( .D(n15953), .CP(wclk), .Q(ram[11712]) );
  DFF ram_reg_591__7_ ( .D(n15896), .CP(wclk), .Q(ram[11655]) );
  DFF ram_reg_591__6_ ( .D(n15895), .CP(wclk), .Q(ram[11654]) );
  DFF ram_reg_591__5_ ( .D(n15894), .CP(wclk), .Q(ram[11653]) );
  DFF ram_reg_591__4_ ( .D(n15893), .CP(wclk), .Q(ram[11652]) );
  DFF ram_reg_591__3_ ( .D(n15892), .CP(wclk), .Q(ram[11651]) );
  DFF ram_reg_591__2_ ( .D(n15891), .CP(wclk), .Q(ram[11650]) );
  DFF ram_reg_591__1_ ( .D(n15890), .CP(wclk), .Q(ram[11649]) );
  DFF ram_reg_591__0_ ( .D(n15889), .CP(wclk), .Q(ram[11648]) );
  DFF ram_reg_595__7_ ( .D(n15864), .CP(wclk), .Q(ram[11623]) );
  DFF ram_reg_595__6_ ( .D(n15863), .CP(wclk), .Q(ram[11622]) );
  DFF ram_reg_595__5_ ( .D(n15862), .CP(wclk), .Q(ram[11621]) );
  DFF ram_reg_595__4_ ( .D(n15861), .CP(wclk), .Q(ram[11620]) );
  DFF ram_reg_595__3_ ( .D(n15860), .CP(wclk), .Q(ram[11619]) );
  DFF ram_reg_595__2_ ( .D(n15859), .CP(wclk), .Q(ram[11618]) );
  DFF ram_reg_595__1_ ( .D(n15858), .CP(wclk), .Q(ram[11617]) );
  DFF ram_reg_595__0_ ( .D(n15857), .CP(wclk), .Q(ram[11616]) );
  DFF ram_reg_599__7_ ( .D(n15832), .CP(wclk), .Q(ram[11591]) );
  DFF ram_reg_599__6_ ( .D(n15831), .CP(wclk), .Q(ram[11590]) );
  DFF ram_reg_599__5_ ( .D(n15830), .CP(wclk), .Q(ram[11589]) );
  DFF ram_reg_599__4_ ( .D(n15829), .CP(wclk), .Q(ram[11588]) );
  DFF ram_reg_599__3_ ( .D(n15828), .CP(wclk), .Q(ram[11587]) );
  DFF ram_reg_599__2_ ( .D(n15827), .CP(wclk), .Q(ram[11586]) );
  DFF ram_reg_599__1_ ( .D(n15826), .CP(wclk), .Q(ram[11585]) );
  DFF ram_reg_599__0_ ( .D(n15825), .CP(wclk), .Q(ram[11584]) );
  DFF ram_reg_603__7_ ( .D(n15800), .CP(wclk), .Q(ram[11559]) );
  DFF ram_reg_603__6_ ( .D(n15799), .CP(wclk), .Q(ram[11558]) );
  DFF ram_reg_603__5_ ( .D(n15798), .CP(wclk), .Q(ram[11557]) );
  DFF ram_reg_603__4_ ( .D(n15797), .CP(wclk), .Q(ram[11556]) );
  DFF ram_reg_603__3_ ( .D(n15796), .CP(wclk), .Q(ram[11555]) );
  DFF ram_reg_603__2_ ( .D(n15795), .CP(wclk), .Q(ram[11554]) );
  DFF ram_reg_603__1_ ( .D(n15794), .CP(wclk), .Q(ram[11553]) );
  DFF ram_reg_603__0_ ( .D(n15793), .CP(wclk), .Q(ram[11552]) );
  DFF ram_reg_607__7_ ( .D(n15768), .CP(wclk), .Q(ram[11527]) );
  DFF ram_reg_607__6_ ( .D(n15767), .CP(wclk), .Q(ram[11526]) );
  DFF ram_reg_607__5_ ( .D(n15766), .CP(wclk), .Q(ram[11525]) );
  DFF ram_reg_607__4_ ( .D(n15765), .CP(wclk), .Q(ram[11524]) );
  DFF ram_reg_607__3_ ( .D(n15764), .CP(wclk), .Q(ram[11523]) );
  DFF ram_reg_607__2_ ( .D(n15763), .CP(wclk), .Q(ram[11522]) );
  DFF ram_reg_607__1_ ( .D(n15762), .CP(wclk), .Q(ram[11521]) );
  DFF ram_reg_607__0_ ( .D(n15761), .CP(wclk), .Q(ram[11520]) );
  DFF ram_reg_611__7_ ( .D(n15736), .CP(wclk), .Q(ram[11495]) );
  DFF ram_reg_611__6_ ( .D(n15735), .CP(wclk), .Q(ram[11494]) );
  DFF ram_reg_611__5_ ( .D(n15734), .CP(wclk), .Q(ram[11493]) );
  DFF ram_reg_611__4_ ( .D(n15733), .CP(wclk), .Q(ram[11492]) );
  DFF ram_reg_611__3_ ( .D(n15732), .CP(wclk), .Q(ram[11491]) );
  DFF ram_reg_611__2_ ( .D(n15731), .CP(wclk), .Q(ram[11490]) );
  DFF ram_reg_611__1_ ( .D(n15730), .CP(wclk), .Q(ram[11489]) );
  DFF ram_reg_611__0_ ( .D(n15729), .CP(wclk), .Q(ram[11488]) );
  DFF ram_reg_615__7_ ( .D(n15704), .CP(wclk), .Q(ram[11463]) );
  DFF ram_reg_615__6_ ( .D(n15703), .CP(wclk), .Q(ram[11462]) );
  DFF ram_reg_615__5_ ( .D(n15702), .CP(wclk), .Q(ram[11461]) );
  DFF ram_reg_615__4_ ( .D(n15701), .CP(wclk), .Q(ram[11460]) );
  DFF ram_reg_615__3_ ( .D(n15700), .CP(wclk), .Q(ram[11459]) );
  DFF ram_reg_615__2_ ( .D(n15699), .CP(wclk), .Q(ram[11458]) );
  DFF ram_reg_615__1_ ( .D(n15698), .CP(wclk), .Q(ram[11457]) );
  DFF ram_reg_615__0_ ( .D(n15697), .CP(wclk), .Q(ram[11456]) );
  DFF ram_reg_627__7_ ( .D(n15608), .CP(wclk), .Q(ram[11367]) );
  DFF ram_reg_627__6_ ( .D(n15607), .CP(wclk), .Q(ram[11366]) );
  DFF ram_reg_627__5_ ( .D(n15606), .CP(wclk), .Q(ram[11365]) );
  DFF ram_reg_627__4_ ( .D(n15605), .CP(wclk), .Q(ram[11364]) );
  DFF ram_reg_627__3_ ( .D(n15604), .CP(wclk), .Q(ram[11363]) );
  DFF ram_reg_627__2_ ( .D(n15603), .CP(wclk), .Q(ram[11362]) );
  DFF ram_reg_627__1_ ( .D(n15602), .CP(wclk), .Q(ram[11361]) );
  DFF ram_reg_627__0_ ( .D(n15601), .CP(wclk), .Q(ram[11360]) );
  DFF ram_reg_631__7_ ( .D(n15576), .CP(wclk), .Q(ram[11335]) );
  DFF ram_reg_631__6_ ( .D(n15575), .CP(wclk), .Q(ram[11334]) );
  DFF ram_reg_631__5_ ( .D(n15574), .CP(wclk), .Q(ram[11333]) );
  DFF ram_reg_631__4_ ( .D(n15573), .CP(wclk), .Q(ram[11332]) );
  DFF ram_reg_631__3_ ( .D(n15572), .CP(wclk), .Q(ram[11331]) );
  DFF ram_reg_631__2_ ( .D(n15571), .CP(wclk), .Q(ram[11330]) );
  DFF ram_reg_631__1_ ( .D(n15570), .CP(wclk), .Q(ram[11329]) );
  DFF ram_reg_631__0_ ( .D(n15569), .CP(wclk), .Q(ram[11328]) );
  DFF ram_reg_663__7_ ( .D(n15320), .CP(wclk), .Q(ram[11079]) );
  DFF ram_reg_663__6_ ( .D(n15319), .CP(wclk), .Q(ram[11078]) );
  DFF ram_reg_663__5_ ( .D(n15318), .CP(wclk), .Q(ram[11077]) );
  DFF ram_reg_663__4_ ( .D(n15317), .CP(wclk), .Q(ram[11076]) );
  DFF ram_reg_663__3_ ( .D(n15316), .CP(wclk), .Q(ram[11075]) );
  DFF ram_reg_663__2_ ( .D(n15315), .CP(wclk), .Q(ram[11074]) );
  DFF ram_reg_663__1_ ( .D(n15314), .CP(wclk), .Q(ram[11073]) );
  DFF ram_reg_663__0_ ( .D(n15313), .CP(wclk), .Q(ram[11072]) );
  DFF ram_reg_711__7_ ( .D(n14936), .CP(wclk), .Q(ram[10695]) );
  DFF ram_reg_711__6_ ( .D(n14935), .CP(wclk), .Q(ram[10694]) );
  DFF ram_reg_711__5_ ( .D(n14934), .CP(wclk), .Q(ram[10693]) );
  DFF ram_reg_711__4_ ( .D(n14933), .CP(wclk), .Q(ram[10692]) );
  DFF ram_reg_711__3_ ( .D(n14932), .CP(wclk), .Q(ram[10691]) );
  DFF ram_reg_711__2_ ( .D(n14931), .CP(wclk), .Q(ram[10690]) );
  DFF ram_reg_711__1_ ( .D(n14930), .CP(wclk), .Q(ram[10689]) );
  DFF ram_reg_711__0_ ( .D(n14929), .CP(wclk), .Q(ram[10688]) );
  DFF ram_reg_727__7_ ( .D(n14808), .CP(wclk), .Q(ram[10567]) );
  DFF ram_reg_727__6_ ( .D(n14807), .CP(wclk), .Q(ram[10566]) );
  DFF ram_reg_727__5_ ( .D(n14806), .CP(wclk), .Q(ram[10565]) );
  DFF ram_reg_727__4_ ( .D(n14805), .CP(wclk), .Q(ram[10564]) );
  DFF ram_reg_727__3_ ( .D(n14804), .CP(wclk), .Q(ram[10563]) );
  DFF ram_reg_727__2_ ( .D(n14803), .CP(wclk), .Q(ram[10562]) );
  DFF ram_reg_727__1_ ( .D(n14802), .CP(wclk), .Q(ram[10561]) );
  DFF ram_reg_727__0_ ( .D(n14801), .CP(wclk), .Q(ram[10560]) );
  DFF ram_reg_775__7_ ( .D(n14424), .CP(wclk), .Q(ram[10183]) );
  DFF ram_reg_775__6_ ( .D(n14423), .CP(wclk), .Q(ram[10182]) );
  DFF ram_reg_775__5_ ( .D(n14422), .CP(wclk), .Q(ram[10181]) );
  DFF ram_reg_775__4_ ( .D(n14421), .CP(wclk), .Q(ram[10180]) );
  DFF ram_reg_775__3_ ( .D(n14420), .CP(wclk), .Q(ram[10179]) );
  DFF ram_reg_775__2_ ( .D(n14419), .CP(wclk), .Q(ram[10178]) );
  DFF ram_reg_775__1_ ( .D(n14418), .CP(wclk), .Q(ram[10177]) );
  DFF ram_reg_775__0_ ( .D(n14417), .CP(wclk), .Q(ram[10176]) );
  DFF ram_reg_787__7_ ( .D(n14328), .CP(wclk), .Q(ram[10087]) );
  DFF ram_reg_787__6_ ( .D(n14327), .CP(wclk), .Q(ram[10086]) );
  DFF ram_reg_787__5_ ( .D(n14326), .CP(wclk), .Q(ram[10085]) );
  DFF ram_reg_787__4_ ( .D(n14325), .CP(wclk), .Q(ram[10084]) );
  DFF ram_reg_787__3_ ( .D(n14324), .CP(wclk), .Q(ram[10083]) );
  DFF ram_reg_787__2_ ( .D(n14323), .CP(wclk), .Q(ram[10082]) );
  DFF ram_reg_787__1_ ( .D(n14322), .CP(wclk), .Q(ram[10081]) );
  DFF ram_reg_787__0_ ( .D(n14321), .CP(wclk), .Q(ram[10080]) );
  DFF ram_reg_791__7_ ( .D(n14296), .CP(wclk), .Q(ram[10055]) );
  DFF ram_reg_791__6_ ( .D(n14295), .CP(wclk), .Q(ram[10054]) );
  DFF ram_reg_791__5_ ( .D(n14294), .CP(wclk), .Q(ram[10053]) );
  DFF ram_reg_791__4_ ( .D(n14293), .CP(wclk), .Q(ram[10052]) );
  DFF ram_reg_791__3_ ( .D(n14292), .CP(wclk), .Q(ram[10051]) );
  DFF ram_reg_791__2_ ( .D(n14291), .CP(wclk), .Q(ram[10050]) );
  DFF ram_reg_791__1_ ( .D(n14290), .CP(wclk), .Q(ram[10049]) );
  DFF ram_reg_791__0_ ( .D(n14289), .CP(wclk), .Q(ram[10048]) );
  DFF ram_reg_807__7_ ( .D(n14168), .CP(wclk), .Q(ram[9927]) );
  DFF ram_reg_807__6_ ( .D(n14167), .CP(wclk), .Q(ram[9926]) );
  DFF ram_reg_807__5_ ( .D(n14166), .CP(wclk), .Q(ram[9925]) );
  DFF ram_reg_807__4_ ( .D(n14165), .CP(wclk), .Q(ram[9924]) );
  DFF ram_reg_807__3_ ( .D(n14164), .CP(wclk), .Q(ram[9923]) );
  DFF ram_reg_807__2_ ( .D(n14163), .CP(wclk), .Q(ram[9922]) );
  DFF ram_reg_807__1_ ( .D(n14162), .CP(wclk), .Q(ram[9921]) );
  DFF ram_reg_807__0_ ( .D(n14161), .CP(wclk), .Q(ram[9920]) );
  DFF ram_reg_823__7_ ( .D(n14040), .CP(wclk), .Q(ram[9799]) );
  DFF ram_reg_823__6_ ( .D(n14039), .CP(wclk), .Q(ram[9798]) );
  DFF ram_reg_823__5_ ( .D(n14038), .CP(wclk), .Q(ram[9797]) );
  DFF ram_reg_823__4_ ( .D(n14037), .CP(wclk), .Q(ram[9796]) );
  DFF ram_reg_823__3_ ( .D(n14036), .CP(wclk), .Q(ram[9795]) );
  DFF ram_reg_823__2_ ( .D(n14035), .CP(wclk), .Q(ram[9794]) );
  DFF ram_reg_823__1_ ( .D(n14034), .CP(wclk), .Q(ram[9793]) );
  DFF ram_reg_823__0_ ( .D(n14033), .CP(wclk), .Q(ram[9792]) );
  DFF ram_reg_835__7_ ( .D(n13944), .CP(wclk), .Q(ram[9703]) );
  DFF ram_reg_835__6_ ( .D(n13943), .CP(wclk), .Q(ram[9702]) );
  DFF ram_reg_835__5_ ( .D(n13942), .CP(wclk), .Q(ram[9701]) );
  DFF ram_reg_835__4_ ( .D(n13941), .CP(wclk), .Q(ram[9700]) );
  DFF ram_reg_835__3_ ( .D(n13940), .CP(wclk), .Q(ram[9699]) );
  DFF ram_reg_835__2_ ( .D(n13939), .CP(wclk), .Q(ram[9698]) );
  DFF ram_reg_835__1_ ( .D(n13938), .CP(wclk), .Q(ram[9697]) );
  DFF ram_reg_835__0_ ( .D(n13937), .CP(wclk), .Q(ram[9696]) );
  DFF ram_reg_839__7_ ( .D(n13912), .CP(wclk), .Q(ram[9671]) );
  DFF ram_reg_839__6_ ( .D(n13911), .CP(wclk), .Q(ram[9670]) );
  DFF ram_reg_839__5_ ( .D(n13910), .CP(wclk), .Q(ram[9669]) );
  DFF ram_reg_839__4_ ( .D(n13909), .CP(wclk), .Q(ram[9668]) );
  DFF ram_reg_839__3_ ( .D(n13908), .CP(wclk), .Q(ram[9667]) );
  DFF ram_reg_839__2_ ( .D(n13907), .CP(wclk), .Q(ram[9666]) );
  DFF ram_reg_839__1_ ( .D(n13906), .CP(wclk), .Q(ram[9665]) );
  DFF ram_reg_839__0_ ( .D(n13905), .CP(wclk), .Q(ram[9664]) );
  DFF ram_reg_847__7_ ( .D(n13848), .CP(wclk), .Q(ram[9607]) );
  DFF ram_reg_847__6_ ( .D(n13847), .CP(wclk), .Q(ram[9606]) );
  DFF ram_reg_847__5_ ( .D(n13846), .CP(wclk), .Q(ram[9605]) );
  DFF ram_reg_847__4_ ( .D(n13845), .CP(wclk), .Q(ram[9604]) );
  DFF ram_reg_847__3_ ( .D(n13844), .CP(wclk), .Q(ram[9603]) );
  DFF ram_reg_847__2_ ( .D(n13843), .CP(wclk), .Q(ram[9602]) );
  DFF ram_reg_847__1_ ( .D(n13842), .CP(wclk), .Q(ram[9601]) );
  DFF ram_reg_847__0_ ( .D(n13841), .CP(wclk), .Q(ram[9600]) );
  DFF ram_reg_851__7_ ( .D(n13816), .CP(wclk), .Q(ram[9575]) );
  DFF ram_reg_851__6_ ( .D(n13815), .CP(wclk), .Q(ram[9574]) );
  DFF ram_reg_851__5_ ( .D(n13814), .CP(wclk), .Q(ram[9573]) );
  DFF ram_reg_851__4_ ( .D(n13813), .CP(wclk), .Q(ram[9572]) );
  DFF ram_reg_851__3_ ( .D(n13812), .CP(wclk), .Q(ram[9571]) );
  DFF ram_reg_851__2_ ( .D(n13811), .CP(wclk), .Q(ram[9570]) );
  DFF ram_reg_851__1_ ( .D(n13810), .CP(wclk), .Q(ram[9569]) );
  DFF ram_reg_851__0_ ( .D(n13809), .CP(wclk), .Q(ram[9568]) );
  DFF ram_reg_855__7_ ( .D(n13784), .CP(wclk), .Q(ram[9543]) );
  DFF ram_reg_855__6_ ( .D(n13783), .CP(wclk), .Q(ram[9542]) );
  DFF ram_reg_855__5_ ( .D(n13782), .CP(wclk), .Q(ram[9541]) );
  DFF ram_reg_855__4_ ( .D(n13781), .CP(wclk), .Q(ram[9540]) );
  DFF ram_reg_855__3_ ( .D(n13780), .CP(wclk), .Q(ram[9539]) );
  DFF ram_reg_855__2_ ( .D(n13779), .CP(wclk), .Q(ram[9538]) );
  DFF ram_reg_855__1_ ( .D(n13778), .CP(wclk), .Q(ram[9537]) );
  DFF ram_reg_855__0_ ( .D(n13777), .CP(wclk), .Q(ram[9536]) );
  DFF ram_reg_863__7_ ( .D(n13720), .CP(wclk), .Q(ram[9479]) );
  DFF ram_reg_863__6_ ( .D(n13719), .CP(wclk), .Q(ram[9478]) );
  DFF ram_reg_863__5_ ( .D(n13718), .CP(wclk), .Q(ram[9477]) );
  DFF ram_reg_863__4_ ( .D(n13717), .CP(wclk), .Q(ram[9476]) );
  DFF ram_reg_863__3_ ( .D(n13716), .CP(wclk), .Q(ram[9475]) );
  DFF ram_reg_863__2_ ( .D(n13715), .CP(wclk), .Q(ram[9474]) );
  DFF ram_reg_863__1_ ( .D(n13714), .CP(wclk), .Q(ram[9473]) );
  DFF ram_reg_863__0_ ( .D(n13713), .CP(wclk), .Q(ram[9472]) );
  DFF ram_reg_867__7_ ( .D(n13688), .CP(wclk), .Q(ram[9447]) );
  DFF ram_reg_867__6_ ( .D(n13687), .CP(wclk), .Q(ram[9446]) );
  DFF ram_reg_867__5_ ( .D(n13686), .CP(wclk), .Q(ram[9445]) );
  DFF ram_reg_867__4_ ( .D(n13685), .CP(wclk), .Q(ram[9444]) );
  DFF ram_reg_867__3_ ( .D(n13684), .CP(wclk), .Q(ram[9443]) );
  DFF ram_reg_867__2_ ( .D(n13683), .CP(wclk), .Q(ram[9442]) );
  DFF ram_reg_867__1_ ( .D(n13682), .CP(wclk), .Q(ram[9441]) );
  DFF ram_reg_867__0_ ( .D(n13681), .CP(wclk), .Q(ram[9440]) );
  DFF ram_reg_871__7_ ( .D(n13656), .CP(wclk), .Q(ram[9415]) );
  DFF ram_reg_871__6_ ( .D(n13655), .CP(wclk), .Q(ram[9414]) );
  DFF ram_reg_871__5_ ( .D(n13654), .CP(wclk), .Q(ram[9413]) );
  DFF ram_reg_871__4_ ( .D(n13653), .CP(wclk), .Q(ram[9412]) );
  DFF ram_reg_871__3_ ( .D(n13652), .CP(wclk), .Q(ram[9411]) );
  DFF ram_reg_871__2_ ( .D(n13651), .CP(wclk), .Q(ram[9410]) );
  DFF ram_reg_871__1_ ( .D(n13650), .CP(wclk), .Q(ram[9409]) );
  DFF ram_reg_871__0_ ( .D(n13649), .CP(wclk), .Q(ram[9408]) );
  DFF ram_reg_883__7_ ( .D(n13560), .CP(wclk), .Q(ram[9319]) );
  DFF ram_reg_883__6_ ( .D(n13559), .CP(wclk), .Q(ram[9318]) );
  DFF ram_reg_883__5_ ( .D(n13558), .CP(wclk), .Q(ram[9317]) );
  DFF ram_reg_883__4_ ( .D(n13557), .CP(wclk), .Q(ram[9316]) );
  DFF ram_reg_883__3_ ( .D(n13556), .CP(wclk), .Q(ram[9315]) );
  DFF ram_reg_883__2_ ( .D(n13555), .CP(wclk), .Q(ram[9314]) );
  DFF ram_reg_883__1_ ( .D(n13554), .CP(wclk), .Q(ram[9313]) );
  DFF ram_reg_883__0_ ( .D(n13553), .CP(wclk), .Q(ram[9312]) );
  DFF ram_reg_887__7_ ( .D(n13528), .CP(wclk), .Q(ram[9287]) );
  DFF ram_reg_887__6_ ( .D(n13527), .CP(wclk), .Q(ram[9286]) );
  DFF ram_reg_887__5_ ( .D(n13526), .CP(wclk), .Q(ram[9285]) );
  DFF ram_reg_887__4_ ( .D(n13525), .CP(wclk), .Q(ram[9284]) );
  DFF ram_reg_887__3_ ( .D(n13524), .CP(wclk), .Q(ram[9283]) );
  DFF ram_reg_887__2_ ( .D(n13523), .CP(wclk), .Q(ram[9282]) );
  DFF ram_reg_887__1_ ( .D(n13522), .CP(wclk), .Q(ram[9281]) );
  DFF ram_reg_887__0_ ( .D(n13521), .CP(wclk), .Q(ram[9280]) );
  DFF ram_reg_967__7_ ( .D(n12888), .CP(wclk), .Q(ram[8647]) );
  DFF ram_reg_967__6_ ( .D(n12887), .CP(wclk), .Q(ram[8646]) );
  DFF ram_reg_967__5_ ( .D(n12886), .CP(wclk), .Q(ram[8645]) );
  DFF ram_reg_967__4_ ( .D(n12885), .CP(wclk), .Q(ram[8644]) );
  DFF ram_reg_967__3_ ( .D(n12884), .CP(wclk), .Q(ram[8643]) );
  DFF ram_reg_967__2_ ( .D(n12883), .CP(wclk), .Q(ram[8642]) );
  DFF ram_reg_967__1_ ( .D(n12882), .CP(wclk), .Q(ram[8641]) );
  DFF ram_reg_967__0_ ( .D(n12881), .CP(wclk), .Q(ram[8640]) );
  DFF ram_reg_983__7_ ( .D(n12760), .CP(wclk), .Q(ram[8519]) );
  DFF ram_reg_983__6_ ( .D(n12759), .CP(wclk), .Q(ram[8518]) );
  DFF ram_reg_983__5_ ( .D(n12758), .CP(wclk), .Q(ram[8517]) );
  DFF ram_reg_983__4_ ( .D(n12757), .CP(wclk), .Q(ram[8516]) );
  DFF ram_reg_983__3_ ( .D(n12756), .CP(wclk), .Q(ram[8515]) );
  DFF ram_reg_983__2_ ( .D(n12755), .CP(wclk), .Q(ram[8514]) );
  DFF ram_reg_983__1_ ( .D(n12754), .CP(wclk), .Q(ram[8513]) );
  DFF ram_reg_983__0_ ( .D(n12753), .CP(wclk), .Q(ram[8512]) );
  DFF ram_reg_1027__7_ ( .D(n12408), .CP(wclk), .Q(ram[8167]) );
  DFF ram_reg_1027__6_ ( .D(n12407), .CP(wclk), .Q(ram[8166]) );
  DFF ram_reg_1027__5_ ( .D(n12406), .CP(wclk), .Q(ram[8165]) );
  DFF ram_reg_1027__4_ ( .D(n12405), .CP(wclk), .Q(ram[8164]) );
  DFF ram_reg_1027__3_ ( .D(n12404), .CP(wclk), .Q(ram[8163]) );
  DFF ram_reg_1027__2_ ( .D(n12403), .CP(wclk), .Q(ram[8162]) );
  DFF ram_reg_1027__1_ ( .D(n12402), .CP(wclk), .Q(ram[8161]) );
  DFF ram_reg_1027__0_ ( .D(n12401), .CP(wclk), .Q(ram[8160]) );
  DFF ram_reg_1031__7_ ( .D(n12376), .CP(wclk), .Q(ram[8135]) );
  DFF ram_reg_1031__6_ ( .D(n12375), .CP(wclk), .Q(ram[8134]) );
  DFF ram_reg_1031__5_ ( .D(n12374), .CP(wclk), .Q(ram[8133]) );
  DFF ram_reg_1031__4_ ( .D(n12373), .CP(wclk), .Q(ram[8132]) );
  DFF ram_reg_1031__3_ ( .D(n12372), .CP(wclk), .Q(ram[8131]) );
  DFF ram_reg_1031__2_ ( .D(n12371), .CP(wclk), .Q(ram[8130]) );
  DFF ram_reg_1031__1_ ( .D(n12370), .CP(wclk), .Q(ram[8129]) );
  DFF ram_reg_1031__0_ ( .D(n12369), .CP(wclk), .Q(ram[8128]) );
  DFF ram_reg_1043__7_ ( .D(n12280), .CP(wclk), .Q(ram[8039]) );
  DFF ram_reg_1043__6_ ( .D(n12279), .CP(wclk), .Q(ram[8038]) );
  DFF ram_reg_1043__5_ ( .D(n12278), .CP(wclk), .Q(ram[8037]) );
  DFF ram_reg_1043__4_ ( .D(n12277), .CP(wclk), .Q(ram[8036]) );
  DFF ram_reg_1043__3_ ( .D(n12276), .CP(wclk), .Q(ram[8035]) );
  DFF ram_reg_1043__2_ ( .D(n12275), .CP(wclk), .Q(ram[8034]) );
  DFF ram_reg_1043__1_ ( .D(n12274), .CP(wclk), .Q(ram[8033]) );
  DFF ram_reg_1043__0_ ( .D(n12273), .CP(wclk), .Q(ram[8032]) );
  DFF ram_reg_1047__7_ ( .D(n12248), .CP(wclk), .Q(ram[8007]) );
  DFF ram_reg_1047__6_ ( .D(n12247), .CP(wclk), .Q(ram[8006]) );
  DFF ram_reg_1047__5_ ( .D(n12246), .CP(wclk), .Q(ram[8005]) );
  DFF ram_reg_1047__4_ ( .D(n12245), .CP(wclk), .Q(ram[8004]) );
  DFF ram_reg_1047__3_ ( .D(n12244), .CP(wclk), .Q(ram[8003]) );
  DFF ram_reg_1047__2_ ( .D(n12243), .CP(wclk), .Q(ram[8002]) );
  DFF ram_reg_1047__1_ ( .D(n12242), .CP(wclk), .Q(ram[8001]) );
  DFF ram_reg_1047__0_ ( .D(n12241), .CP(wclk), .Q(ram[8000]) );
  DFF ram_reg_1055__7_ ( .D(n12184), .CP(wclk), .Q(ram[7943]) );
  DFF ram_reg_1055__6_ ( .D(n12183), .CP(wclk), .Q(ram[7942]) );
  DFF ram_reg_1055__5_ ( .D(n12182), .CP(wclk), .Q(ram[7941]) );
  DFF ram_reg_1055__4_ ( .D(n12181), .CP(wclk), .Q(ram[7940]) );
  DFF ram_reg_1055__3_ ( .D(n12180), .CP(wclk), .Q(ram[7939]) );
  DFF ram_reg_1055__2_ ( .D(n12179), .CP(wclk), .Q(ram[7938]) );
  DFF ram_reg_1055__1_ ( .D(n12178), .CP(wclk), .Q(ram[7937]) );
  DFF ram_reg_1055__0_ ( .D(n12177), .CP(wclk), .Q(ram[7936]) );
  DFF ram_reg_1063__7_ ( .D(n12120), .CP(wclk), .Q(ram[7879]) );
  DFF ram_reg_1063__6_ ( .D(n12119), .CP(wclk), .Q(ram[7878]) );
  DFF ram_reg_1063__5_ ( .D(n12118), .CP(wclk), .Q(ram[7877]) );
  DFF ram_reg_1063__4_ ( .D(n12117), .CP(wclk), .Q(ram[7876]) );
  DFF ram_reg_1063__3_ ( .D(n12116), .CP(wclk), .Q(ram[7875]) );
  DFF ram_reg_1063__2_ ( .D(n12115), .CP(wclk), .Q(ram[7874]) );
  DFF ram_reg_1063__1_ ( .D(n12114), .CP(wclk), .Q(ram[7873]) );
  DFF ram_reg_1063__0_ ( .D(n12113), .CP(wclk), .Q(ram[7872]) );
  DFF ram_reg_1079__7_ ( .D(n11992), .CP(wclk), .Q(ram[7751]) );
  DFF ram_reg_1079__6_ ( .D(n11991), .CP(wclk), .Q(ram[7750]) );
  DFF ram_reg_1079__5_ ( .D(n11990), .CP(wclk), .Q(ram[7749]) );
  DFF ram_reg_1079__4_ ( .D(n11989), .CP(wclk), .Q(ram[7748]) );
  DFF ram_reg_1079__3_ ( .D(n11988), .CP(wclk), .Q(ram[7747]) );
  DFF ram_reg_1079__2_ ( .D(n11987), .CP(wclk), .Q(ram[7746]) );
  DFF ram_reg_1079__1_ ( .D(n11986), .CP(wclk), .Q(ram[7745]) );
  DFF ram_reg_1079__0_ ( .D(n11985), .CP(wclk), .Q(ram[7744]) );
  DFF ram_reg_1091__7_ ( .D(n11896), .CP(wclk), .Q(ram[7655]) );
  DFF ram_reg_1091__6_ ( .D(n11895), .CP(wclk), .Q(ram[7654]) );
  DFF ram_reg_1091__5_ ( .D(n11894), .CP(wclk), .Q(ram[7653]) );
  DFF ram_reg_1091__4_ ( .D(n11893), .CP(wclk), .Q(ram[7652]) );
  DFF ram_reg_1091__3_ ( .D(n11892), .CP(wclk), .Q(ram[7651]) );
  DFF ram_reg_1091__2_ ( .D(n11891), .CP(wclk), .Q(ram[7650]) );
  DFF ram_reg_1091__1_ ( .D(n11890), .CP(wclk), .Q(ram[7649]) );
  DFF ram_reg_1091__0_ ( .D(n11889), .CP(wclk), .Q(ram[7648]) );
  DFF ram_reg_1095__7_ ( .D(n11864), .CP(wclk), .Q(ram[7623]) );
  DFF ram_reg_1095__6_ ( .D(n11863), .CP(wclk), .Q(ram[7622]) );
  DFF ram_reg_1095__5_ ( .D(n11862), .CP(wclk), .Q(ram[7621]) );
  DFF ram_reg_1095__4_ ( .D(n11861), .CP(wclk), .Q(ram[7620]) );
  DFF ram_reg_1095__3_ ( .D(n11860), .CP(wclk), .Q(ram[7619]) );
  DFF ram_reg_1095__2_ ( .D(n11859), .CP(wclk), .Q(ram[7618]) );
  DFF ram_reg_1095__1_ ( .D(n11858), .CP(wclk), .Q(ram[7617]) );
  DFF ram_reg_1095__0_ ( .D(n11857), .CP(wclk), .Q(ram[7616]) );
  DFF ram_reg_1099__7_ ( .D(n11832), .CP(wclk), .Q(ram[7591]) );
  DFF ram_reg_1099__6_ ( .D(n11831), .CP(wclk), .Q(ram[7590]) );
  DFF ram_reg_1099__5_ ( .D(n11830), .CP(wclk), .Q(ram[7589]) );
  DFF ram_reg_1099__4_ ( .D(n11829), .CP(wclk), .Q(ram[7588]) );
  DFF ram_reg_1099__3_ ( .D(n11828), .CP(wclk), .Q(ram[7587]) );
  DFF ram_reg_1099__2_ ( .D(n11827), .CP(wclk), .Q(ram[7586]) );
  DFF ram_reg_1099__1_ ( .D(n11826), .CP(wclk), .Q(ram[7585]) );
  DFF ram_reg_1099__0_ ( .D(n11825), .CP(wclk), .Q(ram[7584]) );
  DFF ram_reg_1103__7_ ( .D(n11800), .CP(wclk), .Q(ram[7559]) );
  DFF ram_reg_1103__6_ ( .D(n11799), .CP(wclk), .Q(ram[7558]) );
  DFF ram_reg_1103__5_ ( .D(n11798), .CP(wclk), .Q(ram[7557]) );
  DFF ram_reg_1103__4_ ( .D(n11797), .CP(wclk), .Q(ram[7556]) );
  DFF ram_reg_1103__3_ ( .D(n11796), .CP(wclk), .Q(ram[7555]) );
  DFF ram_reg_1103__2_ ( .D(n11795), .CP(wclk), .Q(ram[7554]) );
  DFF ram_reg_1103__1_ ( .D(n11794), .CP(wclk), .Q(ram[7553]) );
  DFF ram_reg_1103__0_ ( .D(n11793), .CP(wclk), .Q(ram[7552]) );
  DFF ram_reg_1107__7_ ( .D(n11768), .CP(wclk), .Q(ram[7527]) );
  DFF ram_reg_1107__6_ ( .D(n11767), .CP(wclk), .Q(ram[7526]) );
  DFF ram_reg_1107__5_ ( .D(n11766), .CP(wclk), .Q(ram[7525]) );
  DFF ram_reg_1107__4_ ( .D(n11765), .CP(wclk), .Q(ram[7524]) );
  DFF ram_reg_1107__3_ ( .D(n11764), .CP(wclk), .Q(ram[7523]) );
  DFF ram_reg_1107__2_ ( .D(n11763), .CP(wclk), .Q(ram[7522]) );
  DFF ram_reg_1107__1_ ( .D(n11762), .CP(wclk), .Q(ram[7521]) );
  DFF ram_reg_1107__0_ ( .D(n11761), .CP(wclk), .Q(ram[7520]) );
  DFF ram_reg_1111__7_ ( .D(n11736), .CP(wclk), .Q(ram[7495]) );
  DFF ram_reg_1111__6_ ( .D(n11735), .CP(wclk), .Q(ram[7494]) );
  DFF ram_reg_1111__5_ ( .D(n11734), .CP(wclk), .Q(ram[7493]) );
  DFF ram_reg_1111__4_ ( .D(n11733), .CP(wclk), .Q(ram[7492]) );
  DFF ram_reg_1111__3_ ( .D(n11732), .CP(wclk), .Q(ram[7491]) );
  DFF ram_reg_1111__2_ ( .D(n11731), .CP(wclk), .Q(ram[7490]) );
  DFF ram_reg_1111__1_ ( .D(n11730), .CP(wclk), .Q(ram[7489]) );
  DFF ram_reg_1111__0_ ( .D(n11729), .CP(wclk), .Q(ram[7488]) );
  DFF ram_reg_1115__7_ ( .D(n11704), .CP(wclk), .Q(ram[7463]) );
  DFF ram_reg_1115__6_ ( .D(n11703), .CP(wclk), .Q(ram[7462]) );
  DFF ram_reg_1115__5_ ( .D(n11702), .CP(wclk), .Q(ram[7461]) );
  DFF ram_reg_1115__4_ ( .D(n11701), .CP(wclk), .Q(ram[7460]) );
  DFF ram_reg_1115__3_ ( .D(n11700), .CP(wclk), .Q(ram[7459]) );
  DFF ram_reg_1115__2_ ( .D(n11699), .CP(wclk), .Q(ram[7458]) );
  DFF ram_reg_1115__1_ ( .D(n11698), .CP(wclk), .Q(ram[7457]) );
  DFF ram_reg_1115__0_ ( .D(n11697), .CP(wclk), .Q(ram[7456]) );
  DFF ram_reg_1119__7_ ( .D(n11672), .CP(wclk), .Q(ram[7431]) );
  DFF ram_reg_1119__6_ ( .D(n11671), .CP(wclk), .Q(ram[7430]) );
  DFF ram_reg_1119__5_ ( .D(n11670), .CP(wclk), .Q(ram[7429]) );
  DFF ram_reg_1119__4_ ( .D(n11669), .CP(wclk), .Q(ram[7428]) );
  DFF ram_reg_1119__3_ ( .D(n11668), .CP(wclk), .Q(ram[7427]) );
  DFF ram_reg_1119__2_ ( .D(n11667), .CP(wclk), .Q(ram[7426]) );
  DFF ram_reg_1119__1_ ( .D(n11666), .CP(wclk), .Q(ram[7425]) );
  DFF ram_reg_1119__0_ ( .D(n11665), .CP(wclk), .Q(ram[7424]) );
  DFF ram_reg_1123__7_ ( .D(n11640), .CP(wclk), .Q(ram[7399]) );
  DFF ram_reg_1123__6_ ( .D(n11639), .CP(wclk), .Q(ram[7398]) );
  DFF ram_reg_1123__5_ ( .D(n11638), .CP(wclk), .Q(ram[7397]) );
  DFF ram_reg_1123__4_ ( .D(n11637), .CP(wclk), .Q(ram[7396]) );
  DFF ram_reg_1123__3_ ( .D(n11636), .CP(wclk), .Q(ram[7395]) );
  DFF ram_reg_1123__2_ ( .D(n11635), .CP(wclk), .Q(ram[7394]) );
  DFF ram_reg_1123__1_ ( .D(n11634), .CP(wclk), .Q(ram[7393]) );
  DFF ram_reg_1123__0_ ( .D(n11633), .CP(wclk), .Q(ram[7392]) );
  DFF ram_reg_1127__7_ ( .D(n11608), .CP(wclk), .Q(ram[7367]) );
  DFF ram_reg_1127__6_ ( .D(n11607), .CP(wclk), .Q(ram[7366]) );
  DFF ram_reg_1127__5_ ( .D(n11606), .CP(wclk), .Q(ram[7365]) );
  DFF ram_reg_1127__4_ ( .D(n11605), .CP(wclk), .Q(ram[7364]) );
  DFF ram_reg_1127__3_ ( .D(n11604), .CP(wclk), .Q(ram[7363]) );
  DFF ram_reg_1127__2_ ( .D(n11603), .CP(wclk), .Q(ram[7362]) );
  DFF ram_reg_1127__1_ ( .D(n11602), .CP(wclk), .Q(ram[7361]) );
  DFF ram_reg_1127__0_ ( .D(n11601), .CP(wclk), .Q(ram[7360]) );
  DFF ram_reg_1135__7_ ( .D(n11544), .CP(wclk), .Q(ram[7303]) );
  DFF ram_reg_1135__6_ ( .D(n11543), .CP(wclk), .Q(ram[7302]) );
  DFF ram_reg_1135__5_ ( .D(n11542), .CP(wclk), .Q(ram[7301]) );
  DFF ram_reg_1135__4_ ( .D(n11541), .CP(wclk), .Q(ram[7300]) );
  DFF ram_reg_1135__3_ ( .D(n11540), .CP(wclk), .Q(ram[7299]) );
  DFF ram_reg_1135__2_ ( .D(n11539), .CP(wclk), .Q(ram[7298]) );
  DFF ram_reg_1135__1_ ( .D(n11538), .CP(wclk), .Q(ram[7297]) );
  DFF ram_reg_1135__0_ ( .D(n11537), .CP(wclk), .Q(ram[7296]) );
  DFF ram_reg_1139__7_ ( .D(n11512), .CP(wclk), .Q(ram[7271]) );
  DFF ram_reg_1139__6_ ( .D(n11511), .CP(wclk), .Q(ram[7270]) );
  DFF ram_reg_1139__5_ ( .D(n11510), .CP(wclk), .Q(ram[7269]) );
  DFF ram_reg_1139__4_ ( .D(n11509), .CP(wclk), .Q(ram[7268]) );
  DFF ram_reg_1139__3_ ( .D(n11508), .CP(wclk), .Q(ram[7267]) );
  DFF ram_reg_1139__2_ ( .D(n11507), .CP(wclk), .Q(ram[7266]) );
  DFF ram_reg_1139__1_ ( .D(n11506), .CP(wclk), .Q(ram[7265]) );
  DFF ram_reg_1139__0_ ( .D(n11505), .CP(wclk), .Q(ram[7264]) );
  DFF ram_reg_1143__7_ ( .D(n11480), .CP(wclk), .Q(ram[7239]) );
  DFF ram_reg_1143__6_ ( .D(n11479), .CP(wclk), .Q(ram[7238]) );
  DFF ram_reg_1143__5_ ( .D(n11478), .CP(wclk), .Q(ram[7237]) );
  DFF ram_reg_1143__4_ ( .D(n11477), .CP(wclk), .Q(ram[7236]) );
  DFF ram_reg_1143__3_ ( .D(n11476), .CP(wclk), .Q(ram[7235]) );
  DFF ram_reg_1143__2_ ( .D(n11475), .CP(wclk), .Q(ram[7234]) );
  DFF ram_reg_1143__1_ ( .D(n11474), .CP(wclk), .Q(ram[7233]) );
  DFF ram_reg_1143__0_ ( .D(n11473), .CP(wclk), .Q(ram[7232]) );
  DFF ram_reg_1159__7_ ( .D(n11352), .CP(wclk), .Q(ram[7111]) );
  DFF ram_reg_1159__6_ ( .D(n11351), .CP(wclk), .Q(ram[7110]) );
  DFF ram_reg_1159__5_ ( .D(n11350), .CP(wclk), .Q(ram[7109]) );
  DFF ram_reg_1159__4_ ( .D(n11349), .CP(wclk), .Q(ram[7108]) );
  DFF ram_reg_1159__3_ ( .D(n11348), .CP(wclk), .Q(ram[7107]) );
  DFF ram_reg_1159__2_ ( .D(n11347), .CP(wclk), .Q(ram[7106]) );
  DFF ram_reg_1159__1_ ( .D(n11346), .CP(wclk), .Q(ram[7105]) );
  DFF ram_reg_1159__0_ ( .D(n11345), .CP(wclk), .Q(ram[7104]) );
  DFF ram_reg_1175__7_ ( .D(n11224), .CP(wclk), .Q(ram[6983]) );
  DFF ram_reg_1175__6_ ( .D(n11223), .CP(wclk), .Q(ram[6982]) );
  DFF ram_reg_1175__5_ ( .D(n11222), .CP(wclk), .Q(ram[6981]) );
  DFF ram_reg_1175__4_ ( .D(n11221), .CP(wclk), .Q(ram[6980]) );
  DFF ram_reg_1175__3_ ( .D(n11220), .CP(wclk), .Q(ram[6979]) );
  DFF ram_reg_1175__2_ ( .D(n11219), .CP(wclk), .Q(ram[6978]) );
  DFF ram_reg_1175__1_ ( .D(n11218), .CP(wclk), .Q(ram[6977]) );
  DFF ram_reg_1175__0_ ( .D(n11217), .CP(wclk), .Q(ram[6976]) );
  DFF ram_reg_1223__7_ ( .D(n10840), .CP(wclk), .Q(ram[6599]) );
  DFF ram_reg_1223__6_ ( .D(n10839), .CP(wclk), .Q(ram[6598]) );
  DFF ram_reg_1223__5_ ( .D(n10838), .CP(wclk), .Q(ram[6597]) );
  DFF ram_reg_1223__4_ ( .D(n10837), .CP(wclk), .Q(ram[6596]) );
  DFF ram_reg_1223__3_ ( .D(n10836), .CP(wclk), .Q(ram[6595]) );
  DFF ram_reg_1223__2_ ( .D(n10835), .CP(wclk), .Q(ram[6594]) );
  DFF ram_reg_1223__1_ ( .D(n10834), .CP(wclk), .Q(ram[6593]) );
  DFF ram_reg_1223__0_ ( .D(n10833), .CP(wclk), .Q(ram[6592]) );
  DFF ram_reg_1235__7_ ( .D(n10744), .CP(wclk), .Q(ram[6503]) );
  DFF ram_reg_1235__6_ ( .D(n10743), .CP(wclk), .Q(ram[6502]) );
  DFF ram_reg_1235__5_ ( .D(n10742), .CP(wclk), .Q(ram[6501]) );
  DFF ram_reg_1235__4_ ( .D(n10741), .CP(wclk), .Q(ram[6500]) );
  DFF ram_reg_1235__3_ ( .D(n10740), .CP(wclk), .Q(ram[6499]) );
  DFF ram_reg_1235__2_ ( .D(n10739), .CP(wclk), .Q(ram[6498]) );
  DFF ram_reg_1235__1_ ( .D(n10738), .CP(wclk), .Q(ram[6497]) );
  DFF ram_reg_1235__0_ ( .D(n10737), .CP(wclk), .Q(ram[6496]) );
  DFF ram_reg_1239__7_ ( .D(n10712), .CP(wclk), .Q(ram[6471]) );
  DFF ram_reg_1239__6_ ( .D(n10711), .CP(wclk), .Q(ram[6470]) );
  DFF ram_reg_1239__5_ ( .D(n10710), .CP(wclk), .Q(ram[6469]) );
  DFF ram_reg_1239__4_ ( .D(n10709), .CP(wclk), .Q(ram[6468]) );
  DFF ram_reg_1239__3_ ( .D(n10708), .CP(wclk), .Q(ram[6467]) );
  DFF ram_reg_1239__2_ ( .D(n10707), .CP(wclk), .Q(ram[6466]) );
  DFF ram_reg_1239__1_ ( .D(n10706), .CP(wclk), .Q(ram[6465]) );
  DFF ram_reg_1239__0_ ( .D(n10705), .CP(wclk), .Q(ram[6464]) );
  DFF ram_reg_1255__7_ ( .D(n10584), .CP(wclk), .Q(ram[6343]) );
  DFF ram_reg_1255__6_ ( .D(n10583), .CP(wclk), .Q(ram[6342]) );
  DFF ram_reg_1255__5_ ( .D(n10582), .CP(wclk), .Q(ram[6341]) );
  DFF ram_reg_1255__4_ ( .D(n10581), .CP(wclk), .Q(ram[6340]) );
  DFF ram_reg_1255__3_ ( .D(n10580), .CP(wclk), .Q(ram[6339]) );
  DFF ram_reg_1255__2_ ( .D(n10579), .CP(wclk), .Q(ram[6338]) );
  DFF ram_reg_1255__1_ ( .D(n10578), .CP(wclk), .Q(ram[6337]) );
  DFF ram_reg_1255__0_ ( .D(n10577), .CP(wclk), .Q(ram[6336]) );
  DFF ram_reg_1287__7_ ( .D(n10328), .CP(wclk), .Q(ram[6087]) );
  DFF ram_reg_1287__6_ ( .D(n10327), .CP(wclk), .Q(ram[6086]) );
  DFF ram_reg_1287__5_ ( .D(n10326), .CP(wclk), .Q(ram[6085]) );
  DFF ram_reg_1287__4_ ( .D(n10325), .CP(wclk), .Q(ram[6084]) );
  DFF ram_reg_1287__3_ ( .D(n10324), .CP(wclk), .Q(ram[6083]) );
  DFF ram_reg_1287__2_ ( .D(n10323), .CP(wclk), .Q(ram[6082]) );
  DFF ram_reg_1287__1_ ( .D(n10322), .CP(wclk), .Q(ram[6081]) );
  DFF ram_reg_1287__0_ ( .D(n10321), .CP(wclk), .Q(ram[6080]) );
  DFF ram_reg_1303__7_ ( .D(n10200), .CP(wclk), .Q(ram[5959]) );
  DFF ram_reg_1303__6_ ( .D(n10199), .CP(wclk), .Q(ram[5958]) );
  DFF ram_reg_1303__5_ ( .D(n10198), .CP(wclk), .Q(ram[5957]) );
  DFF ram_reg_1303__4_ ( .D(n10197), .CP(wclk), .Q(ram[5956]) );
  DFF ram_reg_1303__3_ ( .D(n10196), .CP(wclk), .Q(ram[5955]) );
  DFF ram_reg_1303__2_ ( .D(n10195), .CP(wclk), .Q(ram[5954]) );
  DFF ram_reg_1303__1_ ( .D(n10194), .CP(wclk), .Q(ram[5953]) );
  DFF ram_reg_1303__0_ ( .D(n10193), .CP(wclk), .Q(ram[5952]) );
  DFF ram_reg_1319__7_ ( .D(n10072), .CP(wclk), .Q(ram[5831]) );
  DFF ram_reg_1319__6_ ( .D(n10071), .CP(wclk), .Q(ram[5830]) );
  DFF ram_reg_1319__5_ ( .D(n10070), .CP(wclk), .Q(ram[5829]) );
  DFF ram_reg_1319__4_ ( .D(n10069), .CP(wclk), .Q(ram[5828]) );
  DFF ram_reg_1319__3_ ( .D(n10068), .CP(wclk), .Q(ram[5827]) );
  DFF ram_reg_1319__2_ ( .D(n10067), .CP(wclk), .Q(ram[5826]) );
  DFF ram_reg_1319__1_ ( .D(n10066), .CP(wclk), .Q(ram[5825]) );
  DFF ram_reg_1319__0_ ( .D(n10065), .CP(wclk), .Q(ram[5824]) );
  DFF ram_reg_1347__7_ ( .D(n9848), .CP(wclk), .Q(ram[5607]) );
  DFF ram_reg_1347__6_ ( .D(n9847), .CP(wclk), .Q(ram[5606]) );
  DFF ram_reg_1347__5_ ( .D(n9846), .CP(wclk), .Q(ram[5605]) );
  DFF ram_reg_1347__4_ ( .D(n9845), .CP(wclk), .Q(ram[5604]) );
  DFF ram_reg_1347__3_ ( .D(n9844), .CP(wclk), .Q(ram[5603]) );
  DFF ram_reg_1347__2_ ( .D(n9843), .CP(wclk), .Q(ram[5602]) );
  DFF ram_reg_1347__1_ ( .D(n9842), .CP(wclk), .Q(ram[5601]) );
  DFF ram_reg_1347__0_ ( .D(n9841), .CP(wclk), .Q(ram[5600]) );
  DFF ram_reg_1351__7_ ( .D(n9816), .CP(wclk), .Q(ram[5575]) );
  DFF ram_reg_1351__6_ ( .D(n9815), .CP(wclk), .Q(ram[5574]) );
  DFF ram_reg_1351__5_ ( .D(n9814), .CP(wclk), .Q(ram[5573]) );
  DFF ram_reg_1351__4_ ( .D(n9813), .CP(wclk), .Q(ram[5572]) );
  DFF ram_reg_1351__3_ ( .D(n9812), .CP(wclk), .Q(ram[5571]) );
  DFF ram_reg_1351__2_ ( .D(n9811), .CP(wclk), .Q(ram[5570]) );
  DFF ram_reg_1351__1_ ( .D(n9810), .CP(wclk), .Q(ram[5569]) );
  DFF ram_reg_1351__0_ ( .D(n9809), .CP(wclk), .Q(ram[5568]) );
  DFF ram_reg_1363__7_ ( .D(n9720), .CP(wclk), .Q(ram[5479]) );
  DFF ram_reg_1363__6_ ( .D(n9719), .CP(wclk), .Q(ram[5478]) );
  DFF ram_reg_1363__5_ ( .D(n9718), .CP(wclk), .Q(ram[5477]) );
  DFF ram_reg_1363__4_ ( .D(n9717), .CP(wclk), .Q(ram[5476]) );
  DFF ram_reg_1363__3_ ( .D(n9716), .CP(wclk), .Q(ram[5475]) );
  DFF ram_reg_1363__2_ ( .D(n9715), .CP(wclk), .Q(ram[5474]) );
  DFF ram_reg_1363__1_ ( .D(n9714), .CP(wclk), .Q(ram[5473]) );
  DFF ram_reg_1363__0_ ( .D(n9713), .CP(wclk), .Q(ram[5472]) );
  DFF ram_reg_1367__7_ ( .D(n9688), .CP(wclk), .Q(ram[5447]) );
  DFF ram_reg_1367__6_ ( .D(n9687), .CP(wclk), .Q(ram[5446]) );
  DFF ram_reg_1367__5_ ( .D(n9686), .CP(wclk), .Q(ram[5445]) );
  DFF ram_reg_1367__4_ ( .D(n9685), .CP(wclk), .Q(ram[5444]) );
  DFF ram_reg_1367__3_ ( .D(n9684), .CP(wclk), .Q(ram[5443]) );
  DFF ram_reg_1367__2_ ( .D(n9683), .CP(wclk), .Q(ram[5442]) );
  DFF ram_reg_1367__1_ ( .D(n9682), .CP(wclk), .Q(ram[5441]) );
  DFF ram_reg_1367__0_ ( .D(n9681), .CP(wclk), .Q(ram[5440]) );
  DFF ram_reg_1375__7_ ( .D(n9624), .CP(wclk), .Q(ram[5383]) );
  DFF ram_reg_1375__6_ ( .D(n9623), .CP(wclk), .Q(ram[5382]) );
  DFF ram_reg_1375__5_ ( .D(n9622), .CP(wclk), .Q(ram[5381]) );
  DFF ram_reg_1375__4_ ( .D(n9621), .CP(wclk), .Q(ram[5380]) );
  DFF ram_reg_1375__3_ ( .D(n9620), .CP(wclk), .Q(ram[5379]) );
  DFF ram_reg_1375__2_ ( .D(n9619), .CP(wclk), .Q(ram[5378]) );
  DFF ram_reg_1375__1_ ( .D(n9618), .CP(wclk), .Q(ram[5377]) );
  DFF ram_reg_1375__0_ ( .D(n9617), .CP(wclk), .Q(ram[5376]) );
  DFF ram_reg_1379__7_ ( .D(n9592), .CP(wclk), .Q(ram[5351]) );
  DFF ram_reg_1379__6_ ( .D(n9591), .CP(wclk), .Q(ram[5350]) );
  DFF ram_reg_1379__5_ ( .D(n9590), .CP(wclk), .Q(ram[5349]) );
  DFF ram_reg_1379__4_ ( .D(n9589), .CP(wclk), .Q(ram[5348]) );
  DFF ram_reg_1379__3_ ( .D(n9588), .CP(wclk), .Q(ram[5347]) );
  DFF ram_reg_1379__2_ ( .D(n9587), .CP(wclk), .Q(ram[5346]) );
  DFF ram_reg_1379__1_ ( .D(n9586), .CP(wclk), .Q(ram[5345]) );
  DFF ram_reg_1379__0_ ( .D(n9585), .CP(wclk), .Q(ram[5344]) );
  DFF ram_reg_1383__7_ ( .D(n9560), .CP(wclk), .Q(ram[5319]) );
  DFF ram_reg_1383__6_ ( .D(n9559), .CP(wclk), .Q(ram[5318]) );
  DFF ram_reg_1383__5_ ( .D(n9558), .CP(wclk), .Q(ram[5317]) );
  DFF ram_reg_1383__4_ ( .D(n9557), .CP(wclk), .Q(ram[5316]) );
  DFF ram_reg_1383__3_ ( .D(n9556), .CP(wclk), .Q(ram[5315]) );
  DFF ram_reg_1383__2_ ( .D(n9555), .CP(wclk), .Q(ram[5314]) );
  DFF ram_reg_1383__1_ ( .D(n9554), .CP(wclk), .Q(ram[5313]) );
  DFF ram_reg_1383__0_ ( .D(n9553), .CP(wclk), .Q(ram[5312]) );
  DFF ram_reg_1399__7_ ( .D(n9432), .CP(wclk), .Q(ram[5191]) );
  DFF ram_reg_1399__6_ ( .D(n9431), .CP(wclk), .Q(ram[5190]) );
  DFF ram_reg_1399__5_ ( .D(n9430), .CP(wclk), .Q(ram[5189]) );
  DFF ram_reg_1399__4_ ( .D(n9429), .CP(wclk), .Q(ram[5188]) );
  DFF ram_reg_1399__3_ ( .D(n9428), .CP(wclk), .Q(ram[5187]) );
  DFF ram_reg_1399__2_ ( .D(n9427), .CP(wclk), .Q(ram[5186]) );
  DFF ram_reg_1399__1_ ( .D(n9426), .CP(wclk), .Q(ram[5185]) );
  DFF ram_reg_1399__0_ ( .D(n9425), .CP(wclk), .Q(ram[5184]) );
  DFF ram_reg_1495__7_ ( .D(n8664), .CP(wclk), .Q(ram[4423]) );
  DFF ram_reg_1495__6_ ( .D(n8663), .CP(wclk), .Q(ram[4422]) );
  DFF ram_reg_1495__5_ ( .D(n8662), .CP(wclk), .Q(ram[4421]) );
  DFF ram_reg_1495__4_ ( .D(n8661), .CP(wclk), .Q(ram[4420]) );
  DFF ram_reg_1495__3_ ( .D(n8660), .CP(wclk), .Q(ram[4419]) );
  DFF ram_reg_1495__2_ ( .D(n8659), .CP(wclk), .Q(ram[4418]) );
  DFF ram_reg_1495__1_ ( .D(n8658), .CP(wclk), .Q(ram[4417]) );
  DFF ram_reg_1495__0_ ( .D(n8657), .CP(wclk), .Q(ram[4416]) );
  DFF ram_reg_1539__7_ ( .D(n8312), .CP(wclk), .Q(ram[4071]) );
  DFF ram_reg_1539__6_ ( .D(n8311), .CP(wclk), .Q(ram[4070]) );
  DFF ram_reg_1539__5_ ( .D(n8310), .CP(wclk), .Q(ram[4069]) );
  DFF ram_reg_1539__4_ ( .D(n8309), .CP(wclk), .Q(ram[4068]) );
  DFF ram_reg_1539__3_ ( .D(n8308), .CP(wclk), .Q(ram[4067]) );
  DFF ram_reg_1539__2_ ( .D(n8307), .CP(wclk), .Q(ram[4066]) );
  DFF ram_reg_1539__1_ ( .D(n8306), .CP(wclk), .Q(ram[4065]) );
  DFF ram_reg_1539__0_ ( .D(n8305), .CP(wclk), .Q(ram[4064]) );
  DFF ram_reg_1543__7_ ( .D(n8280), .CP(wclk), .Q(ram[4039]) );
  DFF ram_reg_1543__6_ ( .D(n8279), .CP(wclk), .Q(ram[4038]) );
  DFF ram_reg_1543__5_ ( .D(n8278), .CP(wclk), .Q(ram[4037]) );
  DFF ram_reg_1543__4_ ( .D(n8277), .CP(wclk), .Q(ram[4036]) );
  DFF ram_reg_1543__3_ ( .D(n8276), .CP(wclk), .Q(ram[4035]) );
  DFF ram_reg_1543__2_ ( .D(n8275), .CP(wclk), .Q(ram[4034]) );
  DFF ram_reg_1543__1_ ( .D(n8274), .CP(wclk), .Q(ram[4033]) );
  DFF ram_reg_1543__0_ ( .D(n8273), .CP(wclk), .Q(ram[4032]) );
  DFF ram_reg_1555__7_ ( .D(n8184), .CP(wclk), .Q(ram[3943]) );
  DFF ram_reg_1555__6_ ( .D(n8183), .CP(wclk), .Q(ram[3942]) );
  DFF ram_reg_1555__5_ ( .D(n8182), .CP(wclk), .Q(ram[3941]) );
  DFF ram_reg_1555__4_ ( .D(n8181), .CP(wclk), .Q(ram[3940]) );
  DFF ram_reg_1555__3_ ( .D(n8180), .CP(wclk), .Q(ram[3939]) );
  DFF ram_reg_1555__2_ ( .D(n8179), .CP(wclk), .Q(ram[3938]) );
  DFF ram_reg_1555__1_ ( .D(n8178), .CP(wclk), .Q(ram[3937]) );
  DFF ram_reg_1555__0_ ( .D(n8177), .CP(wclk), .Q(ram[3936]) );
  DFF ram_reg_1559__7_ ( .D(n8152), .CP(wclk), .Q(ram[3911]) );
  DFF ram_reg_1559__6_ ( .D(n8151), .CP(wclk), .Q(ram[3910]) );
  DFF ram_reg_1559__5_ ( .D(n8150), .CP(wclk), .Q(ram[3909]) );
  DFF ram_reg_1559__4_ ( .D(n8149), .CP(wclk), .Q(ram[3908]) );
  DFF ram_reg_1559__3_ ( .D(n8148), .CP(wclk), .Q(ram[3907]) );
  DFF ram_reg_1559__2_ ( .D(n8147), .CP(wclk), .Q(ram[3906]) );
  DFF ram_reg_1559__1_ ( .D(n8146), .CP(wclk), .Q(ram[3905]) );
  DFF ram_reg_1559__0_ ( .D(n8145), .CP(wclk), .Q(ram[3904]) );
  DFF ram_reg_1567__7_ ( .D(n8088), .CP(wclk), .Q(ram[3847]) );
  DFF ram_reg_1567__6_ ( .D(n8087), .CP(wclk), .Q(ram[3846]) );
  DFF ram_reg_1567__5_ ( .D(n8086), .CP(wclk), .Q(ram[3845]) );
  DFF ram_reg_1567__4_ ( .D(n8085), .CP(wclk), .Q(ram[3844]) );
  DFF ram_reg_1567__3_ ( .D(n8084), .CP(wclk), .Q(ram[3843]) );
  DFF ram_reg_1567__2_ ( .D(n8083), .CP(wclk), .Q(ram[3842]) );
  DFF ram_reg_1567__1_ ( .D(n8082), .CP(wclk), .Q(ram[3841]) );
  DFF ram_reg_1567__0_ ( .D(n8081), .CP(wclk), .Q(ram[3840]) );
  DFF ram_reg_1575__7_ ( .D(n8024), .CP(wclk), .Q(ram[3783]) );
  DFF ram_reg_1575__6_ ( .D(n8023), .CP(wclk), .Q(ram[3782]) );
  DFF ram_reg_1575__5_ ( .D(n8022), .CP(wclk), .Q(ram[3781]) );
  DFF ram_reg_1575__4_ ( .D(n8021), .CP(wclk), .Q(ram[3780]) );
  DFF ram_reg_1575__3_ ( .D(n8020), .CP(wclk), .Q(ram[3779]) );
  DFF ram_reg_1575__2_ ( .D(n8019), .CP(wclk), .Q(ram[3778]) );
  DFF ram_reg_1575__1_ ( .D(n8018), .CP(wclk), .Q(ram[3777]) );
  DFF ram_reg_1575__0_ ( .D(n8017), .CP(wclk), .Q(ram[3776]) );
  DFF ram_reg_1591__7_ ( .D(n7896), .CP(wclk), .Q(ram[3655]) );
  DFF ram_reg_1591__6_ ( .D(n7895), .CP(wclk), .Q(ram[3654]) );
  DFF ram_reg_1591__5_ ( .D(n7894), .CP(wclk), .Q(ram[3653]) );
  DFF ram_reg_1591__4_ ( .D(n7893), .CP(wclk), .Q(ram[3652]) );
  DFF ram_reg_1591__3_ ( .D(n7892), .CP(wclk), .Q(ram[3651]) );
  DFF ram_reg_1591__2_ ( .D(n7891), .CP(wclk), .Q(ram[3650]) );
  DFF ram_reg_1591__1_ ( .D(n7890), .CP(wclk), .Q(ram[3649]) );
  DFF ram_reg_1591__0_ ( .D(n7889), .CP(wclk), .Q(ram[3648]) );
  DFF ram_reg_1603__7_ ( .D(n7800), .CP(wclk), .Q(ram[3559]) );
  DFF ram_reg_1603__6_ ( .D(n7799), .CP(wclk), .Q(ram[3558]) );
  DFF ram_reg_1603__5_ ( .D(n7798), .CP(wclk), .Q(ram[3557]) );
  DFF ram_reg_1603__4_ ( .D(n7797), .CP(wclk), .Q(ram[3556]) );
  DFF ram_reg_1603__3_ ( .D(n7796), .CP(wclk), .Q(ram[3555]) );
  DFF ram_reg_1603__2_ ( .D(n7795), .CP(wclk), .Q(ram[3554]) );
  DFF ram_reg_1603__1_ ( .D(n7794), .CP(wclk), .Q(ram[3553]) );
  DFF ram_reg_1603__0_ ( .D(n7793), .CP(wclk), .Q(ram[3552]) );
  DFF ram_reg_1607__7_ ( .D(n7768), .CP(wclk), .Q(ram[3527]) );
  DFF ram_reg_1607__6_ ( .D(n7767), .CP(wclk), .Q(ram[3526]) );
  DFF ram_reg_1607__5_ ( .D(n7766), .CP(wclk), .Q(ram[3525]) );
  DFF ram_reg_1607__4_ ( .D(n7765), .CP(wclk), .Q(ram[3524]) );
  DFF ram_reg_1607__3_ ( .D(n7764), .CP(wclk), .Q(ram[3523]) );
  DFF ram_reg_1607__2_ ( .D(n7763), .CP(wclk), .Q(ram[3522]) );
  DFF ram_reg_1607__1_ ( .D(n7762), .CP(wclk), .Q(ram[3521]) );
  DFF ram_reg_1607__0_ ( .D(n7761), .CP(wclk), .Q(ram[3520]) );
  DFF ram_reg_1611__7_ ( .D(n7736), .CP(wclk), .Q(ram[3495]) );
  DFF ram_reg_1611__6_ ( .D(n7735), .CP(wclk), .Q(ram[3494]) );
  DFF ram_reg_1611__5_ ( .D(n7734), .CP(wclk), .Q(ram[3493]) );
  DFF ram_reg_1611__4_ ( .D(n7733), .CP(wclk), .Q(ram[3492]) );
  DFF ram_reg_1611__3_ ( .D(n7732), .CP(wclk), .Q(ram[3491]) );
  DFF ram_reg_1611__2_ ( .D(n7731), .CP(wclk), .Q(ram[3490]) );
  DFF ram_reg_1611__1_ ( .D(n7730), .CP(wclk), .Q(ram[3489]) );
  DFF ram_reg_1611__0_ ( .D(n7729), .CP(wclk), .Q(ram[3488]) );
  DFF ram_reg_1615__7_ ( .D(n7704), .CP(wclk), .Q(ram[3463]) );
  DFF ram_reg_1615__6_ ( .D(n7703), .CP(wclk), .Q(ram[3462]) );
  DFF ram_reg_1615__5_ ( .D(n7702), .CP(wclk), .Q(ram[3461]) );
  DFF ram_reg_1615__4_ ( .D(n7701), .CP(wclk), .Q(ram[3460]) );
  DFF ram_reg_1615__3_ ( .D(n7700), .CP(wclk), .Q(ram[3459]) );
  DFF ram_reg_1615__2_ ( .D(n7699), .CP(wclk), .Q(ram[3458]) );
  DFF ram_reg_1615__1_ ( .D(n7698), .CP(wclk), .Q(ram[3457]) );
  DFF ram_reg_1615__0_ ( .D(n7697), .CP(wclk), .Q(ram[3456]) );
  DFF ram_reg_1619__7_ ( .D(n7672), .CP(wclk), .Q(ram[3431]) );
  DFF ram_reg_1619__6_ ( .D(n7671), .CP(wclk), .Q(ram[3430]) );
  DFF ram_reg_1619__5_ ( .D(n7670), .CP(wclk), .Q(ram[3429]) );
  DFF ram_reg_1619__4_ ( .D(n7669), .CP(wclk), .Q(ram[3428]) );
  DFF ram_reg_1619__3_ ( .D(n7668), .CP(wclk), .Q(ram[3427]) );
  DFF ram_reg_1619__2_ ( .D(n7667), .CP(wclk), .Q(ram[3426]) );
  DFF ram_reg_1619__1_ ( .D(n7666), .CP(wclk), .Q(ram[3425]) );
  DFF ram_reg_1619__0_ ( .D(n7665), .CP(wclk), .Q(ram[3424]) );
  DFF ram_reg_1623__7_ ( .D(n7640), .CP(wclk), .Q(ram[3399]) );
  DFF ram_reg_1623__6_ ( .D(n7639), .CP(wclk), .Q(ram[3398]) );
  DFF ram_reg_1623__5_ ( .D(n7638), .CP(wclk), .Q(ram[3397]) );
  DFF ram_reg_1623__4_ ( .D(n7637), .CP(wclk), .Q(ram[3396]) );
  DFF ram_reg_1623__3_ ( .D(n7636), .CP(wclk), .Q(ram[3395]) );
  DFF ram_reg_1623__2_ ( .D(n7635), .CP(wclk), .Q(ram[3394]) );
  DFF ram_reg_1623__1_ ( .D(n7634), .CP(wclk), .Q(ram[3393]) );
  DFF ram_reg_1623__0_ ( .D(n7633), .CP(wclk), .Q(ram[3392]) );
  DFF ram_reg_1627__7_ ( .D(n7608), .CP(wclk), .Q(ram[3367]) );
  DFF ram_reg_1627__6_ ( .D(n7607), .CP(wclk), .Q(ram[3366]) );
  DFF ram_reg_1627__5_ ( .D(n7606), .CP(wclk), .Q(ram[3365]) );
  DFF ram_reg_1627__4_ ( .D(n7605), .CP(wclk), .Q(ram[3364]) );
  DFF ram_reg_1627__3_ ( .D(n7604), .CP(wclk), .Q(ram[3363]) );
  DFF ram_reg_1627__2_ ( .D(n7603), .CP(wclk), .Q(ram[3362]) );
  DFF ram_reg_1627__1_ ( .D(n7602), .CP(wclk), .Q(ram[3361]) );
  DFF ram_reg_1627__0_ ( .D(n7601), .CP(wclk), .Q(ram[3360]) );
  DFF ram_reg_1631__7_ ( .D(n7576), .CP(wclk), .Q(ram[3335]) );
  DFF ram_reg_1631__6_ ( .D(n7575), .CP(wclk), .Q(ram[3334]) );
  DFF ram_reg_1631__5_ ( .D(n7574), .CP(wclk), .Q(ram[3333]) );
  DFF ram_reg_1631__4_ ( .D(n7573), .CP(wclk), .Q(ram[3332]) );
  DFF ram_reg_1631__3_ ( .D(n7572), .CP(wclk), .Q(ram[3331]) );
  DFF ram_reg_1631__2_ ( .D(n7571), .CP(wclk), .Q(ram[3330]) );
  DFF ram_reg_1631__1_ ( .D(n7570), .CP(wclk), .Q(ram[3329]) );
  DFF ram_reg_1631__0_ ( .D(n7569), .CP(wclk), .Q(ram[3328]) );
  DFF ram_reg_1635__7_ ( .D(n7544), .CP(wclk), .Q(ram[3303]) );
  DFF ram_reg_1635__6_ ( .D(n7543), .CP(wclk), .Q(ram[3302]) );
  DFF ram_reg_1635__5_ ( .D(n7542), .CP(wclk), .Q(ram[3301]) );
  DFF ram_reg_1635__4_ ( .D(n7541), .CP(wclk), .Q(ram[3300]) );
  DFF ram_reg_1635__3_ ( .D(n7540), .CP(wclk), .Q(ram[3299]) );
  DFF ram_reg_1635__2_ ( .D(n7539), .CP(wclk), .Q(ram[3298]) );
  DFF ram_reg_1635__1_ ( .D(n7538), .CP(wclk), .Q(ram[3297]) );
  DFF ram_reg_1635__0_ ( .D(n7537), .CP(wclk), .Q(ram[3296]) );
  DFF ram_reg_1639__7_ ( .D(n7512), .CP(wclk), .Q(ram[3271]) );
  DFF ram_reg_1639__6_ ( .D(n7511), .CP(wclk), .Q(ram[3270]) );
  DFF ram_reg_1639__5_ ( .D(n7510), .CP(wclk), .Q(ram[3269]) );
  DFF ram_reg_1639__4_ ( .D(n7509), .CP(wclk), .Q(ram[3268]) );
  DFF ram_reg_1639__3_ ( .D(n7508), .CP(wclk), .Q(ram[3267]) );
  DFF ram_reg_1639__2_ ( .D(n7507), .CP(wclk), .Q(ram[3266]) );
  DFF ram_reg_1639__1_ ( .D(n7506), .CP(wclk), .Q(ram[3265]) );
  DFF ram_reg_1639__0_ ( .D(n7505), .CP(wclk), .Q(ram[3264]) );
  DFF ram_reg_1647__7_ ( .D(n7448), .CP(wclk), .Q(ram[3207]) );
  DFF ram_reg_1647__6_ ( .D(n7447), .CP(wclk), .Q(ram[3206]) );
  DFF ram_reg_1647__5_ ( .D(n7446), .CP(wclk), .Q(ram[3205]) );
  DFF ram_reg_1647__4_ ( .D(n7445), .CP(wclk), .Q(ram[3204]) );
  DFF ram_reg_1647__3_ ( .D(n7444), .CP(wclk), .Q(ram[3203]) );
  DFF ram_reg_1647__2_ ( .D(n7443), .CP(wclk), .Q(ram[3202]) );
  DFF ram_reg_1647__1_ ( .D(n7442), .CP(wclk), .Q(ram[3201]) );
  DFF ram_reg_1647__0_ ( .D(n7441), .CP(wclk), .Q(ram[3200]) );
  DFF ram_reg_1651__7_ ( .D(n7416), .CP(wclk), .Q(ram[3175]) );
  DFF ram_reg_1651__6_ ( .D(n7415), .CP(wclk), .Q(ram[3174]) );
  DFF ram_reg_1651__5_ ( .D(n7414), .CP(wclk), .Q(ram[3173]) );
  DFF ram_reg_1651__4_ ( .D(n7413), .CP(wclk), .Q(ram[3172]) );
  DFF ram_reg_1651__3_ ( .D(n7412), .CP(wclk), .Q(ram[3171]) );
  DFF ram_reg_1651__2_ ( .D(n7411), .CP(wclk), .Q(ram[3170]) );
  DFF ram_reg_1651__1_ ( .D(n7410), .CP(wclk), .Q(ram[3169]) );
  DFF ram_reg_1651__0_ ( .D(n7409), .CP(wclk), .Q(ram[3168]) );
  DFF ram_reg_1655__7_ ( .D(n7384), .CP(wclk), .Q(ram[3143]) );
  DFF ram_reg_1655__6_ ( .D(n7383), .CP(wclk), .Q(ram[3142]) );
  DFF ram_reg_1655__5_ ( .D(n7382), .CP(wclk), .Q(ram[3141]) );
  DFF ram_reg_1655__4_ ( .D(n7381), .CP(wclk), .Q(ram[3140]) );
  DFF ram_reg_1655__3_ ( .D(n7380), .CP(wclk), .Q(ram[3139]) );
  DFF ram_reg_1655__2_ ( .D(n7379), .CP(wclk), .Q(ram[3138]) );
  DFF ram_reg_1655__1_ ( .D(n7378), .CP(wclk), .Q(ram[3137]) );
  DFF ram_reg_1655__0_ ( .D(n7377), .CP(wclk), .Q(ram[3136]) );
  DFF ram_reg_1671__7_ ( .D(n7256), .CP(wclk), .Q(ram[3015]) );
  DFF ram_reg_1671__6_ ( .D(n7255), .CP(wclk), .Q(ram[3014]) );
  DFF ram_reg_1671__5_ ( .D(n7254), .CP(wclk), .Q(ram[3013]) );
  DFF ram_reg_1671__4_ ( .D(n7253), .CP(wclk), .Q(ram[3012]) );
  DFF ram_reg_1671__3_ ( .D(n7252), .CP(wclk), .Q(ram[3011]) );
  DFF ram_reg_1671__2_ ( .D(n7251), .CP(wclk), .Q(ram[3010]) );
  DFF ram_reg_1671__1_ ( .D(n7250), .CP(wclk), .Q(ram[3009]) );
  DFF ram_reg_1671__0_ ( .D(n7249), .CP(wclk), .Q(ram[3008]) );
  DFF ram_reg_1687__7_ ( .D(n7128), .CP(wclk), .Q(ram[2887]) );
  DFF ram_reg_1687__6_ ( .D(n7127), .CP(wclk), .Q(ram[2886]) );
  DFF ram_reg_1687__5_ ( .D(n7126), .CP(wclk), .Q(ram[2885]) );
  DFF ram_reg_1687__4_ ( .D(n7125), .CP(wclk), .Q(ram[2884]) );
  DFF ram_reg_1687__3_ ( .D(n7124), .CP(wclk), .Q(ram[2883]) );
  DFF ram_reg_1687__2_ ( .D(n7123), .CP(wclk), .Q(ram[2882]) );
  DFF ram_reg_1687__1_ ( .D(n7122), .CP(wclk), .Q(ram[2881]) );
  DFF ram_reg_1687__0_ ( .D(n7121), .CP(wclk), .Q(ram[2880]) );
  DFF ram_reg_1735__7_ ( .D(n6744), .CP(wclk), .Q(ram[2503]) );
  DFF ram_reg_1735__6_ ( .D(n6743), .CP(wclk), .Q(ram[2502]) );
  DFF ram_reg_1735__5_ ( .D(n6742), .CP(wclk), .Q(ram[2501]) );
  DFF ram_reg_1735__4_ ( .D(n6741), .CP(wclk), .Q(ram[2500]) );
  DFF ram_reg_1735__3_ ( .D(n6740), .CP(wclk), .Q(ram[2499]) );
  DFF ram_reg_1735__2_ ( .D(n6739), .CP(wclk), .Q(ram[2498]) );
  DFF ram_reg_1735__1_ ( .D(n6738), .CP(wclk), .Q(ram[2497]) );
  DFF ram_reg_1735__0_ ( .D(n6737), .CP(wclk), .Q(ram[2496]) );
  DFF ram_reg_1747__7_ ( .D(n6648), .CP(wclk), .Q(ram[2407]) );
  DFF ram_reg_1747__6_ ( .D(n6647), .CP(wclk), .Q(ram[2406]) );
  DFF ram_reg_1747__5_ ( .D(n6646), .CP(wclk), .Q(ram[2405]) );
  DFF ram_reg_1747__4_ ( .D(n6645), .CP(wclk), .Q(ram[2404]) );
  DFF ram_reg_1747__3_ ( .D(n6644), .CP(wclk), .Q(ram[2403]) );
  DFF ram_reg_1747__2_ ( .D(n6643), .CP(wclk), .Q(ram[2402]) );
  DFF ram_reg_1747__1_ ( .D(n6642), .CP(wclk), .Q(ram[2401]) );
  DFF ram_reg_1747__0_ ( .D(n6641), .CP(wclk), .Q(ram[2400]) );
  DFF ram_reg_1751__7_ ( .D(n6616), .CP(wclk), .Q(ram[2375]) );
  DFF ram_reg_1751__6_ ( .D(n6615), .CP(wclk), .Q(ram[2374]) );
  DFF ram_reg_1751__5_ ( .D(n6614), .CP(wclk), .Q(ram[2373]) );
  DFF ram_reg_1751__4_ ( .D(n6613), .CP(wclk), .Q(ram[2372]) );
  DFF ram_reg_1751__3_ ( .D(n6612), .CP(wclk), .Q(ram[2371]) );
  DFF ram_reg_1751__2_ ( .D(n6611), .CP(wclk), .Q(ram[2370]) );
  DFF ram_reg_1751__1_ ( .D(n6610), .CP(wclk), .Q(ram[2369]) );
  DFF ram_reg_1751__0_ ( .D(n6609), .CP(wclk), .Q(ram[2368]) );
  DFF ram_reg_1767__7_ ( .D(n6488), .CP(wclk), .Q(ram[2247]) );
  DFF ram_reg_1767__6_ ( .D(n6487), .CP(wclk), .Q(ram[2246]) );
  DFF ram_reg_1767__5_ ( .D(n6486), .CP(wclk), .Q(ram[2245]) );
  DFF ram_reg_1767__4_ ( .D(n6485), .CP(wclk), .Q(ram[2244]) );
  DFF ram_reg_1767__3_ ( .D(n6484), .CP(wclk), .Q(ram[2243]) );
  DFF ram_reg_1767__2_ ( .D(n6483), .CP(wclk), .Q(ram[2242]) );
  DFF ram_reg_1767__1_ ( .D(n6482), .CP(wclk), .Q(ram[2241]) );
  DFF ram_reg_1767__0_ ( .D(n6481), .CP(wclk), .Q(ram[2240]) );
  DFF ram_reg_1795__7_ ( .D(n6264), .CP(wclk), .Q(ram[2023]) );
  DFF ram_reg_1795__6_ ( .D(n6263), .CP(wclk), .Q(ram[2022]) );
  DFF ram_reg_1795__5_ ( .D(n6262), .CP(wclk), .Q(ram[2021]) );
  DFF ram_reg_1795__4_ ( .D(n6261), .CP(wclk), .Q(ram[2020]) );
  DFF ram_reg_1795__3_ ( .D(n6260), .CP(wclk), .Q(ram[2019]) );
  DFF ram_reg_1795__2_ ( .D(n6259), .CP(wclk), .Q(ram[2018]) );
  DFF ram_reg_1795__1_ ( .D(n6258), .CP(wclk), .Q(ram[2017]) );
  DFF ram_reg_1795__0_ ( .D(n6257), .CP(wclk), .Q(ram[2016]) );
  DFF ram_reg_1799__7_ ( .D(n6232), .CP(wclk), .Q(ram[1991]) );
  DFF ram_reg_1799__6_ ( .D(n6231), .CP(wclk), .Q(ram[1990]) );
  DFF ram_reg_1799__5_ ( .D(n6230), .CP(wclk), .Q(ram[1989]) );
  DFF ram_reg_1799__4_ ( .D(n6229), .CP(wclk), .Q(ram[1988]) );
  DFF ram_reg_1799__3_ ( .D(n6228), .CP(wclk), .Q(ram[1987]) );
  DFF ram_reg_1799__2_ ( .D(n6227), .CP(wclk), .Q(ram[1986]) );
  DFF ram_reg_1799__1_ ( .D(n6226), .CP(wclk), .Q(ram[1985]) );
  DFF ram_reg_1799__0_ ( .D(n6225), .CP(wclk), .Q(ram[1984]) );
  DFF ram_reg_1811__7_ ( .D(n6136), .CP(wclk), .Q(ram[1895]) );
  DFF ram_reg_1811__6_ ( .D(n6135), .CP(wclk), .Q(ram[1894]) );
  DFF ram_reg_1811__5_ ( .D(n6134), .CP(wclk), .Q(ram[1893]) );
  DFF ram_reg_1811__4_ ( .D(n6133), .CP(wclk), .Q(ram[1892]) );
  DFF ram_reg_1811__3_ ( .D(n6132), .CP(wclk), .Q(ram[1891]) );
  DFF ram_reg_1811__2_ ( .D(n6131), .CP(wclk), .Q(ram[1890]) );
  DFF ram_reg_1811__1_ ( .D(n6130), .CP(wclk), .Q(ram[1889]) );
  DFF ram_reg_1811__0_ ( .D(n6129), .CP(wclk), .Q(ram[1888]) );
  DFF ram_reg_1815__7_ ( .D(n6104), .CP(wclk), .Q(ram[1863]) );
  DFF ram_reg_1815__6_ ( .D(n6103), .CP(wclk), .Q(ram[1862]) );
  DFF ram_reg_1815__5_ ( .D(n6102), .CP(wclk), .Q(ram[1861]) );
  DFF ram_reg_1815__4_ ( .D(n6101), .CP(wclk), .Q(ram[1860]) );
  DFF ram_reg_1815__3_ ( .D(n6100), .CP(wclk), .Q(ram[1859]) );
  DFF ram_reg_1815__2_ ( .D(n6099), .CP(wclk), .Q(ram[1858]) );
  DFF ram_reg_1815__1_ ( .D(n6098), .CP(wclk), .Q(ram[1857]) );
  DFF ram_reg_1815__0_ ( .D(n6097), .CP(wclk), .Q(ram[1856]) );
  DFF ram_reg_1831__7_ ( .D(n5976), .CP(wclk), .Q(ram[1735]) );
  DFF ram_reg_1831__6_ ( .D(n5975), .CP(wclk), .Q(ram[1734]) );
  DFF ram_reg_1831__5_ ( .D(n5974), .CP(wclk), .Q(ram[1733]) );
  DFF ram_reg_1831__4_ ( .D(n5973), .CP(wclk), .Q(ram[1732]) );
  DFF ram_reg_1831__3_ ( .D(n5972), .CP(wclk), .Q(ram[1731]) );
  DFF ram_reg_1831__2_ ( .D(n5971), .CP(wclk), .Q(ram[1730]) );
  DFF ram_reg_1831__1_ ( .D(n5970), .CP(wclk), .Q(ram[1729]) );
  DFF ram_reg_1831__0_ ( .D(n5969), .CP(wclk), .Q(ram[1728]) );
  DFF ram_reg_1847__7_ ( .D(n5848), .CP(wclk), .Q(ram[1607]) );
  DFF ram_reg_1847__6_ ( .D(n5847), .CP(wclk), .Q(ram[1606]) );
  DFF ram_reg_1847__5_ ( .D(n5846), .CP(wclk), .Q(ram[1605]) );
  DFF ram_reg_1847__4_ ( .D(n5845), .CP(wclk), .Q(ram[1604]) );
  DFF ram_reg_1847__3_ ( .D(n5844), .CP(wclk), .Q(ram[1603]) );
  DFF ram_reg_1847__2_ ( .D(n5843), .CP(wclk), .Q(ram[1602]) );
  DFF ram_reg_1847__1_ ( .D(n5842), .CP(wclk), .Q(ram[1601]) );
  DFF ram_reg_1847__0_ ( .D(n5841), .CP(wclk), .Q(ram[1600]) );
  DFF ram_reg_1859__7_ ( .D(n5752), .CP(wclk), .Q(ram[1511]) );
  DFF ram_reg_1859__6_ ( .D(n5751), .CP(wclk), .Q(ram[1510]) );
  DFF ram_reg_1859__5_ ( .D(n5750), .CP(wclk), .Q(ram[1509]) );
  DFF ram_reg_1859__4_ ( .D(n5749), .CP(wclk), .Q(ram[1508]) );
  DFF ram_reg_1859__3_ ( .D(n5748), .CP(wclk), .Q(ram[1507]) );
  DFF ram_reg_1859__2_ ( .D(n5747), .CP(wclk), .Q(ram[1506]) );
  DFF ram_reg_1859__1_ ( .D(n5746), .CP(wclk), .Q(ram[1505]) );
  DFF ram_reg_1859__0_ ( .D(n5745), .CP(wclk), .Q(ram[1504]) );
  DFF ram_reg_1863__7_ ( .D(n5720), .CP(wclk), .Q(ram[1479]) );
  DFF ram_reg_1863__6_ ( .D(n5719), .CP(wclk), .Q(ram[1478]) );
  DFF ram_reg_1863__5_ ( .D(n5718), .CP(wclk), .Q(ram[1477]) );
  DFF ram_reg_1863__4_ ( .D(n5717), .CP(wclk), .Q(ram[1476]) );
  DFF ram_reg_1863__3_ ( .D(n5716), .CP(wclk), .Q(ram[1475]) );
  DFF ram_reg_1863__2_ ( .D(n5715), .CP(wclk), .Q(ram[1474]) );
  DFF ram_reg_1863__1_ ( .D(n5714), .CP(wclk), .Q(ram[1473]) );
  DFF ram_reg_1863__0_ ( .D(n5713), .CP(wclk), .Q(ram[1472]) );
  DFF ram_reg_1871__7_ ( .D(n5656), .CP(wclk), .Q(ram[1415]) );
  DFF ram_reg_1871__6_ ( .D(n5655), .CP(wclk), .Q(ram[1414]) );
  DFF ram_reg_1871__5_ ( .D(n5654), .CP(wclk), .Q(ram[1413]) );
  DFF ram_reg_1871__4_ ( .D(n5653), .CP(wclk), .Q(ram[1412]) );
  DFF ram_reg_1871__3_ ( .D(n5652), .CP(wclk), .Q(ram[1411]) );
  DFF ram_reg_1871__2_ ( .D(n5651), .CP(wclk), .Q(ram[1410]) );
  DFF ram_reg_1871__1_ ( .D(n5650), .CP(wclk), .Q(ram[1409]) );
  DFF ram_reg_1871__0_ ( .D(n5649), .CP(wclk), .Q(ram[1408]) );
  DFF ram_reg_1875__7_ ( .D(n5624), .CP(wclk), .Q(ram[1383]) );
  DFF ram_reg_1875__6_ ( .D(n5623), .CP(wclk), .Q(ram[1382]) );
  DFF ram_reg_1875__5_ ( .D(n5622), .CP(wclk), .Q(ram[1381]) );
  DFF ram_reg_1875__4_ ( .D(n5621), .CP(wclk), .Q(ram[1380]) );
  DFF ram_reg_1875__3_ ( .D(n5620), .CP(wclk), .Q(ram[1379]) );
  DFF ram_reg_1875__2_ ( .D(n5619), .CP(wclk), .Q(ram[1378]) );
  DFF ram_reg_1875__1_ ( .D(n5618), .CP(wclk), .Q(ram[1377]) );
  DFF ram_reg_1875__0_ ( .D(n5617), .CP(wclk), .Q(ram[1376]) );
  DFF ram_reg_1879__7_ ( .D(n5592), .CP(wclk), .Q(ram[1351]) );
  DFF ram_reg_1879__6_ ( .D(n5591), .CP(wclk), .Q(ram[1350]) );
  DFF ram_reg_1879__5_ ( .D(n5590), .CP(wclk), .Q(ram[1349]) );
  DFF ram_reg_1879__4_ ( .D(n5589), .CP(wclk), .Q(ram[1348]) );
  DFF ram_reg_1879__3_ ( .D(n5588), .CP(wclk), .Q(ram[1347]) );
  DFF ram_reg_1879__2_ ( .D(n5587), .CP(wclk), .Q(ram[1346]) );
  DFF ram_reg_1879__1_ ( .D(n5586), .CP(wclk), .Q(ram[1345]) );
  DFF ram_reg_1879__0_ ( .D(n5585), .CP(wclk), .Q(ram[1344]) );
  DFF ram_reg_1883__7_ ( .D(n5560), .CP(wclk), .Q(ram[1319]) );
  DFF ram_reg_1883__6_ ( .D(n5559), .CP(wclk), .Q(ram[1318]) );
  DFF ram_reg_1883__5_ ( .D(n5558), .CP(wclk), .Q(ram[1317]) );
  DFF ram_reg_1883__4_ ( .D(n5557), .CP(wclk), .Q(ram[1316]) );
  DFF ram_reg_1883__3_ ( .D(n5556), .CP(wclk), .Q(ram[1315]) );
  DFF ram_reg_1883__2_ ( .D(n5555), .CP(wclk), .Q(ram[1314]) );
  DFF ram_reg_1883__1_ ( .D(n5554), .CP(wclk), .Q(ram[1313]) );
  DFF ram_reg_1883__0_ ( .D(n5553), .CP(wclk), .Q(ram[1312]) );
  DFF ram_reg_1887__7_ ( .D(n5528), .CP(wclk), .Q(ram[1287]) );
  DFF ram_reg_1887__6_ ( .D(n5527), .CP(wclk), .Q(ram[1286]) );
  DFF ram_reg_1887__5_ ( .D(n5526), .CP(wclk), .Q(ram[1285]) );
  DFF ram_reg_1887__4_ ( .D(n5525), .CP(wclk), .Q(ram[1284]) );
  DFF ram_reg_1887__3_ ( .D(n5524), .CP(wclk), .Q(ram[1283]) );
  DFF ram_reg_1887__2_ ( .D(n5523), .CP(wclk), .Q(ram[1282]) );
  DFF ram_reg_1887__1_ ( .D(n5522), .CP(wclk), .Q(ram[1281]) );
  DFF ram_reg_1887__0_ ( .D(n5521), .CP(wclk), .Q(ram[1280]) );
  DFF ram_reg_1891__7_ ( .D(n5496), .CP(wclk), .Q(ram[1255]) );
  DFF ram_reg_1891__6_ ( .D(n5495), .CP(wclk), .Q(ram[1254]) );
  DFF ram_reg_1891__5_ ( .D(n5494), .CP(wclk), .Q(ram[1253]) );
  DFF ram_reg_1891__4_ ( .D(n5493), .CP(wclk), .Q(ram[1252]) );
  DFF ram_reg_1891__3_ ( .D(n5492), .CP(wclk), .Q(ram[1251]) );
  DFF ram_reg_1891__2_ ( .D(n5491), .CP(wclk), .Q(ram[1250]) );
  DFF ram_reg_1891__1_ ( .D(n5490), .CP(wclk), .Q(ram[1249]) );
  DFF ram_reg_1891__0_ ( .D(n5489), .CP(wclk), .Q(ram[1248]) );
  DFF ram_reg_1895__7_ ( .D(n5464), .CP(wclk), .Q(ram[1223]) );
  DFF ram_reg_1895__6_ ( .D(n5463), .CP(wclk), .Q(ram[1222]) );
  DFF ram_reg_1895__5_ ( .D(n5462), .CP(wclk), .Q(ram[1221]) );
  DFF ram_reg_1895__4_ ( .D(n5461), .CP(wclk), .Q(ram[1220]) );
  DFF ram_reg_1895__3_ ( .D(n5460), .CP(wclk), .Q(ram[1219]) );
  DFF ram_reg_1895__2_ ( .D(n5459), .CP(wclk), .Q(ram[1218]) );
  DFF ram_reg_1895__1_ ( .D(n5458), .CP(wclk), .Q(ram[1217]) );
  DFF ram_reg_1895__0_ ( .D(n5457), .CP(wclk), .Q(ram[1216]) );
  DFF ram_reg_1907__7_ ( .D(n5368), .CP(wclk), .Q(ram[1127]) );
  DFF ram_reg_1907__6_ ( .D(n5367), .CP(wclk), .Q(ram[1126]) );
  DFF ram_reg_1907__5_ ( .D(n5366), .CP(wclk), .Q(ram[1125]) );
  DFF ram_reg_1907__4_ ( .D(n5365), .CP(wclk), .Q(ram[1124]) );
  DFF ram_reg_1907__3_ ( .D(n5364), .CP(wclk), .Q(ram[1123]) );
  DFF ram_reg_1907__2_ ( .D(n5363), .CP(wclk), .Q(ram[1122]) );
  DFF ram_reg_1907__1_ ( .D(n5362), .CP(wclk), .Q(ram[1121]) );
  DFF ram_reg_1907__0_ ( .D(n5361), .CP(wclk), .Q(ram[1120]) );
  DFF ram_reg_1911__7_ ( .D(n5336), .CP(wclk), .Q(ram[1095]) );
  DFF ram_reg_1911__6_ ( .D(n5335), .CP(wclk), .Q(ram[1094]) );
  DFF ram_reg_1911__5_ ( .D(n5334), .CP(wclk), .Q(ram[1093]) );
  DFF ram_reg_1911__4_ ( .D(n5333), .CP(wclk), .Q(ram[1092]) );
  DFF ram_reg_1911__3_ ( .D(n5332), .CP(wclk), .Q(ram[1091]) );
  DFF ram_reg_1911__2_ ( .D(n5331), .CP(wclk), .Q(ram[1090]) );
  DFF ram_reg_1911__1_ ( .D(n5330), .CP(wclk), .Q(ram[1089]) );
  DFF ram_reg_1911__0_ ( .D(n5329), .CP(wclk), .Q(ram[1088]) );
  DFF ram_reg_1943__7_ ( .D(n5080), .CP(wclk), .Q(ram[839]) );
  DFF ram_reg_1943__6_ ( .D(n5079), .CP(wclk), .Q(ram[838]) );
  DFF ram_reg_1943__5_ ( .D(n5078), .CP(wclk), .Q(ram[837]) );
  DFF ram_reg_1943__4_ ( .D(n5077), .CP(wclk), .Q(ram[836]) );
  DFF ram_reg_1943__3_ ( .D(n5076), .CP(wclk), .Q(ram[835]) );
  DFF ram_reg_1943__2_ ( .D(n5075), .CP(wclk), .Q(ram[834]) );
  DFF ram_reg_1943__1_ ( .D(n5074), .CP(wclk), .Q(ram[833]) );
  DFF ram_reg_1943__0_ ( .D(n5073), .CP(wclk), .Q(ram[832]) );
  DFF ram_reg_1991__7_ ( .D(n4696), .CP(wclk), .Q(ram[455]) );
  DFF ram_reg_1991__6_ ( .D(n4695), .CP(wclk), .Q(ram[454]) );
  DFF ram_reg_1991__5_ ( .D(n4694), .CP(wclk), .Q(ram[453]) );
  DFF ram_reg_1991__4_ ( .D(n4693), .CP(wclk), .Q(ram[452]) );
  DFF ram_reg_1991__3_ ( .D(n4692), .CP(wclk), .Q(ram[451]) );
  DFF ram_reg_1991__2_ ( .D(n4691), .CP(wclk), .Q(ram[450]) );
  DFF ram_reg_1991__1_ ( .D(n4690), .CP(wclk), .Q(ram[449]) );
  DFF ram_reg_1991__0_ ( .D(n4689), .CP(wclk), .Q(ram[448]) );
  DFF ram_reg_2007__7_ ( .D(n4568), .CP(wclk), .Q(ram[327]) );
  DFF ram_reg_2007__6_ ( .D(n4567), .CP(wclk), .Q(ram[326]) );
  DFF ram_reg_2007__5_ ( .D(n4566), .CP(wclk), .Q(ram[325]) );
  DFF ram_reg_2007__4_ ( .D(n4565), .CP(wclk), .Q(ram[324]) );
  DFF ram_reg_2007__3_ ( .D(n4564), .CP(wclk), .Q(ram[323]) );
  DFF ram_reg_2007__2_ ( .D(n4563), .CP(wclk), .Q(ram[322]) );
  DFF ram_reg_2007__1_ ( .D(n4562), .CP(wclk), .Q(ram[321]) );
  DFF ram_reg_2007__0_ ( .D(n4561), .CP(wclk), .Q(ram[320]) );
  AND2 U2 ( .A1(n4226), .A2(n4112), .Z(n1) );
  AND2 U3 ( .A1(n4226), .A2(n4115), .Z(n2) );
  AND2 U4 ( .A1(n4226), .A2(n4118), .Z(n3) );
  AND2 U5 ( .A1(n4226), .A2(n4121), .Z(n4) );
  AND2 U6 ( .A1(n4103), .A2(n4100), .Z(n5) );
  AND2 U7 ( .A1(n4106), .A2(n4100), .Z(n6) );
  AND2 U8 ( .A1(n4109), .A2(n4100), .Z(n7) );
  AND2 U9 ( .A1(n4112), .A2(n4100), .Z(n8) );
  AND2 U10 ( .A1(n4115), .A2(n4100), .Z(n9) );
  AND2 U11 ( .A1(n4209), .A2(n4099), .Z(n10) );
  AND2 U12 ( .A1(n4209), .A2(n4103), .Z(n11) );
  AND2 U13 ( .A1(n4209), .A2(n4106), .Z(n12) );
  AND2 U14 ( .A1(n4209), .A2(n4109), .Z(n24) );
  AND2 U15 ( .A1(n4209), .A2(n4112), .Z(n27) );
  AND2 U16 ( .A1(n4209), .A2(n4115), .Z(n30) );
  AND2 U17 ( .A1(n4209), .A2(n4118), .Z(n33) );
  AND2 U18 ( .A1(n4209), .A2(n4121), .Z(n36) );
  AND2 U19 ( .A1(n4226), .A2(n4099), .Z(n39) );
  AND2 U20 ( .A1(n4226), .A2(n4103), .Z(n168) );
  AND2 U21 ( .A1(n4226), .A2(n4106), .Z(n171) );
  AND2 U22 ( .A1(n4226), .A2(n4109), .Z(n174) );
  NAND2 U23 ( .A1(n345), .A2(n215), .ZN(n177) );
  NAND2 U24 ( .A1(n475), .A2(n215), .ZN(n180) );
  NAND2 U25 ( .A1(n605), .A2(n215), .ZN(n183) );
  NAND2 U26 ( .A1(n735), .A2(n215), .ZN(n186) );
  NAND2 U27 ( .A1(n865), .A2(n215), .ZN(n189) );
  NAND2 U28 ( .A1(n995), .A2(n215), .ZN(n192) );
  NAND2 U29 ( .A1(n1125), .A2(n215), .ZN(n195) );
  NAND2 U30 ( .A1(n214), .A2(n215), .ZN(n198) );
  NAND2 U31 ( .A1(n1255), .A2(n214), .ZN(n201) );
  NAND2 U32 ( .A1(n1255), .A2(n345), .ZN(n204) );
  NAND2 U33 ( .A1(n1255), .A2(n475), .ZN(n207) );
  NAND2 U34 ( .A1(n1255), .A2(n605), .ZN(n210) );
  NAND2 U35 ( .A1(n1255), .A2(n735), .ZN(n213) );
  NAND2 U36 ( .A1(n1255), .A2(n865), .ZN(n218) );
  NAND2 U37 ( .A1(n1255), .A2(n995), .ZN(n348) );
  NAND2 U38 ( .A1(n1255), .A2(n1125), .ZN(n478) );
  NAND2 U39 ( .A1(n2288), .A2(n214), .ZN(n608) );
  NAND2 U40 ( .A1(n2288), .A2(n345), .ZN(n738) );
  NAND2 U41 ( .A1(n2288), .A2(n475), .ZN(n868) );
  NAND2 U42 ( .A1(n2288), .A2(n605), .ZN(n998) );
  NAND2 U43 ( .A1(n2288), .A2(n735), .ZN(n1128) );
  NAND2 U44 ( .A1(n2288), .A2(n865), .ZN(n1258) );
  NAND2 U45 ( .A1(n2288), .A2(n995), .ZN(n1387) );
  NAND2 U46 ( .A1(n2288), .A2(n1125), .ZN(n1516) );
  NAND2 U47 ( .A1(n3321), .A2(n214), .ZN(n1645) );
  NAND2 U48 ( .A1(n3321), .A2(n345), .ZN(n1774) );
  NAND2 U49 ( .A1(n3321), .A2(n475), .ZN(n1903) );
  NAND2 U50 ( .A1(n3321), .A2(n605), .ZN(n2032) );
  NAND2 U51 ( .A1(n3321), .A2(n735), .ZN(n2161) );
  NAND2 U52 ( .A1(n3321), .A2(n865), .ZN(n2291) );
  NAND2 U53 ( .A1(n3321), .A2(n995), .ZN(n2420) );
  NAND2 U54 ( .A1(n3321), .A2(n1125), .ZN(n2549) );
  MUX31 U55 ( .I0(n21296), .I1(n21125), .I2(n20954), .S0(raddr[9]), .S1(
        raddr[10]), .Z(N36) );
  MUX31 U56 ( .I0(n20949), .I1(n20864), .I2(n20783), .S0(n29321), .S1(
        raddr[9]), .Z(n20954) );
  MUX31 U57 ( .I0(n21980), .I1(n21809), .I2(n21638), .S0(raddr[9]), .S1(
        raddr[10]), .Z(N35) );
  MUX31 U58 ( .I0(n21633), .I1(n21548), .I2(n21467), .S0(n29321), .S1(
        raddr[9]), .Z(n21638) );
  MUX31 U59 ( .I0(n22664), .I1(n22493), .I2(n22322), .S0(raddr[9]), .S1(
        raddr[10]), .Z(N34) );
  MUX31 U60 ( .I0(n22317), .I1(n22232), .I2(n22151), .S0(n29321), .S1(
        raddr[9]), .Z(n22322) );
  MUX31 U61 ( .I0(n23348), .I1(n23177), .I2(n23006), .S0(raddr[9]), .S1(
        raddr[10]), .Z(N33) );
  MUX31 U62 ( .I0(n23001), .I1(n22916), .I2(n22835), .S0(n29321), .S1(
        raddr[9]), .Z(n23006) );
  MUX31 U63 ( .I0(n24032), .I1(n23861), .I2(n23690), .S0(raddr[9]), .S1(
        raddr[10]), .Z(N32) );
  MUX31 U64 ( .I0(n23685), .I1(n23600), .I2(n23519), .S0(n29321), .S1(
        raddr[9]), .Z(n23690) );
  MUX31 U65 ( .I0(n24716), .I1(n24545), .I2(n24374), .S0(raddr[9]), .S1(
        raddr[10]), .Z(N31) );
  MUX31 U66 ( .I0(n24369), .I1(n24284), .I2(n24203), .S0(n29321), .S1(
        raddr[9]), .Z(n24374) );
  MUX31 U67 ( .I0(n25400), .I1(n25229), .I2(n25058), .S0(raddr[9]), .S1(
        raddr[10]), .Z(N30) );
  MUX31 U68 ( .I0(n25053), .I1(n24968), .I2(n24887), .S0(n29321), .S1(
        raddr[9]), .Z(n25058) );
  MUX31 U69 ( .I0(n26084), .I1(n25913), .I2(n25742), .S0(raddr[9]), .S1(
        raddr[10]), .Z(N29) );
  MUX31 U70 ( .I0(n25737), .I1(n25652), .I2(n25571), .S0(n29321), .S1(
        raddr[9]), .Z(n25742) );
  INV U71 ( .I(n177), .ZN(n27431) );
  INV U72 ( .I(n177), .ZN(n27432) );
  INV U73 ( .I(n177), .ZN(n27433) );
  INV U74 ( .I(n180), .ZN(n27428) );
  INV U75 ( .I(n180), .ZN(n27429) );
  INV U76 ( .I(n180), .ZN(n27430) );
  INV U77 ( .I(n183), .ZN(n27425) );
  INV U78 ( .I(n183), .ZN(n27426) );
  INV U79 ( .I(n183), .ZN(n27427) );
  INV U80 ( .I(n186), .ZN(n27422) );
  INV U81 ( .I(n186), .ZN(n27423) );
  INV U82 ( .I(n186), .ZN(n27424) );
  INV U83 ( .I(n189), .ZN(n27419) );
  INV U84 ( .I(n189), .ZN(n27420) );
  INV U85 ( .I(n189), .ZN(n27421) );
  INV U86 ( .I(n192), .ZN(n27416) );
  INV U87 ( .I(n192), .ZN(n27417) );
  INV U88 ( .I(n192), .ZN(n27418) );
  INV U89 ( .I(n195), .ZN(n27413) );
  INV U90 ( .I(n195), .ZN(n27414) );
  INV U91 ( .I(n195), .ZN(n27415) );
  INV U92 ( .I(n201), .ZN(n27410) );
  INV U93 ( .I(n201), .ZN(n27411) );
  INV U94 ( .I(n201), .ZN(n27412) );
  INV U95 ( .I(n204), .ZN(n27407) );
  INV U96 ( .I(n204), .ZN(n27408) );
  INV U97 ( .I(n204), .ZN(n27409) );
  INV U98 ( .I(n207), .ZN(n27404) );
  INV U99 ( .I(n207), .ZN(n27405) );
  INV U100 ( .I(n207), .ZN(n27406) );
  INV U101 ( .I(n210), .ZN(n27401) );
  INV U102 ( .I(n210), .ZN(n27402) );
  INV U103 ( .I(n210), .ZN(n27403) );
  INV U104 ( .I(n213), .ZN(n27398) );
  INV U105 ( .I(n213), .ZN(n27399) );
  INV U106 ( .I(n213), .ZN(n27400) );
  INV U107 ( .I(n218), .ZN(n27395) );
  INV U108 ( .I(n218), .ZN(n27396) );
  INV U109 ( .I(n218), .ZN(n27397) );
  INV U110 ( .I(n348), .ZN(n27392) );
  INV U111 ( .I(n348), .ZN(n27393) );
  INV U112 ( .I(n348), .ZN(n27394) );
  INV U113 ( .I(n478), .ZN(n27389) );
  INV U114 ( .I(n478), .ZN(n27390) );
  INV U115 ( .I(n478), .ZN(n27391) );
  INV U116 ( .I(n608), .ZN(n27386) );
  INV U117 ( .I(n608), .ZN(n27387) );
  INV U118 ( .I(n608), .ZN(n27388) );
  INV U119 ( .I(n738), .ZN(n27383) );
  INV U120 ( .I(n738), .ZN(n27384) );
  INV U121 ( .I(n738), .ZN(n27385) );
  INV U122 ( .I(n868), .ZN(n27380) );
  INV U123 ( .I(n868), .ZN(n27381) );
  INV U124 ( .I(n868), .ZN(n27382) );
  INV U125 ( .I(n998), .ZN(n27377) );
  INV U126 ( .I(n998), .ZN(n27378) );
  INV U127 ( .I(n998), .ZN(n27379) );
  INV U128 ( .I(n1516), .ZN(n27365) );
  INV U129 ( .I(n1516), .ZN(n27366) );
  INV U130 ( .I(n1516), .ZN(n27367) );
  INV U131 ( .I(n2549), .ZN(n27341) );
  INV U132 ( .I(n2549), .ZN(n27342) );
  INV U133 ( .I(n2549), .ZN(n27343) );
  NOR3 U134 ( .A1(waddr[1]), .A2(waddr[2]), .A3(n29582), .ZN(n4118) );
  NOR3 U135 ( .A1(waddr[1]), .A2(waddr[2]), .A3(waddr[0]), .ZN(n4121) );
  NOR3 U136 ( .A1(waddr[0]), .A2(waddr[1]), .A3(n29584), .ZN(n4109) );
  NOR3 U137 ( .A1(waddr[0]), .A2(waddr[2]), .A3(n29583), .ZN(n4115) );
  NOR3 U138 ( .A1(n29582), .A2(waddr[1]), .A3(n29584), .ZN(n4106) );
  NOR3 U139 ( .A1(n29583), .A2(waddr[0]), .A3(n29584), .ZN(n4103) );
  NOR3 U140 ( .A1(n29582), .A2(waddr[2]), .A3(n29583), .ZN(n4112) );
  I_NAND2 U141 ( .A1(n13), .B1(n29407), .ZN(n15) );
  BUF U142 ( .I(n29533), .Z(n29376) );
  BUF U143 ( .I(n29532), .Z(n29377) );
  BUF U144 ( .I(n29532), .Z(n29378) );
  BUF U145 ( .I(n29532), .Z(n29379) );
  BUF U146 ( .I(n29531), .Z(n29380) );
  BUF U147 ( .I(n29531), .Z(n29381) );
  BUF U148 ( .I(n29531), .Z(n29382) );
  BUF U149 ( .I(n29530), .Z(n29383) );
  BUF U150 ( .I(n29530), .Z(n29384) );
  BUF U151 ( .I(n29530), .Z(n29385) );
  BUF U152 ( .I(n29536), .Z(n29365) );
  BUF U153 ( .I(n29536), .Z(n29366) );
  BUF U154 ( .I(n29536), .Z(n29367) );
  BUF U155 ( .I(n29535), .Z(n29368) );
  BUF U156 ( .I(n29535), .Z(n29369) );
  BUF U157 ( .I(n29535), .Z(n29370) );
  BUF U158 ( .I(n29534), .Z(n29371) );
  BUF U159 ( .I(n29534), .Z(n29372) );
  BUF U160 ( .I(n29534), .Z(n29373) );
  BUF U161 ( .I(n29533), .Z(n29374) );
  BUF U162 ( .I(n29533), .Z(n29375) );
  BUF U163 ( .I(n29526), .Z(n29397) );
  BUF U164 ( .I(n29525), .Z(n29398) );
  BUF U165 ( .I(n29525), .Z(n29399) );
  BUF U166 ( .I(n29525), .Z(n29400) );
  BUF U167 ( .I(n29524), .Z(n29401) );
  BUF U168 ( .I(n29524), .Z(n29402) );
  BUF U169 ( .I(n29524), .Z(n29403) );
  BUF U170 ( .I(n29523), .Z(n29404) );
  BUF U171 ( .I(n29523), .Z(n29405) );
  BUF U172 ( .I(n29523), .Z(n29406) );
  BUF U173 ( .I(n29529), .Z(n29386) );
  BUF U174 ( .I(n29529), .Z(n29387) );
  BUF U175 ( .I(n29529), .Z(n29388) );
  BUF U176 ( .I(n29528), .Z(n29389) );
  BUF U177 ( .I(n29528), .Z(n29390) );
  BUF U178 ( .I(n29528), .Z(n29391) );
  BUF U179 ( .I(n29527), .Z(n29392) );
  BUF U180 ( .I(n29527), .Z(n29393) );
  BUF U181 ( .I(n29527), .Z(n29394) );
  BUF U182 ( .I(n29526), .Z(n29395) );
  BUF U183 ( .I(n29526), .Z(n29396) );
  BUF U184 ( .I(n29547), .Z(n29333) );
  BUF U185 ( .I(n29547), .Z(n29334) );
  BUF U186 ( .I(n29546), .Z(n29335) );
  BUF U187 ( .I(n29546), .Z(n29336) );
  BUF U188 ( .I(n29546), .Z(n29337) );
  BUF U189 ( .I(n29545), .Z(n29338) );
  BUF U190 ( .I(n29545), .Z(n29339) );
  BUF U191 ( .I(n29545), .Z(n29340) );
  BUF U192 ( .I(n29544), .Z(n29341) );
  BUF U193 ( .I(n29544), .Z(n29342) );
  BUF U194 ( .I(n29550), .Z(n29323) );
  BUF U195 ( .I(n29550), .Z(n29324) );
  BUF U196 ( .I(n29550), .Z(n29325) );
  BUF U197 ( .I(n29549), .Z(n29326) );
  BUF U198 ( .I(n29549), .Z(n29327) );
  BUF U199 ( .I(n29549), .Z(n29328) );
  BUF U200 ( .I(n29548), .Z(n29329) );
  BUF U201 ( .I(n29548), .Z(n29330) );
  BUF U202 ( .I(n29548), .Z(n29331) );
  BUF U203 ( .I(n29547), .Z(n29332) );
  BUF U204 ( .I(n29540), .Z(n29355) );
  BUF U205 ( .I(n29539), .Z(n29356) );
  BUF U206 ( .I(n29539), .Z(n29357) );
  BUF U207 ( .I(n29539), .Z(n29358) );
  BUF U208 ( .I(n29538), .Z(n29359) );
  BUF U209 ( .I(n29538), .Z(n29360) );
  BUF U210 ( .I(n29538), .Z(n29361) );
  BUF U211 ( .I(n29537), .Z(n29362) );
  BUF U212 ( .I(n29537), .Z(n29363) );
  BUF U213 ( .I(n29544), .Z(n29343) );
  BUF U214 ( .I(n29543), .Z(n29344) );
  BUF U215 ( .I(n29543), .Z(n29345) );
  BUF U216 ( .I(n29543), .Z(n29346) );
  BUF U217 ( .I(n29542), .Z(n29347) );
  BUF U218 ( .I(n29542), .Z(n29348) );
  BUF U219 ( .I(n29542), .Z(n29349) );
  BUF U220 ( .I(n29541), .Z(n29350) );
  BUF U221 ( .I(n29541), .Z(n29351) );
  BUF U222 ( .I(n29541), .Z(n29352) );
  BUF U223 ( .I(n29540), .Z(n29353) );
  BUF U224 ( .I(n29540), .Z(n29354) );
  BUF U225 ( .I(n29537), .Z(n29364) );
  BUF U226 ( .I(n29504), .Z(n29461) );
  BUF U227 ( .I(n29504), .Z(n29462) );
  BUF U228 ( .I(n29504), .Z(n29463) );
  BUF U229 ( .I(n29503), .Z(n29464) );
  BUF U230 ( .I(n29503), .Z(n29465) );
  BUF U231 ( .I(n29503), .Z(n29466) );
  BUF U232 ( .I(n29502), .Z(n29467) );
  BUF U233 ( .I(n29502), .Z(n29468) );
  BUF U234 ( .I(n29502), .Z(n29469) );
  BUF U235 ( .I(n29501), .Z(n29470) );
  BUF U236 ( .I(n29508), .Z(n29451) );
  BUF U237 ( .I(n29507), .Z(n29452) );
  BUF U238 ( .I(n29507), .Z(n29453) );
  BUF U239 ( .I(n29507), .Z(n29454) );
  BUF U240 ( .I(n29506), .Z(n29455) );
  BUF U241 ( .I(n29506), .Z(n29456) );
  BUF U242 ( .I(n29506), .Z(n29457) );
  BUF U243 ( .I(n29505), .Z(n29458) );
  BUF U244 ( .I(n29505), .Z(n29459) );
  BUF U245 ( .I(n29505), .Z(n29460) );
  BUF U246 ( .I(n29501), .Z(n29471) );
  BUF U247 ( .I(n29501), .Z(n29472) );
  BUF U248 ( .I(n29518), .Z(n29419) );
  BUF U249 ( .I(n29518), .Z(n29420) );
  BUF U250 ( .I(n29518), .Z(n29421) );
  BUF U251 ( .I(n29517), .Z(n29422) );
  BUF U252 ( .I(n29517), .Z(n29423) );
  BUF U253 ( .I(n29517), .Z(n29424) );
  BUF U254 ( .I(n29516), .Z(n29425) );
  BUF U255 ( .I(n29516), .Z(n29426) );
  BUF U256 ( .I(n29516), .Z(n29427) );
  BUF U257 ( .I(n29522), .Z(n29407) );
  BUF U258 ( .I(n29522), .Z(n29408) );
  BUF U259 ( .I(n29522), .Z(n29409) );
  BUF U260 ( .I(n29521), .Z(n29410) );
  BUF U261 ( .I(n29521), .Z(n29411) );
  BUF U262 ( .I(n29521), .Z(n29412) );
  BUF U263 ( .I(n29520), .Z(n29413) );
  BUF U264 ( .I(n29520), .Z(n29414) );
  BUF U265 ( .I(n29520), .Z(n29415) );
  BUF U266 ( .I(n29519), .Z(n29416) );
  BUF U267 ( .I(n29519), .Z(n29417) );
  BUF U268 ( .I(n29519), .Z(n29418) );
  BUF U269 ( .I(n29511), .Z(n29440) );
  BUF U270 ( .I(n29511), .Z(n29441) );
  BUF U271 ( .I(n29511), .Z(n29442) );
  BUF U272 ( .I(n29510), .Z(n29443) );
  BUF U273 ( .I(n29510), .Z(n29444) );
  BUF U274 ( .I(n29510), .Z(n29445) );
  BUF U275 ( .I(n29509), .Z(n29446) );
  BUF U276 ( .I(n29509), .Z(n29447) );
  BUF U277 ( .I(n29509), .Z(n29448) );
  BUF U278 ( .I(n29508), .Z(n29449) );
  BUF U279 ( .I(n29508), .Z(n29450) );
  BUF U280 ( .I(n29515), .Z(n29428) );
  BUF U281 ( .I(n29515), .Z(n29429) );
  BUF U282 ( .I(n29515), .Z(n29430) );
  BUF U283 ( .I(n29514), .Z(n29431) );
  BUF U284 ( .I(n29514), .Z(n29432) );
  BUF U285 ( .I(n29514), .Z(n29433) );
  BUF U286 ( .I(n29513), .Z(n29434) );
  BUF U287 ( .I(n29513), .Z(n29435) );
  BUF U288 ( .I(n29513), .Z(n29436) );
  BUF U289 ( .I(n29512), .Z(n29437) );
  BUF U290 ( .I(n29512), .Z(n29438) );
  BUF U291 ( .I(n29512), .Z(n29439) );
  BUF U292 ( .I(n26994), .Z(n27111) );
  BUF U293 ( .I(n26994), .Z(n27110) );
  BUF U294 ( .I(n26995), .Z(n27109) );
  BUF U295 ( .I(n26995), .Z(n27108) );
  BUF U296 ( .I(n26995), .Z(n27107) );
  BUF U297 ( .I(n26996), .Z(n27106) );
  BUF U298 ( .I(n26996), .Z(n27105) );
  BUF U299 ( .I(n26996), .Z(n27104) );
  BUF U300 ( .I(n26997), .Z(n27103) );
  BUF U301 ( .I(n26981), .Z(n27150) );
  BUF U302 ( .I(n26982), .Z(n27147) );
  BUF U303 ( .I(n26981), .Z(n27149) );
  BUF U304 ( .I(n26982), .Z(n27148) );
  BUF U305 ( .I(n26982), .Z(n27146) );
  BUF U306 ( .I(n26983), .Z(n27145) );
  BUF U307 ( .I(n26983), .Z(n27144) );
  BUF U308 ( .I(n26983), .Z(n27143) );
  BUF U309 ( .I(n26968), .Z(n27189) );
  BUF U310 ( .I(n26968), .Z(n27190) );
  BUF U311 ( .I(n26968), .Z(n27188) );
  BUF U312 ( .I(n26969), .Z(n27187) );
  BUF U313 ( .I(n26970), .Z(n27184) );
  BUF U314 ( .I(n26969), .Z(n27186) );
  BUF U315 ( .I(n26969), .Z(n27185) );
  BUF U316 ( .I(n26970), .Z(n27183) );
  BUF U317 ( .I(n26970), .Z(n27182) );
  BUF U318 ( .I(n26955), .Z(n27229) );
  BUF U319 ( .I(n26956), .Z(n27226) );
  BUF U320 ( .I(n26955), .Z(n27228) );
  BUF U321 ( .I(n26955), .Z(n27227) );
  BUF U322 ( .I(n26956), .Z(n27225) );
  BUF U323 ( .I(n26956), .Z(n27224) );
  BUF U324 ( .I(n26957), .Z(n27221) );
  BUF U325 ( .I(n26957), .Z(n27223) );
  BUF U326 ( .I(n26957), .Z(n27222) );
  BUF U327 ( .I(n26941), .Z(n27269) );
  BUF U328 ( .I(n26942), .Z(n27268) );
  BUF U329 ( .I(n26942), .Z(n27267) );
  BUF U330 ( .I(n26942), .Z(n27266) );
  BUF U331 ( .I(n26943), .Z(n27265) );
  BUF U332 ( .I(n26943), .Z(n27263) );
  BUF U333 ( .I(n26943), .Z(n27264) );
  BUF U334 ( .I(n26944), .Z(n27262) );
  BUF U335 ( .I(n26944), .Z(n27261) );
  BUF U336 ( .I(n26929), .Z(n27307) );
  BUF U337 ( .I(n26928), .Z(n27308) );
  BUF U338 ( .I(n26929), .Z(n27306) );
  BUF U339 ( .I(n26929), .Z(n27305) );
  BUF U340 ( .I(n26930), .Z(n27304) );
  BUF U341 ( .I(n26930), .Z(n27303) );
  BUF U342 ( .I(n26930), .Z(n27302) );
  BUF U343 ( .I(n26931), .Z(n27301) );
  BUF U344 ( .I(n26931), .Z(n27300) );
  BUF U345 ( .I(n26997), .Z(n27102) );
  BUF U346 ( .I(n26997), .Z(n27101) );
  BUF U347 ( .I(n26998), .Z(n27100) );
  BUF U348 ( .I(n26998), .Z(n27099) );
  BUF U349 ( .I(n26998), .Z(n27098) );
  BUF U350 ( .I(n26984), .Z(n27142) );
  BUF U351 ( .I(n26984), .Z(n27141) );
  BUF U352 ( .I(n26984), .Z(n27140) );
  BUF U353 ( .I(n26985), .Z(n27139) );
  BUF U354 ( .I(n26985), .Z(n27138) );
  BUF U355 ( .I(n26985), .Z(n27137) );
  BUF U356 ( .I(n26986), .Z(n27136) );
  BUF U357 ( .I(n26986), .Z(n27135) );
  BUF U358 ( .I(n26986), .Z(n27134) );
  BUF U359 ( .I(n26987), .Z(n27133) );
  BUF U360 ( .I(n26991), .Z(n27120) );
  BUF U361 ( .I(n26991), .Z(n27121) );
  BUF U362 ( .I(n26991), .Z(n27119) );
  BUF U363 ( .I(n26992), .Z(n27118) );
  BUF U364 ( .I(n26993), .Z(n27115) );
  BUF U365 ( .I(n26992), .Z(n27117) );
  BUF U366 ( .I(n26992), .Z(n27116) );
  BUF U367 ( .I(n26994), .Z(n27112) );
  BUF U368 ( .I(n26993), .Z(n27114) );
  BUF U369 ( .I(n26993), .Z(n27113) );
  BUF U370 ( .I(n26988), .Z(n27130) );
  BUF U371 ( .I(n26987), .Z(n27132) );
  BUF U372 ( .I(n26987), .Z(n27131) );
  BUF U373 ( .I(n26988), .Z(n27129) );
  BUF U374 ( .I(n26988), .Z(n27128) );
  BUF U375 ( .I(n26989), .Z(n27125) );
  BUF U376 ( .I(n26989), .Z(n27127) );
  BUF U377 ( .I(n26989), .Z(n27126) );
  BUF U378 ( .I(n26990), .Z(n27122) );
  BUF U379 ( .I(n26990), .Z(n27124) );
  BUF U380 ( .I(n26990), .Z(n27123) );
  BUF U381 ( .I(n26971), .Z(n27179) );
  BUF U382 ( .I(n26971), .Z(n27181) );
  BUF U383 ( .I(n26971), .Z(n27180) );
  BUF U384 ( .I(n26972), .Z(n27178) );
  BUF U385 ( .I(n26972), .Z(n27177) );
  BUF U386 ( .I(n26972), .Z(n27176) );
  BUF U387 ( .I(n26973), .Z(n27175) );
  BUF U388 ( .I(n26973), .Z(n27174) );
  BUF U389 ( .I(n26973), .Z(n27173) );
  BUF U390 ( .I(n26974), .Z(n27172) );
  BUF U391 ( .I(n26978), .Z(n27160) );
  BUF U392 ( .I(n26979), .Z(n27157) );
  BUF U393 ( .I(n26978), .Z(n27159) );
  BUF U394 ( .I(n26978), .Z(n27158) );
  BUF U395 ( .I(n26979), .Z(n27156) );
  BUF U396 ( .I(n26979), .Z(n27155) );
  BUF U397 ( .I(n26981), .Z(n27151) );
  BUF U398 ( .I(n26980), .Z(n27152) );
  BUF U399 ( .I(n26980), .Z(n27154) );
  BUF U400 ( .I(n26980), .Z(n27153) );
  BUF U401 ( .I(n26974), .Z(n27171) );
  BUF U402 ( .I(n26974), .Z(n27170) );
  BUF U403 ( .I(n26975), .Z(n27169) );
  BUF U404 ( .I(n26975), .Z(n27167) );
  BUF U405 ( .I(n26975), .Z(n27168) );
  BUF U406 ( .I(n26976), .Z(n27166) );
  BUF U407 ( .I(n26976), .Z(n27165) );
  BUF U408 ( .I(n26977), .Z(n27162) );
  BUF U409 ( .I(n26977), .Z(n27161) );
  BUF U410 ( .I(n26976), .Z(n27164) );
  BUF U411 ( .I(n26977), .Z(n27163) );
  BUF U412 ( .I(n26958), .Z(n27220) );
  BUF U413 ( .I(n26958), .Z(n27219) );
  BUF U414 ( .I(n26958), .Z(n27218) );
  BUF U415 ( .I(n26959), .Z(n27217) );
  BUF U416 ( .I(n26959), .Z(n27216) );
  BUF U417 ( .I(n26959), .Z(n27215) );
  BUF U418 ( .I(n26960), .Z(n27214) );
  BUF U419 ( .I(n26960), .Z(n27213) );
  BUF U420 ( .I(n26960), .Z(n27212) );
  BUF U421 ( .I(n26961), .Z(n27211) );
  BUF U422 ( .I(n26965), .Z(n27199) );
  BUF U423 ( .I(n26964), .Z(n27200) );
  BUF U424 ( .I(n26965), .Z(n27198) );
  BUF U425 ( .I(n26965), .Z(n27197) );
  BUF U426 ( .I(n26966), .Z(n27194) );
  BUF U427 ( .I(n26966), .Z(n27196) );
  BUF U428 ( .I(n26966), .Z(n27195) );
  BUF U429 ( .I(n26967), .Z(n27191) );
  BUF U430 ( .I(n26967), .Z(n27193) );
  BUF U431 ( .I(n26967), .Z(n27192) );
  BUF U432 ( .I(n26961), .Z(n27210) );
  BUF U433 ( .I(n26961), .Z(n27209) );
  BUF U434 ( .I(n26962), .Z(n27208) );
  BUF U435 ( .I(n26962), .Z(n27207) );
  BUF U436 ( .I(n26962), .Z(n27206) );
  BUF U437 ( .I(n26963), .Z(n27205) );
  BUF U438 ( .I(n26963), .Z(n27204) );
  BUF U439 ( .I(n26964), .Z(n27201) );
  BUF U440 ( .I(n26963), .Z(n27203) );
  BUF U441 ( .I(n26964), .Z(n27202) );
  BUF U442 ( .I(n26945), .Z(n27258) );
  BUF U443 ( .I(n26944), .Z(n27260) );
  BUF U444 ( .I(n26945), .Z(n27259) );
  BUF U445 ( .I(n26945), .Z(n27257) );
  BUF U446 ( .I(n26946), .Z(n27256) );
  BUF U447 ( .I(n26947), .Z(n27253) );
  BUF U448 ( .I(n26946), .Z(n27255) );
  BUF U449 ( .I(n26946), .Z(n27254) );
  BUF U450 ( .I(n26947), .Z(n27252) );
  BUF U451 ( .I(n26947), .Z(n27251) );
  BUF U452 ( .I(n26951), .Z(n27239) );
  BUF U453 ( .I(n26952), .Z(n27238) );
  BUF U454 ( .I(n26952), .Z(n27237) );
  BUF U455 ( .I(n26952), .Z(n27236) );
  BUF U456 ( .I(n26953), .Z(n27235) );
  BUF U457 ( .I(n26953), .Z(n27234) );
  BUF U458 ( .I(n26954), .Z(n27230) );
  BUF U459 ( .I(n26953), .Z(n27233) );
  BUF U460 ( .I(n26954), .Z(n27231) );
  BUF U461 ( .I(n26954), .Z(n27232) );
  BUF U462 ( .I(n26948), .Z(n27248) );
  BUF U463 ( .I(n26948), .Z(n27250) );
  BUF U464 ( .I(n26948), .Z(n27249) );
  BUF U465 ( .I(n26949), .Z(n27247) );
  BUF U466 ( .I(n26949), .Z(n27246) );
  BUF U467 ( .I(n26950), .Z(n27243) );
  BUF U468 ( .I(n26949), .Z(n27245) );
  BUF U469 ( .I(n26950), .Z(n27244) );
  BUF U470 ( .I(n26951), .Z(n27240) );
  BUF U471 ( .I(n26950), .Z(n27242) );
  BUF U472 ( .I(n26951), .Z(n27241) );
  BUF U473 ( .I(n26931), .Z(n27299) );
  BUF U474 ( .I(n26932), .Z(n27298) );
  BUF U475 ( .I(n26932), .Z(n27297) );
  BUF U476 ( .I(n26932), .Z(n27296) );
  BUF U477 ( .I(n26933), .Z(n27295) );
  BUF U478 ( .I(n26933), .Z(n27294) );
  BUF U479 ( .I(n26933), .Z(n27293) );
  BUF U480 ( .I(n26934), .Z(n27292) );
  BUF U481 ( .I(n26934), .Z(n27291) );
  BUF U482 ( .I(n26934), .Z(n27290) );
  BUF U483 ( .I(n26938), .Z(n27278) );
  BUF U484 ( .I(n26939), .Z(n27275) );
  BUF U485 ( .I(n26939), .Z(n27277) );
  BUF U486 ( .I(n26939), .Z(n27276) );
  BUF U487 ( .I(n26940), .Z(n27274) );
  BUF U488 ( .I(n26940), .Z(n27273) );
  BUF U489 ( .I(n26941), .Z(n27270) );
  BUF U490 ( .I(n26940), .Z(n27272) );
  BUF U491 ( .I(n26941), .Z(n27271) );
  BUF U492 ( .I(n26935), .Z(n27289) );
  BUF U493 ( .I(n26935), .Z(n27288) );
  BUF U494 ( .I(n26936), .Z(n27285) );
  BUF U495 ( .I(n26935), .Z(n27287) );
  BUF U496 ( .I(n26936), .Z(n27286) );
  BUF U497 ( .I(n26936), .Z(n27284) );
  BUF U498 ( .I(n26937), .Z(n27283) );
  BUF U499 ( .I(n26938), .Z(n27279) );
  BUF U500 ( .I(n26938), .Z(n27280) );
  BUF U501 ( .I(n26937), .Z(n27282) );
  BUF U502 ( .I(n26937), .Z(n27281) );
  BUF U503 ( .I(n26919), .Z(n27337) );
  BUF U504 ( .I(n26919), .Z(n27336) );
  BUF U505 ( .I(n26919), .Z(n27335) );
  BUF U506 ( .I(n26920), .Z(n27334) );
  BUF U507 ( .I(n26920), .Z(n27333) );
  BUF U508 ( .I(n26920), .Z(n27332) );
  BUF U509 ( .I(n26921), .Z(n27331) );
  BUF U510 ( .I(n26921), .Z(n27330) );
  BUF U511 ( .I(n26925), .Z(n27317) );
  BUF U512 ( .I(n26925), .Z(n27318) );
  BUF U513 ( .I(n26926), .Z(n27316) );
  BUF U514 ( .I(n26926), .Z(n27315) );
  BUF U515 ( .I(n26927), .Z(n27312) );
  BUF U516 ( .I(n26926), .Z(n27314) );
  BUF U517 ( .I(n26927), .Z(n27313) );
  BUF U518 ( .I(n26928), .Z(n27309) );
  BUF U519 ( .I(n26927), .Z(n27311) );
  BUF U520 ( .I(n26928), .Z(n27310) );
  BUF U521 ( .I(n26921), .Z(n27329) );
  BUF U522 ( .I(n26922), .Z(n27327) );
  BUF U523 ( .I(n26922), .Z(n27328) );
  BUF U524 ( .I(n26922), .Z(n27326) );
  BUF U525 ( .I(n26923), .Z(n27325) );
  BUF U526 ( .I(n26924), .Z(n27322) );
  BUF U527 ( .I(n26923), .Z(n27324) );
  BUF U528 ( .I(n26923), .Z(n27323) );
  BUF U529 ( .I(n26925), .Z(n27319) );
  BUF U530 ( .I(n26924), .Z(n27321) );
  BUF U531 ( .I(n26924), .Z(n27320) );
  BUF U532 ( .I(n26519), .Z(n26635) );
  BUF U533 ( .I(n26506), .Z(n26675) );
  BUF U534 ( .I(n26493), .Z(n26714) );
  BUF U535 ( .I(n26480), .Z(n26754) );
  BUF U536 ( .I(n26467), .Z(n26793) );
  BUF U537 ( .I(n26454), .Z(n26832) );
  BUF U538 ( .I(n26522), .Z(n26626) );
  BUF U539 ( .I(n26509), .Z(n26665) );
  BUF U540 ( .I(n26511), .Z(n26660) );
  BUF U541 ( .I(n26516), .Z(n26645) );
  BUF U542 ( .I(n26496), .Z(n26704) );
  BUF U543 ( .I(n26496), .Z(n26705) );
  BUF U544 ( .I(n26498), .Z(n26699) );
  BUF U545 ( .I(n26503), .Z(n26685) );
  BUF U546 ( .I(n26483), .Z(n26744) );
  BUF U547 ( .I(n26485), .Z(n26739) );
  BUF U548 ( .I(n26490), .Z(n26724) );
  BUF U549 ( .I(n26470), .Z(n26783) );
  BUF U550 ( .I(n26472), .Z(n26778) );
  BUF U551 ( .I(n26477), .Z(n26763) );
  BUF U552 ( .I(n26457), .Z(n26823) );
  BUF U553 ( .I(n26457), .Z(n26822) );
  BUF U554 ( .I(n26458), .Z(n26818) );
  BUF U555 ( .I(n26463), .Z(n26803) );
  BUF U556 ( .I(n26444), .Z(n26862) );
  BUF U557 ( .I(n26445), .Z(n26857) );
  BUF U558 ( .I(n26450), .Z(n26842) );
  BUF U559 ( .I(n26519), .Z(n26636) );
  BUF U560 ( .I(n26520), .Z(n26634) );
  BUF U561 ( .I(n26520), .Z(n26633) );
  BUF U562 ( .I(n26520), .Z(n26632) );
  BUF U563 ( .I(n26521), .Z(n26631) );
  BUF U564 ( .I(n26521), .Z(n26630) );
  BUF U565 ( .I(n26521), .Z(n26629) );
  BUF U566 ( .I(n26522), .Z(n26628) );
  BUF U567 ( .I(n26507), .Z(n26672) );
  BUF U568 ( .I(n26506), .Z(n26674) );
  BUF U569 ( .I(n26507), .Z(n26673) );
  BUF U570 ( .I(n26507), .Z(n26671) );
  BUF U571 ( .I(n26508), .Z(n26670) );
  BUF U572 ( .I(n26508), .Z(n26669) );
  BUF U573 ( .I(n26508), .Z(n26668) );
  BUF U574 ( .I(n26493), .Z(n26715) );
  BUF U575 ( .I(n26493), .Z(n26713) );
  BUF U576 ( .I(n26494), .Z(n26712) );
  BUF U577 ( .I(n26495), .Z(n26709) );
  BUF U578 ( .I(n26494), .Z(n26711) );
  BUF U579 ( .I(n26494), .Z(n26710) );
  BUF U580 ( .I(n26495), .Z(n26708) );
  BUF U581 ( .I(n26495), .Z(n26707) );
  BUF U582 ( .I(n26481), .Z(n26751) );
  BUF U583 ( .I(n26480), .Z(n26753) );
  BUF U584 ( .I(n26480), .Z(n26752) );
  BUF U585 ( .I(n26481), .Z(n26750) );
  BUF U586 ( .I(n26481), .Z(n26749) );
  BUF U587 ( .I(n26482), .Z(n26746) );
  BUF U588 ( .I(n26482), .Z(n26748) );
  BUF U589 ( .I(n26482), .Z(n26747) );
  BUF U590 ( .I(n26466), .Z(n26794) );
  BUF U591 ( .I(n26467), .Z(n26792) );
  BUF U592 ( .I(n26467), .Z(n26791) );
  BUF U593 ( .I(n26468), .Z(n26790) );
  BUF U594 ( .I(n26468), .Z(n26788) );
  BUF U595 ( .I(n26468), .Z(n26789) );
  BUF U596 ( .I(n26469), .Z(n26787) );
  BUF U597 ( .I(n26469), .Z(n26786) );
  BUF U598 ( .I(n26453), .Z(n26833) );
  BUF U599 ( .I(n26454), .Z(n26831) );
  BUF U600 ( .I(n26454), .Z(n26830) );
  BUF U601 ( .I(n26455), .Z(n26829) );
  BUF U602 ( .I(n26455), .Z(n26828) );
  BUF U603 ( .I(n26455), .Z(n26827) );
  BUF U604 ( .I(n26456), .Z(n26826) );
  BUF U605 ( .I(n26456), .Z(n26825) );
  BUF U606 ( .I(n26522), .Z(n26627) );
  BUF U607 ( .I(n26523), .Z(n26625) );
  BUF U608 ( .I(n26523), .Z(n26624) );
  BUF U609 ( .I(n26523), .Z(n26623) );
  BUF U610 ( .I(n26509), .Z(n26667) );
  BUF U611 ( .I(n26509), .Z(n26666) );
  BUF U612 ( .I(n26510), .Z(n26664) );
  BUF U613 ( .I(n26510), .Z(n26663) );
  BUF U614 ( .I(n26510), .Z(n26662) );
  BUF U615 ( .I(n26511), .Z(n26661) );
  BUF U616 ( .I(n26511), .Z(n26659) );
  BUF U617 ( .I(n26512), .Z(n26658) );
  BUF U618 ( .I(n26516), .Z(n26646) );
  BUF U619 ( .I(n26516), .Z(n26644) );
  BUF U620 ( .I(n26517), .Z(n26643) );
  BUF U621 ( .I(n26518), .Z(n26640) );
  BUF U622 ( .I(n26517), .Z(n26642) );
  BUF U623 ( .I(n26517), .Z(n26641) );
  BUF U624 ( .I(n26519), .Z(n26637) );
  BUF U625 ( .I(n26518), .Z(n26639) );
  BUF U626 ( .I(n26518), .Z(n26638) );
  BUF U627 ( .I(n26513), .Z(n26655) );
  BUF U628 ( .I(n26512), .Z(n26657) );
  BUF U629 ( .I(n26512), .Z(n26656) );
  BUF U630 ( .I(n26513), .Z(n26654) );
  BUF U631 ( .I(n26513), .Z(n26653) );
  BUF U632 ( .I(n26514), .Z(n26650) );
  BUF U633 ( .I(n26514), .Z(n26652) );
  BUF U634 ( .I(n26514), .Z(n26651) );
  BUF U635 ( .I(n26515), .Z(n26647) );
  BUF U636 ( .I(n26515), .Z(n26649) );
  BUF U637 ( .I(n26515), .Z(n26648) );
  BUF U638 ( .I(n26496), .Z(n26706) );
  BUF U639 ( .I(n26497), .Z(n26703) );
  BUF U640 ( .I(n26497), .Z(n26702) );
  BUF U641 ( .I(n26497), .Z(n26701) );
  BUF U642 ( .I(n26498), .Z(n26700) );
  BUF U643 ( .I(n26498), .Z(n26698) );
  BUF U644 ( .I(n26499), .Z(n26697) );
  BUF U645 ( .I(n26504), .Z(n26682) );
  BUF U646 ( .I(n26503), .Z(n26684) );
  BUF U647 ( .I(n26503), .Z(n26683) );
  BUF U648 ( .I(n26504), .Z(n26681) );
  BUF U649 ( .I(n26504), .Z(n26680) );
  BUF U650 ( .I(n26506), .Z(n26676) );
  BUF U651 ( .I(n26505), .Z(n26677) );
  BUF U652 ( .I(n26505), .Z(n26679) );
  BUF U653 ( .I(n26505), .Z(n26678) );
  BUF U654 ( .I(n26499), .Z(n26696) );
  BUF U655 ( .I(n26499), .Z(n26695) );
  BUF U656 ( .I(n26500), .Z(n26694) );
  BUF U657 ( .I(n26500), .Z(n26692) );
  BUF U658 ( .I(n26500), .Z(n26693) );
  BUF U659 ( .I(n26501), .Z(n26691) );
  BUF U660 ( .I(n26501), .Z(n26690) );
  BUF U661 ( .I(n26502), .Z(n26687) );
  BUF U662 ( .I(n26502), .Z(n26686) );
  BUF U663 ( .I(n26501), .Z(n26689) );
  BUF U664 ( .I(n26502), .Z(n26688) );
  BUF U665 ( .I(n26483), .Z(n26745) );
  BUF U666 ( .I(n26483), .Z(n26743) );
  BUF U667 ( .I(n26484), .Z(n26742) );
  BUF U668 ( .I(n26484), .Z(n26741) );
  BUF U669 ( .I(n26484), .Z(n26740) );
  BUF U670 ( .I(n26485), .Z(n26738) );
  BUF U671 ( .I(n26485), .Z(n26737) );
  BUF U672 ( .I(n26486), .Z(n26736) );
  BUF U673 ( .I(n26489), .Z(n26725) );
  BUF U674 ( .I(n26490), .Z(n26723) );
  BUF U675 ( .I(n26490), .Z(n26722) );
  BUF U676 ( .I(n26491), .Z(n26719) );
  BUF U677 ( .I(n26491), .Z(n26721) );
  BUF U678 ( .I(n26491), .Z(n26720) );
  BUF U679 ( .I(n26492), .Z(n26716) );
  BUF U680 ( .I(n26492), .Z(n26718) );
  BUF U681 ( .I(n26492), .Z(n26717) );
  BUF U682 ( .I(n26486), .Z(n26735) );
  BUF U683 ( .I(n26486), .Z(n26734) );
  BUF U684 ( .I(n26487), .Z(n26733) );
  BUF U685 ( .I(n26487), .Z(n26732) );
  BUF U686 ( .I(n26487), .Z(n26731) );
  BUF U687 ( .I(n26488), .Z(n26730) );
  BUF U688 ( .I(n26488), .Z(n26729) );
  BUF U689 ( .I(n26489), .Z(n26726) );
  BUF U690 ( .I(n26488), .Z(n26728) );
  BUF U691 ( .I(n26489), .Z(n26727) );
  BUF U692 ( .I(n26469), .Z(n26785) );
  BUF U693 ( .I(n26470), .Z(n26784) );
  BUF U694 ( .I(n26470), .Z(n26782) );
  BUF U695 ( .I(n26471), .Z(n26781) );
  BUF U696 ( .I(n26471), .Z(n26780) );
  BUF U697 ( .I(n26471), .Z(n26779) );
  BUF U698 ( .I(n26472), .Z(n26777) );
  BUF U699 ( .I(n26472), .Z(n26776) );
  BUF U700 ( .I(n26476), .Z(n26764) );
  BUF U701 ( .I(n26477), .Z(n26762) );
  BUF U702 ( .I(n26477), .Z(n26761) );
  BUF U703 ( .I(n26478), .Z(n26760) );
  BUF U704 ( .I(n26478), .Z(n26759) );
  BUF U705 ( .I(n26479), .Z(n26755) );
  BUF U706 ( .I(n26478), .Z(n26758) );
  BUF U707 ( .I(n26479), .Z(n26756) );
  BUF U708 ( .I(n26479), .Z(n26757) );
  BUF U709 ( .I(n26473), .Z(n26773) );
  BUF U710 ( .I(n26473), .Z(n26775) );
  BUF U711 ( .I(n26473), .Z(n26774) );
  BUF U712 ( .I(n26474), .Z(n26772) );
  BUF U713 ( .I(n26474), .Z(n26771) );
  BUF U714 ( .I(n26475), .Z(n26768) );
  BUF U715 ( .I(n26474), .Z(n26770) );
  BUF U716 ( .I(n26475), .Z(n26769) );
  BUF U717 ( .I(n26476), .Z(n26765) );
  BUF U718 ( .I(n26475), .Z(n26767) );
  BUF U719 ( .I(n26476), .Z(n26766) );
  BUF U720 ( .I(n26456), .Z(n26824) );
  BUF U721 ( .I(n26457), .Z(n26821) );
  BUF U722 ( .I(n26458), .Z(n26820) );
  BUF U723 ( .I(n26458), .Z(n26819) );
  BUF U724 ( .I(n26459), .Z(n26817) );
  BUF U725 ( .I(n26459), .Z(n26816) );
  BUF U726 ( .I(n26459), .Z(n26815) );
  BUF U727 ( .I(n26464), .Z(n26800) );
  BUF U728 ( .I(n26464), .Z(n26802) );
  BUF U729 ( .I(n26464), .Z(n26801) );
  BUF U730 ( .I(n26465), .Z(n26799) );
  BUF U731 ( .I(n26465), .Z(n26798) );
  BUF U732 ( .I(n26466), .Z(n26795) );
  BUF U733 ( .I(n26465), .Z(n26797) );
  BUF U734 ( .I(n26466), .Z(n26796) );
  BUF U735 ( .I(n26460), .Z(n26814) );
  BUF U736 ( .I(n26460), .Z(n26813) );
  BUF U737 ( .I(n26461), .Z(n26810) );
  BUF U738 ( .I(n26460), .Z(n26812) );
  BUF U739 ( .I(n26461), .Z(n26811) );
  BUF U740 ( .I(n26461), .Z(n26809) );
  BUF U741 ( .I(n26462), .Z(n26808) );
  BUF U742 ( .I(n26463), .Z(n26804) );
  BUF U743 ( .I(n26463), .Z(n26805) );
  BUF U744 ( .I(n26462), .Z(n26807) );
  BUF U745 ( .I(n26462), .Z(n26806) );
  BUF U746 ( .I(n26444), .Z(n26861) );
  BUF U747 ( .I(n26444), .Z(n26860) );
  BUF U748 ( .I(n26445), .Z(n26859) );
  BUF U749 ( .I(n26445), .Z(n26858) );
  BUF U750 ( .I(n26446), .Z(n26856) );
  BUF U751 ( .I(n26446), .Z(n26855) );
  BUF U752 ( .I(n26450), .Z(n26843) );
  BUF U753 ( .I(n26451), .Z(n26841) );
  BUF U754 ( .I(n26451), .Z(n26840) );
  BUF U755 ( .I(n26452), .Z(n26837) );
  BUF U756 ( .I(n26451), .Z(n26839) );
  BUF U757 ( .I(n26452), .Z(n26838) );
  BUF U758 ( .I(n26453), .Z(n26834) );
  BUF U759 ( .I(n26452), .Z(n26836) );
  BUF U760 ( .I(n26453), .Z(n26835) );
  BUF U761 ( .I(n26446), .Z(n26854) );
  BUF U762 ( .I(n26447), .Z(n26852) );
  BUF U763 ( .I(n26447), .Z(n26853) );
  BUF U764 ( .I(n26447), .Z(n26851) );
  BUF U765 ( .I(n26448), .Z(n26850) );
  BUF U766 ( .I(n26449), .Z(n26847) );
  BUF U767 ( .I(n26448), .Z(n26849) );
  BUF U768 ( .I(n26448), .Z(n26848) );
  BUF U769 ( .I(n26450), .Z(n26844) );
  BUF U770 ( .I(n26449), .Z(n26846) );
  BUF U771 ( .I(n26449), .Z(n26845) );
  I_NAND2 U772 ( .A1(n25), .B1(n29322), .ZN(n26) );
  I_NAND2 U773 ( .A1(n28), .B1(n29386), .ZN(n29) );
  I_NAND2 U774 ( .A1(n31), .B1(n29380), .ZN(n32) );
  I_NAND2 U775 ( .A1(n34), .B1(n29375), .ZN(n35) );
  I_NAND2 U776 ( .A1(n37), .B1(n29375), .ZN(n38) );
  I_NAND2 U777 ( .A1(n40), .B1(n29375), .ZN(n41) );
  I_NAND2 U778 ( .A1(n43), .B1(n29375), .ZN(n44) );
  I_NAND2 U779 ( .A1(n46), .B1(n29375), .ZN(n47) );
  I_NAND2 U780 ( .A1(n49), .B1(n29375), .ZN(n50) );
  I_NAND2 U781 ( .A1(n52), .B1(n29376), .ZN(n53) );
  I_NAND2 U782 ( .A1(n55), .B1(n29376), .ZN(n56) );
  I_NAND2 U783 ( .A1(n58), .B1(n29376), .ZN(n59) );
  I_NAND2 U784 ( .A1(n61), .B1(n29376), .ZN(n62) );
  I_NAND2 U785 ( .A1(n64), .B1(n29376), .ZN(n65) );
  I_NAND2 U786 ( .A1(n67), .B1(n29376), .ZN(n68) );
  I_NAND2 U787 ( .A1(n70), .B1(n29376), .ZN(n71) );
  I_NAND2 U788 ( .A1(n73), .B1(n29376), .ZN(n74) );
  I_NAND2 U789 ( .A1(n76), .B1(n29376), .ZN(n77) );
  I_NAND2 U790 ( .A1(n79), .B1(n29376), .ZN(n80) );
  I_NAND2 U791 ( .A1(n82), .B1(n29376), .ZN(n83) );
  I_NAND2 U792 ( .A1(n85), .B1(n29376), .ZN(n86) );
  I_NAND2 U793 ( .A1(n88), .B1(n29377), .ZN(n89) );
  I_NAND2 U794 ( .A1(n91), .B1(n29377), .ZN(n92) );
  I_NAND2 U795 ( .A1(n94), .B1(n29377), .ZN(n95) );
  I_NAND2 U796 ( .A1(n97), .B1(n29377), .ZN(n98) );
  I_NAND2 U797 ( .A1(n100), .B1(n29377), .ZN(n101) );
  I_NAND2 U798 ( .A1(n103), .B1(n29377), .ZN(n104) );
  I_NAND2 U799 ( .A1(n106), .B1(n29377), .ZN(n107) );
  I_NAND2 U800 ( .A1(n109), .B1(n29377), .ZN(n110) );
  I_NAND2 U801 ( .A1(n112), .B1(n29377), .ZN(n113) );
  I_NAND2 U802 ( .A1(n115), .B1(n29377), .ZN(n116) );
  I_NAND2 U803 ( .A1(n118), .B1(n29377), .ZN(n119) );
  I_NAND2 U804 ( .A1(n121), .B1(n29377), .ZN(n122) );
  I_NAND2 U805 ( .A1(n124), .B1(n29378), .ZN(n125) );
  I_NAND2 U806 ( .A1(n127), .B1(n29378), .ZN(n128) );
  I_NAND2 U807 ( .A1(n130), .B1(n29378), .ZN(n131) );
  I_NAND2 U808 ( .A1(n133), .B1(n29378), .ZN(n134) );
  I_NAND2 U809 ( .A1(n136), .B1(n29378), .ZN(n137) );
  I_NAND2 U810 ( .A1(n139), .B1(n29378), .ZN(n140) );
  I_NAND2 U811 ( .A1(n142), .B1(n29378), .ZN(n143) );
  I_NAND2 U812 ( .A1(n145), .B1(n29378), .ZN(n146) );
  I_NAND2 U813 ( .A1(n148), .B1(n29378), .ZN(n149) );
  I_NAND2 U814 ( .A1(n151), .B1(n29378), .ZN(n152) );
  I_NAND2 U815 ( .A1(n154), .B1(n29378), .ZN(n155) );
  I_NAND2 U816 ( .A1(n157), .B1(n29378), .ZN(n158) );
  I_NAND2 U817 ( .A1(n160), .B1(n29379), .ZN(n161) );
  I_NAND2 U818 ( .A1(n163), .B1(n29379), .ZN(n164) );
  I_NAND2 U819 ( .A1(n166), .B1(n29379), .ZN(n167) );
  I_NAND2 U820 ( .A1(n169), .B1(n29379), .ZN(n170) );
  I_NAND2 U821 ( .A1(n172), .B1(n29379), .ZN(n173) );
  I_NAND2 U822 ( .A1(n175), .B1(n29379), .ZN(n176) );
  I_NAND2 U823 ( .A1(n178), .B1(n29379), .ZN(n179) );
  I_NAND2 U824 ( .A1(n181), .B1(n29379), .ZN(n182) );
  I_NAND2 U825 ( .A1(n184), .B1(n29379), .ZN(n185) );
  I_NAND2 U826 ( .A1(n187), .B1(n29379), .ZN(n188) );
  I_NAND2 U827 ( .A1(n190), .B1(n29379), .ZN(n191) );
  I_NAND2 U828 ( .A1(n193), .B1(n29379), .ZN(n194) );
  I_NAND2 U829 ( .A1(n196), .B1(n29380), .ZN(n197) );
  I_NAND2 U830 ( .A1(n199), .B1(n29380), .ZN(n200) );
  I_NAND2 U831 ( .A1(n202), .B1(n29380), .ZN(n203) );
  I_NAND2 U832 ( .A1(n205), .B1(n29380), .ZN(n206) );
  I_NAND2 U833 ( .A1(n208), .B1(n29380), .ZN(n209) );
  I_NAND2 U834 ( .A1(n211), .B1(n29380), .ZN(n212) );
  I_NAND2 U835 ( .A1(n216), .B1(n29380), .ZN(n217) );
  I_NAND2 U836 ( .A1(n219), .B1(n29380), .ZN(n220) );
  I_NAND2 U837 ( .A1(n221), .B1(n29380), .ZN(n222) );
  I_NAND2 U838 ( .A1(n223), .B1(n29380), .ZN(n224) );
  I_NAND2 U839 ( .A1(n225), .B1(n29380), .ZN(n226) );
  I_NAND2 U840 ( .A1(n227), .B1(n29381), .ZN(n228) );
  I_NAND2 U841 ( .A1(n229), .B1(n29381), .ZN(n230) );
  I_NAND2 U842 ( .A1(n231), .B1(n29381), .ZN(n232) );
  I_NAND2 U843 ( .A1(n233), .B1(n29381), .ZN(n234) );
  I_NAND2 U844 ( .A1(n235), .B1(n29381), .ZN(n236) );
  I_NAND2 U845 ( .A1(n237), .B1(n29381), .ZN(n238) );
  I_NAND2 U846 ( .A1(n239), .B1(n29381), .ZN(n240) );
  I_NAND2 U847 ( .A1(n241), .B1(n29381), .ZN(n242) );
  I_NAND2 U848 ( .A1(n243), .B1(n29381), .ZN(n244) );
  I_NAND2 U849 ( .A1(n245), .B1(n29381), .ZN(n246) );
  I_NAND2 U850 ( .A1(n247), .B1(n29381), .ZN(n248) );
  I_NAND2 U851 ( .A1(n249), .B1(n29381), .ZN(n250) );
  I_NAND2 U852 ( .A1(n251), .B1(n29382), .ZN(n252) );
  I_NAND2 U853 ( .A1(n253), .B1(n29382), .ZN(n254) );
  I_NAND2 U854 ( .A1(n255), .B1(n29382), .ZN(n256) );
  I_NAND2 U855 ( .A1(n257), .B1(n29382), .ZN(n258) );
  I_NAND2 U856 ( .A1(n259), .B1(n29382), .ZN(n260) );
  I_NAND2 U857 ( .A1(n261), .B1(n29382), .ZN(n262) );
  I_NAND2 U858 ( .A1(n263), .B1(n29382), .ZN(n264) );
  I_NAND2 U859 ( .A1(n265), .B1(n29382), .ZN(n266) );
  I_NAND2 U860 ( .A1(n267), .B1(n29382), .ZN(n268) );
  I_NAND2 U861 ( .A1(n269), .B1(n29382), .ZN(n270) );
  I_NAND2 U862 ( .A1(n271), .B1(n29382), .ZN(n272) );
  I_NAND2 U863 ( .A1(n273), .B1(n29382), .ZN(n274) );
  I_NAND2 U864 ( .A1(n275), .B1(n29383), .ZN(n276) );
  I_NAND2 U865 ( .A1(n277), .B1(n29383), .ZN(n278) );
  I_NAND2 U866 ( .A1(n279), .B1(n29383), .ZN(n280) );
  I_NAND2 U867 ( .A1(n281), .B1(n29383), .ZN(n282) );
  I_NAND2 U868 ( .A1(n283), .B1(n29383), .ZN(n284) );
  I_NAND2 U869 ( .A1(n285), .B1(n29383), .ZN(n286) );
  I_NAND2 U870 ( .A1(n287), .B1(n29383), .ZN(n288) );
  I_NAND2 U871 ( .A1(n289), .B1(n29383), .ZN(n290) );
  I_NAND2 U872 ( .A1(n291), .B1(n29383), .ZN(n292) );
  I_NAND2 U873 ( .A1(n293), .B1(n29383), .ZN(n294) );
  I_NAND2 U874 ( .A1(n295), .B1(n29383), .ZN(n296) );
  I_NAND2 U875 ( .A1(n297), .B1(n29383), .ZN(n298) );
  I_NAND2 U876 ( .A1(n299), .B1(n29384), .ZN(n300) );
  I_NAND2 U877 ( .A1(n301), .B1(n29384), .ZN(n302) );
  I_NAND2 U878 ( .A1(n303), .B1(n29384), .ZN(n304) );
  I_NAND2 U879 ( .A1(n305), .B1(n29384), .ZN(n306) );
  I_NAND2 U880 ( .A1(n307), .B1(n29384), .ZN(n308) );
  I_NAND2 U881 ( .A1(n309), .B1(n29384), .ZN(n310) );
  I_NAND2 U882 ( .A1(n311), .B1(n29384), .ZN(n312) );
  I_NAND2 U883 ( .A1(n313), .B1(n29384), .ZN(n314) );
  I_NAND2 U884 ( .A1(n315), .B1(n29384), .ZN(n316) );
  I_NAND2 U885 ( .A1(n317), .B1(n29384), .ZN(n318) );
  I_NAND2 U886 ( .A1(n319), .B1(n29384), .ZN(n320) );
  I_NAND2 U887 ( .A1(n321), .B1(n29384), .ZN(n322) );
  I_NAND2 U888 ( .A1(n323), .B1(n29385), .ZN(n324) );
  I_NAND2 U889 ( .A1(n325), .B1(n29385), .ZN(n326) );
  I_NAND2 U890 ( .A1(n327), .B1(n29385), .ZN(n328) );
  I_NAND2 U891 ( .A1(n329), .B1(n29385), .ZN(n330) );
  I_NAND2 U892 ( .A1(n331), .B1(n29385), .ZN(n332) );
  I_NAND2 U893 ( .A1(n333), .B1(n29385), .ZN(n334) );
  I_NAND2 U894 ( .A1(n335), .B1(n29385), .ZN(n336) );
  I_NAND2 U895 ( .A1(n337), .B1(n29385), .ZN(n338) );
  I_NAND2 U896 ( .A1(n339), .B1(n29385), .ZN(n340) );
  I_NAND2 U897 ( .A1(n341), .B1(n29385), .ZN(n342) );
  I_NAND2 U898 ( .A1(n343), .B1(n29385), .ZN(n344) );
  I_NAND2 U899 ( .A1(n346), .B1(n29385), .ZN(n347) );
  I_NAND2 U900 ( .A1(n349), .B1(n29386), .ZN(n350) );
  I_NAND2 U901 ( .A1(n351), .B1(n29386), .ZN(n352) );
  I_NAND2 U902 ( .A1(n353), .B1(n29370), .ZN(n354) );
  I_NAND2 U903 ( .A1(n355), .B1(n29364), .ZN(n356) );
  I_NAND2 U904 ( .A1(n357), .B1(n29364), .ZN(n358) );
  I_NAND2 U905 ( .A1(n359), .B1(n29365), .ZN(n360) );
  I_NAND2 U906 ( .A1(n361), .B1(n29365), .ZN(n362) );
  I_NAND2 U907 ( .A1(n363), .B1(n29365), .ZN(n364) );
  I_NAND2 U908 ( .A1(n365), .B1(n29365), .ZN(n366) );
  I_NAND2 U909 ( .A1(n367), .B1(n29365), .ZN(n368) );
  I_NAND2 U910 ( .A1(n369), .B1(n29365), .ZN(n370) );
  I_NAND2 U911 ( .A1(n371), .B1(n29365), .ZN(n372) );
  I_NAND2 U912 ( .A1(n373), .B1(n29365), .ZN(n374) );
  I_NAND2 U913 ( .A1(n375), .B1(n29365), .ZN(n376) );
  I_NAND2 U914 ( .A1(n377), .B1(n29365), .ZN(n378) );
  I_NAND2 U915 ( .A1(n379), .B1(n29365), .ZN(n380) );
  I_NAND2 U916 ( .A1(n381), .B1(n29365), .ZN(n382) );
  I_NAND2 U917 ( .A1(n383), .B1(n29366), .ZN(n384) );
  I_NAND2 U918 ( .A1(n385), .B1(n29366), .ZN(n386) );
  I_NAND2 U919 ( .A1(n387), .B1(n29366), .ZN(n388) );
  I_NAND2 U920 ( .A1(n389), .B1(n29366), .ZN(n390) );
  I_NAND2 U921 ( .A1(n391), .B1(n29366), .ZN(n392) );
  I_NAND2 U922 ( .A1(n393), .B1(n29366), .ZN(n394) );
  I_NAND2 U923 ( .A1(n395), .B1(n29366), .ZN(n396) );
  I_NAND2 U924 ( .A1(n397), .B1(n29366), .ZN(n398) );
  I_NAND2 U925 ( .A1(n399), .B1(n29366), .ZN(n400) );
  I_NAND2 U926 ( .A1(n401), .B1(n29366), .ZN(n402) );
  I_NAND2 U927 ( .A1(n403), .B1(n29366), .ZN(n404) );
  I_NAND2 U928 ( .A1(n405), .B1(n29366), .ZN(n406) );
  I_NAND2 U929 ( .A1(n407), .B1(n29367), .ZN(n408) );
  I_NAND2 U930 ( .A1(n409), .B1(n29367), .ZN(n410) );
  I_NAND2 U931 ( .A1(n411), .B1(n29367), .ZN(n412) );
  I_NAND2 U932 ( .A1(n413), .B1(n29367), .ZN(n414) );
  I_NAND2 U933 ( .A1(n415), .B1(n29367), .ZN(n416) );
  I_NAND2 U934 ( .A1(n417), .B1(n29367), .ZN(n418) );
  I_NAND2 U935 ( .A1(n419), .B1(n29367), .ZN(n420) );
  I_NAND2 U936 ( .A1(n421), .B1(n29367), .ZN(n422) );
  I_NAND2 U937 ( .A1(n423), .B1(n29367), .ZN(n424) );
  I_NAND2 U938 ( .A1(n425), .B1(n29367), .ZN(n426) );
  I_NAND2 U939 ( .A1(n427), .B1(n29367), .ZN(n428) );
  I_NAND2 U940 ( .A1(n429), .B1(n29367), .ZN(n430) );
  I_NAND2 U941 ( .A1(n431), .B1(n29368), .ZN(n432) );
  I_NAND2 U942 ( .A1(n433), .B1(n29368), .ZN(n434) );
  I_NAND2 U943 ( .A1(n435), .B1(n29368), .ZN(n436) );
  I_NAND2 U944 ( .A1(n437), .B1(n29368), .ZN(n438) );
  I_NAND2 U945 ( .A1(n439), .B1(n29368), .ZN(n440) );
  I_NAND2 U946 ( .A1(n441), .B1(n29368), .ZN(n442) );
  I_NAND2 U947 ( .A1(n443), .B1(n29368), .ZN(n444) );
  I_NAND2 U948 ( .A1(n445), .B1(n29368), .ZN(n446) );
  I_NAND2 U949 ( .A1(n447), .B1(n29368), .ZN(n448) );
  I_NAND2 U950 ( .A1(n449), .B1(n29368), .ZN(n450) );
  I_NAND2 U951 ( .A1(n451), .B1(n29368), .ZN(n452) );
  I_NAND2 U952 ( .A1(n453), .B1(n29368), .ZN(n454) );
  I_NAND2 U953 ( .A1(n455), .B1(n29369), .ZN(n456) );
  I_NAND2 U954 ( .A1(n457), .B1(n29369), .ZN(n458) );
  I_NAND2 U955 ( .A1(n459), .B1(n29369), .ZN(n460) );
  I_NAND2 U956 ( .A1(n461), .B1(n29369), .ZN(n462) );
  I_NAND2 U957 ( .A1(n463), .B1(n29369), .ZN(n464) );
  I_NAND2 U958 ( .A1(n465), .B1(n29369), .ZN(n466) );
  I_NAND2 U959 ( .A1(n467), .B1(n29369), .ZN(n468) );
  I_NAND2 U960 ( .A1(n469), .B1(n29369), .ZN(n470) );
  I_NAND2 U961 ( .A1(n471), .B1(n29369), .ZN(n472) );
  I_NAND2 U962 ( .A1(n473), .B1(n29369), .ZN(n474) );
  I_NAND2 U963 ( .A1(n476), .B1(n29369), .ZN(n477) );
  I_NAND2 U964 ( .A1(n479), .B1(n29369), .ZN(n480) );
  I_NAND2 U965 ( .A1(n481), .B1(n29370), .ZN(n482) );
  I_NAND2 U966 ( .A1(n483), .B1(n29370), .ZN(n484) );
  I_NAND2 U967 ( .A1(n485), .B1(n29370), .ZN(n486) );
  I_NAND2 U968 ( .A1(n487), .B1(n29370), .ZN(n488) );
  I_NAND2 U969 ( .A1(n489), .B1(n29370), .ZN(n490) );
  I_NAND2 U970 ( .A1(n491), .B1(n29370), .ZN(n492) );
  I_NAND2 U971 ( .A1(n493), .B1(n29370), .ZN(n494) );
  I_NAND2 U972 ( .A1(n495), .B1(n29370), .ZN(n496) );
  I_NAND2 U973 ( .A1(n497), .B1(n29370), .ZN(n498) );
  I_NAND2 U974 ( .A1(n499), .B1(n29370), .ZN(n500) );
  I_NAND2 U975 ( .A1(n501), .B1(n29370), .ZN(n502) );
  I_NAND2 U976 ( .A1(n503), .B1(n29371), .ZN(n504) );
  I_NAND2 U977 ( .A1(n505), .B1(n29371), .ZN(n506) );
  I_NAND2 U978 ( .A1(n507), .B1(n29371), .ZN(n508) );
  I_NAND2 U979 ( .A1(n509), .B1(n29371), .ZN(n510) );
  I_NAND2 U980 ( .A1(n511), .B1(n29371), .ZN(n512) );
  I_NAND2 U981 ( .A1(n513), .B1(n29371), .ZN(n514) );
  I_NAND2 U982 ( .A1(n515), .B1(n29371), .ZN(n516) );
  I_NAND2 U983 ( .A1(n517), .B1(n29371), .ZN(n518) );
  I_NAND2 U984 ( .A1(n519), .B1(n29371), .ZN(n520) );
  I_NAND2 U985 ( .A1(n521), .B1(n29371), .ZN(n522) );
  I_NAND2 U986 ( .A1(n523), .B1(n29371), .ZN(n524) );
  I_NAND2 U987 ( .A1(n525), .B1(n29371), .ZN(n526) );
  I_NAND2 U988 ( .A1(n527), .B1(n29372), .ZN(n528) );
  I_NAND2 U989 ( .A1(n529), .B1(n29372), .ZN(n530) );
  I_NAND2 U990 ( .A1(n531), .B1(n29372), .ZN(n532) );
  I_NAND2 U991 ( .A1(n533), .B1(n29372), .ZN(n534) );
  I_NAND2 U992 ( .A1(n535), .B1(n29372), .ZN(n536) );
  I_NAND2 U993 ( .A1(n537), .B1(n29372), .ZN(n538) );
  I_NAND2 U994 ( .A1(n539), .B1(n29372), .ZN(n540) );
  I_NAND2 U995 ( .A1(n541), .B1(n29372), .ZN(n542) );
  I_NAND2 U996 ( .A1(n543), .B1(n29372), .ZN(n544) );
  I_NAND2 U997 ( .A1(n545), .B1(n29372), .ZN(n546) );
  I_NAND2 U998 ( .A1(n547), .B1(n29372), .ZN(n548) );
  I_NAND2 U999 ( .A1(n549), .B1(n29372), .ZN(n550) );
  I_NAND2 U1000 ( .A1(n551), .B1(n29373), .ZN(n552) );
  I_NAND2 U1001 ( .A1(n553), .B1(n29373), .ZN(n554) );
  I_NAND2 U1002 ( .A1(n555), .B1(n29373), .ZN(n556) );
  I_NAND2 U1003 ( .A1(n557), .B1(n29373), .ZN(n558) );
  I_NAND2 U1004 ( .A1(n559), .B1(n29373), .ZN(n560) );
  I_NAND2 U1005 ( .A1(n561), .B1(n29373), .ZN(n562) );
  I_NAND2 U1006 ( .A1(n563), .B1(n29373), .ZN(n564) );
  I_NAND2 U1007 ( .A1(n565), .B1(n29373), .ZN(n566) );
  I_NAND2 U1008 ( .A1(n567), .B1(n29373), .ZN(n568) );
  I_NAND2 U1009 ( .A1(n569), .B1(n29373), .ZN(n570) );
  I_NAND2 U1010 ( .A1(n571), .B1(n29373), .ZN(n572) );
  I_NAND2 U1011 ( .A1(n573), .B1(n29373), .ZN(n574) );
  I_NAND2 U1012 ( .A1(n575), .B1(n29374), .ZN(n576) );
  I_NAND2 U1013 ( .A1(n577), .B1(n29374), .ZN(n578) );
  I_NAND2 U1014 ( .A1(n579), .B1(n29374), .ZN(n580) );
  I_NAND2 U1015 ( .A1(n581), .B1(n29374), .ZN(n582) );
  I_NAND2 U1016 ( .A1(n583), .B1(n29374), .ZN(n584) );
  I_NAND2 U1017 ( .A1(n585), .B1(n29374), .ZN(n586) );
  I_NAND2 U1018 ( .A1(n587), .B1(n29374), .ZN(n588) );
  I_NAND2 U1019 ( .A1(n589), .B1(n29374), .ZN(n590) );
  I_NAND2 U1020 ( .A1(n591), .B1(n29374), .ZN(n592) );
  I_NAND2 U1021 ( .A1(n593), .B1(n29374), .ZN(n594) );
  I_NAND2 U1022 ( .A1(n595), .B1(n29374), .ZN(n596) );
  I_NAND2 U1023 ( .A1(n597), .B1(n29374), .ZN(n598) );
  I_NAND2 U1024 ( .A1(n599), .B1(n29375), .ZN(n600) );
  I_NAND2 U1025 ( .A1(n601), .B1(n29375), .ZN(n602) );
  I_NAND2 U1026 ( .A1(n603), .B1(n29375), .ZN(n604) );
  I_NAND2 U1027 ( .A1(n606), .B1(n29375), .ZN(n607) );
  I_NAND2 U1028 ( .A1(n609), .B1(n29375), .ZN(n610) );
  I_NAND2 U1029 ( .A1(n611), .B1(n29375), .ZN(n612) );
  I_NAND2 U1030 ( .A1(n613), .B1(n29402), .ZN(n614) );
  I_NAND2 U1031 ( .A1(n615), .B1(n29396), .ZN(n616) );
  I_NAND2 U1032 ( .A1(n617), .B1(n29397), .ZN(n618) );
  I_NAND2 U1033 ( .A1(n619), .B1(n29397), .ZN(n620) );
  I_NAND2 U1034 ( .A1(n621), .B1(n29397), .ZN(n622) );
  I_NAND2 U1035 ( .A1(n623), .B1(n29397), .ZN(n624) );
  I_NAND2 U1036 ( .A1(n625), .B1(n29397), .ZN(n626) );
  I_NAND2 U1037 ( .A1(n627), .B1(n29397), .ZN(n628) );
  I_NAND2 U1038 ( .A1(n629), .B1(n29397), .ZN(n630) );
  I_NAND2 U1039 ( .A1(n631), .B1(n29397), .ZN(n632) );
  I_NAND2 U1040 ( .A1(n633), .B1(n29397), .ZN(n634) );
  I_NAND2 U1041 ( .A1(n635), .B1(n29397), .ZN(n636) );
  I_NAND2 U1042 ( .A1(n637), .B1(n29397), .ZN(n638) );
  I_NAND2 U1043 ( .A1(n639), .B1(n29397), .ZN(n640) );
  I_NAND2 U1044 ( .A1(n641), .B1(n29398), .ZN(n642) );
  I_NAND2 U1045 ( .A1(n643), .B1(n29398), .ZN(n644) );
  I_NAND2 U1046 ( .A1(n645), .B1(n29398), .ZN(n646) );
  I_NAND2 U1047 ( .A1(n647), .B1(n29398), .ZN(n648) );
  I_NAND2 U1048 ( .A1(n649), .B1(n29398), .ZN(n650) );
  I_NAND2 U1049 ( .A1(n651), .B1(n29398), .ZN(n652) );
  I_NAND2 U1050 ( .A1(n653), .B1(n29398), .ZN(n654) );
  I_NAND2 U1051 ( .A1(n655), .B1(n29398), .ZN(n656) );
  I_NAND2 U1052 ( .A1(n657), .B1(n29398), .ZN(n658) );
  I_NAND2 U1053 ( .A1(n659), .B1(n29398), .ZN(n660) );
  I_NAND2 U1054 ( .A1(n661), .B1(n29398), .ZN(n662) );
  I_NAND2 U1055 ( .A1(n663), .B1(n29398), .ZN(n664) );
  I_NAND2 U1056 ( .A1(n665), .B1(n29399), .ZN(n666) );
  I_NAND2 U1057 ( .A1(n667), .B1(n29399), .ZN(n668) );
  I_NAND2 U1058 ( .A1(n669), .B1(n29399), .ZN(n670) );
  I_NAND2 U1059 ( .A1(n671), .B1(n29399), .ZN(n672) );
  I_NAND2 U1060 ( .A1(n673), .B1(n29399), .ZN(n674) );
  I_NAND2 U1061 ( .A1(n675), .B1(n29399), .ZN(n676) );
  I_NAND2 U1062 ( .A1(n677), .B1(n29399), .ZN(n678) );
  I_NAND2 U1063 ( .A1(n679), .B1(n29399), .ZN(n680) );
  I_NAND2 U1064 ( .A1(n681), .B1(n29399), .ZN(n682) );
  I_NAND2 U1065 ( .A1(n683), .B1(n29399), .ZN(n684) );
  I_NAND2 U1066 ( .A1(n685), .B1(n29399), .ZN(n686) );
  I_NAND2 U1067 ( .A1(n687), .B1(n29399), .ZN(n688) );
  I_NAND2 U1068 ( .A1(n689), .B1(n29400), .ZN(n690) );
  I_NAND2 U1069 ( .A1(n691), .B1(n29400), .ZN(n692) );
  I_NAND2 U1070 ( .A1(n693), .B1(n29400), .ZN(n694) );
  I_NAND2 U1071 ( .A1(n695), .B1(n29400), .ZN(n696) );
  I_NAND2 U1072 ( .A1(n697), .B1(n29400), .ZN(n698) );
  I_NAND2 U1073 ( .A1(n699), .B1(n29400), .ZN(n700) );
  I_NAND2 U1074 ( .A1(n701), .B1(n29400), .ZN(n702) );
  I_NAND2 U1075 ( .A1(n703), .B1(n29400), .ZN(n704) );
  I_NAND2 U1076 ( .A1(n705), .B1(n29400), .ZN(n706) );
  I_NAND2 U1077 ( .A1(n707), .B1(n29400), .ZN(n708) );
  I_NAND2 U1078 ( .A1(n709), .B1(n29400), .ZN(n710) );
  I_NAND2 U1079 ( .A1(n711), .B1(n29400), .ZN(n712) );
  I_NAND2 U1080 ( .A1(n713), .B1(n29401), .ZN(n714) );
  I_NAND2 U1081 ( .A1(n715), .B1(n29401), .ZN(n716) );
  I_NAND2 U1082 ( .A1(n717), .B1(n29401), .ZN(n718) );
  I_NAND2 U1083 ( .A1(n719), .B1(n29401), .ZN(n720) );
  I_NAND2 U1084 ( .A1(n721), .B1(n29401), .ZN(n722) );
  I_NAND2 U1085 ( .A1(n723), .B1(n29401), .ZN(n724) );
  I_NAND2 U1086 ( .A1(n725), .B1(n29401), .ZN(n726) );
  I_NAND2 U1087 ( .A1(n727), .B1(n29401), .ZN(n728) );
  I_NAND2 U1088 ( .A1(n729), .B1(n29401), .ZN(n730) );
  I_NAND2 U1089 ( .A1(n731), .B1(n29401), .ZN(n732) );
  I_NAND2 U1090 ( .A1(n733), .B1(n29401), .ZN(n734) );
  I_NAND2 U1091 ( .A1(n736), .B1(n29401), .ZN(n737) );
  I_NAND2 U1092 ( .A1(n739), .B1(n29402), .ZN(n740) );
  I_NAND2 U1093 ( .A1(n741), .B1(n29402), .ZN(n742) );
  I_NAND2 U1094 ( .A1(n743), .B1(n29402), .ZN(n744) );
  I_NAND2 U1095 ( .A1(n745), .B1(n29402), .ZN(n746) );
  I_NAND2 U1096 ( .A1(n747), .B1(n29402), .ZN(n748) );
  I_NAND2 U1097 ( .A1(n749), .B1(n29402), .ZN(n750) );
  I_NAND2 U1098 ( .A1(n751), .B1(n29402), .ZN(n752) );
  I_NAND2 U1099 ( .A1(n753), .B1(n29402), .ZN(n754) );
  I_NAND2 U1100 ( .A1(n755), .B1(n29402), .ZN(n756) );
  I_NAND2 U1101 ( .A1(n757), .B1(n29402), .ZN(n758) );
  I_NAND2 U1102 ( .A1(n759), .B1(n29402), .ZN(n760) );
  I_NAND2 U1103 ( .A1(n761), .B1(n29403), .ZN(n762) );
  I_NAND2 U1104 ( .A1(n763), .B1(n29403), .ZN(n764) );
  I_NAND2 U1105 ( .A1(n765), .B1(n29403), .ZN(n766) );
  I_NAND2 U1106 ( .A1(n767), .B1(n29403), .ZN(n768) );
  I_NAND2 U1107 ( .A1(n769), .B1(n29403), .ZN(n770) );
  I_NAND2 U1108 ( .A1(n771), .B1(n29403), .ZN(n772) );
  I_NAND2 U1109 ( .A1(n773), .B1(n29403), .ZN(n774) );
  I_NAND2 U1110 ( .A1(n775), .B1(n29403), .ZN(n776) );
  I_NAND2 U1111 ( .A1(n777), .B1(n29403), .ZN(n778) );
  I_NAND2 U1112 ( .A1(n779), .B1(n29403), .ZN(n780) );
  I_NAND2 U1113 ( .A1(n781), .B1(n29403), .ZN(n782) );
  I_NAND2 U1114 ( .A1(n783), .B1(n29403), .ZN(n784) );
  I_NAND2 U1115 ( .A1(n785), .B1(n29404), .ZN(n786) );
  I_NAND2 U1116 ( .A1(n787), .B1(n29404), .ZN(n788) );
  I_NAND2 U1117 ( .A1(n789), .B1(n29404), .ZN(n790) );
  I_NAND2 U1118 ( .A1(n791), .B1(n29404), .ZN(n792) );
  I_NAND2 U1119 ( .A1(n793), .B1(n29404), .ZN(n794) );
  I_NAND2 U1120 ( .A1(n795), .B1(n29404), .ZN(n796) );
  I_NAND2 U1121 ( .A1(n797), .B1(n29404), .ZN(n798) );
  I_NAND2 U1122 ( .A1(n799), .B1(n29404), .ZN(n800) );
  I_NAND2 U1123 ( .A1(n801), .B1(n29404), .ZN(n802) );
  I_NAND2 U1124 ( .A1(n803), .B1(n29404), .ZN(n804) );
  I_NAND2 U1125 ( .A1(n805), .B1(n29404), .ZN(n806) );
  I_NAND2 U1126 ( .A1(n807), .B1(n29404), .ZN(n808) );
  I_NAND2 U1127 ( .A1(n809), .B1(n29405), .ZN(n810) );
  I_NAND2 U1128 ( .A1(n811), .B1(n29405), .ZN(n812) );
  I_NAND2 U1129 ( .A1(n813), .B1(n29405), .ZN(n814) );
  I_NAND2 U1130 ( .A1(n815), .B1(n29405), .ZN(n816) );
  I_NAND2 U1131 ( .A1(n817), .B1(n29405), .ZN(n818) );
  I_NAND2 U1132 ( .A1(n819), .B1(n29405), .ZN(n820) );
  I_NAND2 U1133 ( .A1(n821), .B1(n29405), .ZN(n822) );
  I_NAND2 U1134 ( .A1(n823), .B1(n29405), .ZN(n824) );
  I_NAND2 U1135 ( .A1(n825), .B1(n29405), .ZN(n826) );
  I_NAND2 U1136 ( .A1(n827), .B1(n29405), .ZN(n828) );
  I_NAND2 U1137 ( .A1(n829), .B1(n29405), .ZN(n830) );
  I_NAND2 U1138 ( .A1(n831), .B1(n29405), .ZN(n832) );
  I_NAND2 U1139 ( .A1(n833), .B1(n29406), .ZN(n834) );
  I_NAND2 U1140 ( .A1(n835), .B1(n29406), .ZN(n836) );
  I_NAND2 U1141 ( .A1(n837), .B1(n29406), .ZN(n838) );
  I_NAND2 U1142 ( .A1(n839), .B1(n29406), .ZN(n840) );
  I_NAND2 U1143 ( .A1(n841), .B1(n29406), .ZN(n842) );
  I_NAND2 U1144 ( .A1(n843), .B1(n29406), .ZN(n844) );
  I_NAND2 U1145 ( .A1(n845), .B1(n29406), .ZN(n846) );
  I_NAND2 U1146 ( .A1(n847), .B1(n29406), .ZN(n848) );
  I_NAND2 U1147 ( .A1(n849), .B1(n29406), .ZN(n850) );
  I_NAND2 U1148 ( .A1(n851), .B1(n29406), .ZN(n852) );
  I_NAND2 U1149 ( .A1(n853), .B1(n29406), .ZN(n854) );
  I_NAND2 U1150 ( .A1(n855), .B1(n29406), .ZN(n856) );
  I_NAND2 U1151 ( .A1(n857), .B1(n29407), .ZN(n858) );
  I_NAND2 U1152 ( .A1(n859), .B1(n29407), .ZN(n860) );
  I_NAND2 U1153 ( .A1(n861), .B1(n29407), .ZN(n862) );
  I_NAND2 U1154 ( .A1(n863), .B1(n29407), .ZN(n864) );
  I_NAND2 U1155 ( .A1(n866), .B1(n29407), .ZN(n867) );
  I_NAND2 U1156 ( .A1(n869), .B1(n29407), .ZN(n870) );
  I_NAND2 U1157 ( .A1(n871), .B1(n29407), .ZN(n872) );
  I_NAND2 U1158 ( .A1(n873), .B1(n29391), .ZN(n874) );
  I_NAND2 U1159 ( .A1(n875), .B1(n29386), .ZN(n876) );
  I_NAND2 U1160 ( .A1(n877), .B1(n29386), .ZN(n878) );
  I_NAND2 U1161 ( .A1(n879), .B1(n29386), .ZN(n880) );
  I_NAND2 U1162 ( .A1(n881), .B1(n29386), .ZN(n882) );
  I_NAND2 U1163 ( .A1(n883), .B1(n29386), .ZN(n884) );
  I_NAND2 U1164 ( .A1(n885), .B1(n29386), .ZN(n886) );
  I_NAND2 U1165 ( .A1(n887), .B1(n29386), .ZN(n888) );
  I_NAND2 U1166 ( .A1(n889), .B1(n29386), .ZN(n890) );
  I_NAND2 U1167 ( .A1(n891), .B1(n29386), .ZN(n892) );
  I_NAND2 U1168 ( .A1(n893), .B1(n29387), .ZN(n894) );
  I_NAND2 U1169 ( .A1(n895), .B1(n29387), .ZN(n896) );
  I_NAND2 U1170 ( .A1(n897), .B1(n29387), .ZN(n898) );
  I_NAND2 U1171 ( .A1(n899), .B1(n29387), .ZN(n900) );
  I_NAND2 U1172 ( .A1(n901), .B1(n29387), .ZN(n902) );
  I_NAND2 U1173 ( .A1(n903), .B1(n29387), .ZN(n904) );
  I_NAND2 U1174 ( .A1(n905), .B1(n29387), .ZN(n906) );
  I_NAND2 U1175 ( .A1(n907), .B1(n29387), .ZN(n908) );
  I_NAND2 U1176 ( .A1(n909), .B1(n29387), .ZN(n910) );
  I_NAND2 U1177 ( .A1(n911), .B1(n29387), .ZN(n912) );
  I_NAND2 U1178 ( .A1(n913), .B1(n29387), .ZN(n914) );
  I_NAND2 U1179 ( .A1(n915), .B1(n29387), .ZN(n916) );
  I_NAND2 U1180 ( .A1(n917), .B1(n29388), .ZN(n918) );
  I_NAND2 U1181 ( .A1(n919), .B1(n29388), .ZN(n920) );
  I_NAND2 U1182 ( .A1(n921), .B1(n29388), .ZN(n922) );
  I_NAND2 U1183 ( .A1(n923), .B1(n29388), .ZN(n924) );
  I_NAND2 U1184 ( .A1(n925), .B1(n29388), .ZN(n926) );
  I_NAND2 U1185 ( .A1(n927), .B1(n29388), .ZN(n928) );
  I_NAND2 U1186 ( .A1(n929), .B1(n29388), .ZN(n930) );
  I_NAND2 U1187 ( .A1(n931), .B1(n29388), .ZN(n932) );
  I_NAND2 U1188 ( .A1(n933), .B1(n29388), .ZN(n934) );
  I_NAND2 U1189 ( .A1(n935), .B1(n29388), .ZN(n936) );
  I_NAND2 U1190 ( .A1(n937), .B1(n29388), .ZN(n938) );
  I_NAND2 U1191 ( .A1(n939), .B1(n29388), .ZN(n940) );
  I_NAND2 U1192 ( .A1(n941), .B1(n29389), .ZN(n942) );
  I_NAND2 U1193 ( .A1(n943), .B1(n29389), .ZN(n944) );
  I_NAND2 U1194 ( .A1(n945), .B1(n29389), .ZN(n946) );
  I_NAND2 U1195 ( .A1(n947), .B1(n29389), .ZN(n948) );
  I_NAND2 U1196 ( .A1(n949), .B1(n29389), .ZN(n950) );
  I_NAND2 U1197 ( .A1(n951), .B1(n29389), .ZN(n952) );
  I_NAND2 U1198 ( .A1(n953), .B1(n29389), .ZN(n954) );
  I_NAND2 U1199 ( .A1(n955), .B1(n29389), .ZN(n956) );
  I_NAND2 U1200 ( .A1(n957), .B1(n29389), .ZN(n958) );
  I_NAND2 U1201 ( .A1(n959), .B1(n29389), .ZN(n960) );
  I_NAND2 U1202 ( .A1(n961), .B1(n29389), .ZN(n962) );
  I_NAND2 U1203 ( .A1(n963), .B1(n29389), .ZN(n964) );
  I_NAND2 U1204 ( .A1(n965), .B1(n29390), .ZN(n966) );
  I_NAND2 U1205 ( .A1(n967), .B1(n29390), .ZN(n968) );
  I_NAND2 U1206 ( .A1(n969), .B1(n29390), .ZN(n970) );
  I_NAND2 U1207 ( .A1(n971), .B1(n29390), .ZN(n972) );
  I_NAND2 U1208 ( .A1(n973), .B1(n29390), .ZN(n974) );
  I_NAND2 U1209 ( .A1(n975), .B1(n29390), .ZN(n976) );
  I_NAND2 U1210 ( .A1(n977), .B1(n29390), .ZN(n978) );
  I_NAND2 U1211 ( .A1(n979), .B1(n29390), .ZN(n980) );
  I_NAND2 U1212 ( .A1(n981), .B1(n29390), .ZN(n982) );
  I_NAND2 U1213 ( .A1(n983), .B1(n29390), .ZN(n984) );
  I_NAND2 U1214 ( .A1(n985), .B1(n29390), .ZN(n986) );
  I_NAND2 U1215 ( .A1(n987), .B1(n29390), .ZN(n988) );
  I_NAND2 U1216 ( .A1(n989), .B1(n29391), .ZN(n990) );
  I_NAND2 U1217 ( .A1(n991), .B1(n29391), .ZN(n992) );
  I_NAND2 U1218 ( .A1(n993), .B1(n29391), .ZN(n994) );
  I_NAND2 U1219 ( .A1(n996), .B1(n29391), .ZN(n997) );
  I_NAND2 U1220 ( .A1(n999), .B1(n29391), .ZN(n1000) );
  I_NAND2 U1221 ( .A1(n1001), .B1(n29391), .ZN(n1002) );
  I_NAND2 U1222 ( .A1(n1003), .B1(n29391), .ZN(n1004) );
  I_NAND2 U1223 ( .A1(n1005), .B1(n29391), .ZN(n1006) );
  I_NAND2 U1224 ( .A1(n1007), .B1(n29391), .ZN(n1008) );
  I_NAND2 U1225 ( .A1(n1009), .B1(n29391), .ZN(n1010) );
  I_NAND2 U1226 ( .A1(n1011), .B1(n29391), .ZN(n1012) );
  I_NAND2 U1227 ( .A1(n1013), .B1(n29392), .ZN(n1014) );
  I_NAND2 U1228 ( .A1(n1015), .B1(n29392), .ZN(n1016) );
  I_NAND2 U1229 ( .A1(n1017), .B1(n29392), .ZN(n1018) );
  I_NAND2 U1230 ( .A1(n1019), .B1(n29392), .ZN(n1020) );
  I_NAND2 U1231 ( .A1(n1021), .B1(n29392), .ZN(n1022) );
  I_NAND2 U1232 ( .A1(n1023), .B1(n29392), .ZN(n1024) );
  I_NAND2 U1233 ( .A1(n1025), .B1(n29392), .ZN(n1026) );
  I_NAND2 U1234 ( .A1(n1027), .B1(n29392), .ZN(n1028) );
  I_NAND2 U1235 ( .A1(n1029), .B1(n29392), .ZN(n1030) );
  I_NAND2 U1236 ( .A1(n1031), .B1(n29392), .ZN(n1032) );
  I_NAND2 U1237 ( .A1(n1033), .B1(n29392), .ZN(n1034) );
  I_NAND2 U1238 ( .A1(n1035), .B1(n29392), .ZN(n1036) );
  I_NAND2 U1239 ( .A1(n1037), .B1(n29393), .ZN(n1038) );
  I_NAND2 U1240 ( .A1(n1039), .B1(n29393), .ZN(n1040) );
  I_NAND2 U1241 ( .A1(n1041), .B1(n29393), .ZN(n1042) );
  I_NAND2 U1242 ( .A1(n1043), .B1(n29393), .ZN(n1044) );
  I_NAND2 U1243 ( .A1(n1045), .B1(n29393), .ZN(n1046) );
  I_NAND2 U1244 ( .A1(n1047), .B1(n29393), .ZN(n1048) );
  I_NAND2 U1245 ( .A1(n1049), .B1(n29393), .ZN(n1050) );
  I_NAND2 U1246 ( .A1(n1051), .B1(n29393), .ZN(n1052) );
  I_NAND2 U1247 ( .A1(n1053), .B1(n29393), .ZN(n1054) );
  I_NAND2 U1248 ( .A1(n1055), .B1(n29393), .ZN(n1056) );
  I_NAND2 U1249 ( .A1(n1057), .B1(n29393), .ZN(n1058) );
  I_NAND2 U1250 ( .A1(n1059), .B1(n29393), .ZN(n1060) );
  I_NAND2 U1251 ( .A1(n1061), .B1(n29394), .ZN(n1062) );
  I_NAND2 U1252 ( .A1(n1063), .B1(n29394), .ZN(n1064) );
  I_NAND2 U1253 ( .A1(n1065), .B1(n29394), .ZN(n1066) );
  I_NAND2 U1254 ( .A1(n1067), .B1(n29394), .ZN(n1068) );
  I_NAND2 U1255 ( .A1(n1069), .B1(n29394), .ZN(n1070) );
  I_NAND2 U1256 ( .A1(n1071), .B1(n29394), .ZN(n1072) );
  I_NAND2 U1257 ( .A1(n1073), .B1(n29394), .ZN(n1074) );
  I_NAND2 U1258 ( .A1(n1075), .B1(n29394), .ZN(n1076) );
  I_NAND2 U1259 ( .A1(n1077), .B1(n29394), .ZN(n1078) );
  I_NAND2 U1260 ( .A1(n1079), .B1(n29394), .ZN(n1080) );
  I_NAND2 U1261 ( .A1(n1081), .B1(n29394), .ZN(n1082) );
  I_NAND2 U1262 ( .A1(n1083), .B1(n29394), .ZN(n1084) );
  I_NAND2 U1263 ( .A1(n1085), .B1(n29395), .ZN(n1086) );
  I_NAND2 U1264 ( .A1(n1087), .B1(n29395), .ZN(n1088) );
  I_NAND2 U1265 ( .A1(n1089), .B1(n29395), .ZN(n1090) );
  I_NAND2 U1266 ( .A1(n1091), .B1(n29395), .ZN(n1092) );
  I_NAND2 U1267 ( .A1(n1093), .B1(n29395), .ZN(n1094) );
  I_NAND2 U1268 ( .A1(n1095), .B1(n29395), .ZN(n1096) );
  I_NAND2 U1269 ( .A1(n1097), .B1(n29395), .ZN(n1098) );
  I_NAND2 U1270 ( .A1(n1099), .B1(n29395), .ZN(n1100) );
  I_NAND2 U1271 ( .A1(n1101), .B1(n29395), .ZN(n1102) );
  I_NAND2 U1272 ( .A1(n1103), .B1(n29395), .ZN(n1104) );
  I_NAND2 U1273 ( .A1(n1105), .B1(n29395), .ZN(n1106) );
  I_NAND2 U1274 ( .A1(n1107), .B1(n29395), .ZN(n1108) );
  I_NAND2 U1275 ( .A1(n1109), .B1(n29396), .ZN(n1110) );
  I_NAND2 U1276 ( .A1(n1111), .B1(n29396), .ZN(n1112) );
  I_NAND2 U1277 ( .A1(n1113), .B1(n29396), .ZN(n1114) );
  I_NAND2 U1278 ( .A1(n1115), .B1(n29396), .ZN(n1116) );
  I_NAND2 U1279 ( .A1(n1117), .B1(n29396), .ZN(n1118) );
  I_NAND2 U1280 ( .A1(n1119), .B1(n29396), .ZN(n1120) );
  I_NAND2 U1281 ( .A1(n1121), .B1(n29396), .ZN(n1122) );
  I_NAND2 U1282 ( .A1(n1126), .B1(n29396), .ZN(n1127) );
  I_NAND2 U1283 ( .A1(n1129), .B1(n29396), .ZN(n1130) );
  I_NAND2 U1284 ( .A1(n1131), .B1(n29396), .ZN(n1132) );
  I_NAND2 U1285 ( .A1(n1133), .B1(n29343), .ZN(n1134) );
  I_NAND2 U1286 ( .A1(n1135), .B1(n29338), .ZN(n1136) );
  I_NAND2 U1287 ( .A1(n1137), .B1(n29332), .ZN(n1138) );
  I_NAND2 U1288 ( .A1(n1139), .B1(n29332), .ZN(n1140) );
  I_NAND2 U1289 ( .A1(n1141), .B1(n29332), .ZN(n1142) );
  I_NAND2 U1290 ( .A1(n1143), .B1(n29333), .ZN(n1144) );
  I_NAND2 U1291 ( .A1(n1145), .B1(n29333), .ZN(n1146) );
  I_NAND2 U1292 ( .A1(n1147), .B1(n29333), .ZN(n1148) );
  I_NAND2 U1293 ( .A1(n1149), .B1(n29333), .ZN(n1150) );
  I_NAND2 U1294 ( .A1(n1151), .B1(n29333), .ZN(n1152) );
  I_NAND2 U1295 ( .A1(n1153), .B1(n29333), .ZN(n1154) );
  I_NAND2 U1296 ( .A1(n1155), .B1(n29333), .ZN(n1156) );
  I_NAND2 U1297 ( .A1(n1157), .B1(n29333), .ZN(n1158) );
  I_NAND2 U1298 ( .A1(n1159), .B1(n29333), .ZN(n1160) );
  I_NAND2 U1299 ( .A1(n1161), .B1(n29333), .ZN(n1162) );
  I_NAND2 U1300 ( .A1(n1163), .B1(n29333), .ZN(n1164) );
  I_NAND2 U1301 ( .A1(n1165), .B1(n29333), .ZN(n1166) );
  I_NAND2 U1302 ( .A1(n1167), .B1(n29334), .ZN(n1168) );
  I_NAND2 U1303 ( .A1(n1169), .B1(n29334), .ZN(n1170) );
  I_NAND2 U1304 ( .A1(n1171), .B1(n29334), .ZN(n1172) );
  I_NAND2 U1305 ( .A1(n1173), .B1(n29334), .ZN(n1174) );
  I_NAND2 U1306 ( .A1(n1175), .B1(n29334), .ZN(n1176) );
  I_NAND2 U1307 ( .A1(n1177), .B1(n29334), .ZN(n1178) );
  I_NAND2 U1308 ( .A1(n1179), .B1(n29334), .ZN(n1180) );
  I_NAND2 U1309 ( .A1(n1181), .B1(n29334), .ZN(n1182) );
  I_NAND2 U1310 ( .A1(n1183), .B1(n29334), .ZN(n1184) );
  I_NAND2 U1311 ( .A1(n1185), .B1(n29334), .ZN(n1186) );
  I_NAND2 U1312 ( .A1(n1187), .B1(n29334), .ZN(n1188) );
  I_NAND2 U1313 ( .A1(n1189), .B1(n29334), .ZN(n1190) );
  I_NAND2 U1314 ( .A1(n1191), .B1(n29335), .ZN(n1192) );
  I_NAND2 U1315 ( .A1(n1193), .B1(n29335), .ZN(n1194) );
  I_NAND2 U1316 ( .A1(n1195), .B1(n29335), .ZN(n1196) );
  I_NAND2 U1317 ( .A1(n1197), .B1(n29335), .ZN(n1198) );
  I_NAND2 U1318 ( .A1(n1199), .B1(n29335), .ZN(n1200) );
  I_NAND2 U1319 ( .A1(n1201), .B1(n29335), .ZN(n1202) );
  I_NAND2 U1320 ( .A1(n1203), .B1(n29335), .ZN(n1204) );
  I_NAND2 U1321 ( .A1(n1205), .B1(n29335), .ZN(n1206) );
  I_NAND2 U1322 ( .A1(n1207), .B1(n29335), .ZN(n1208) );
  I_NAND2 U1323 ( .A1(n1209), .B1(n29335), .ZN(n1210) );
  I_NAND2 U1324 ( .A1(n1211), .B1(n29335), .ZN(n1212) );
  I_NAND2 U1325 ( .A1(n1213), .B1(n29335), .ZN(n1214) );
  I_NAND2 U1326 ( .A1(n1215), .B1(n29336), .ZN(n1216) );
  I_NAND2 U1327 ( .A1(n1217), .B1(n29336), .ZN(n1218) );
  I_NAND2 U1328 ( .A1(n1219), .B1(n29336), .ZN(n1220) );
  I_NAND2 U1329 ( .A1(n1221), .B1(n29336), .ZN(n1222) );
  I_NAND2 U1330 ( .A1(n1223), .B1(n29336), .ZN(n1224) );
  I_NAND2 U1331 ( .A1(n1225), .B1(n29336), .ZN(n1226) );
  I_NAND2 U1332 ( .A1(n1227), .B1(n29336), .ZN(n1228) );
  I_NAND2 U1333 ( .A1(n1229), .B1(n29336), .ZN(n1230) );
  I_NAND2 U1334 ( .A1(n1231), .B1(n29336), .ZN(n1232) );
  I_NAND2 U1335 ( .A1(n1233), .B1(n29336), .ZN(n1234) );
  I_NAND2 U1336 ( .A1(n1235), .B1(n29336), .ZN(n1236) );
  I_NAND2 U1337 ( .A1(n1237), .B1(n29336), .ZN(n1238) );
  I_NAND2 U1338 ( .A1(n1239), .B1(n29337), .ZN(n1240) );
  I_NAND2 U1339 ( .A1(n1241), .B1(n29337), .ZN(n1242) );
  I_NAND2 U1340 ( .A1(n1243), .B1(n29337), .ZN(n1244) );
  I_NAND2 U1341 ( .A1(n1245), .B1(n29337), .ZN(n1246) );
  I_NAND2 U1342 ( .A1(n1247), .B1(n29337), .ZN(n1248) );
  I_NAND2 U1343 ( .A1(n1249), .B1(n29337), .ZN(n1250) );
  I_NAND2 U1344 ( .A1(n1251), .B1(n29337), .ZN(n1252) );
  I_NAND2 U1345 ( .A1(n1253), .B1(n29337), .ZN(n1254) );
  I_NAND2 U1346 ( .A1(n1256), .B1(n29337), .ZN(n1257) );
  I_NAND2 U1347 ( .A1(n1259), .B1(n29337), .ZN(n1260) );
  I_NAND2 U1348 ( .A1(n1261), .B1(n29337), .ZN(n1262) );
  I_NAND2 U1349 ( .A1(n1263), .B1(n29337), .ZN(n1264) );
  I_NAND2 U1350 ( .A1(n1265), .B1(n29338), .ZN(n1266) );
  I_NAND2 U1351 ( .A1(n1267), .B1(n29338), .ZN(n1268) );
  I_NAND2 U1352 ( .A1(n1269), .B1(n29338), .ZN(n1270) );
  I_NAND2 U1353 ( .A1(n1271), .B1(n29338), .ZN(n1272) );
  I_NAND2 U1354 ( .A1(n1273), .B1(n29338), .ZN(n1274) );
  I_NAND2 U1355 ( .A1(n1275), .B1(n29338), .ZN(n1276) );
  I_NAND2 U1356 ( .A1(n1277), .B1(n29338), .ZN(n1278) );
  I_NAND2 U1357 ( .A1(n1279), .B1(n29338), .ZN(n1280) );
  I_NAND2 U1358 ( .A1(n1281), .B1(n29338), .ZN(n1282) );
  I_NAND2 U1359 ( .A1(n1283), .B1(n29338), .ZN(n1284) );
  I_NAND2 U1360 ( .A1(n1285), .B1(n29338), .ZN(n1286) );
  I_NAND2 U1361 ( .A1(n1287), .B1(n29339), .ZN(n1288) );
  I_NAND2 U1362 ( .A1(n1289), .B1(n29339), .ZN(n1290) );
  I_NAND2 U1363 ( .A1(n1291), .B1(n29339), .ZN(n1292) );
  I_NAND2 U1364 ( .A1(n1293), .B1(n29339), .ZN(n1294) );
  I_NAND2 U1365 ( .A1(n1295), .B1(n29339), .ZN(n1296) );
  I_NAND2 U1366 ( .A1(n1297), .B1(n29339), .ZN(n1298) );
  I_NAND2 U1367 ( .A1(n1299), .B1(n29339), .ZN(n1300) );
  I_NAND2 U1368 ( .A1(n1301), .B1(n29339), .ZN(n1302) );
  I_NAND2 U1369 ( .A1(n1303), .B1(n29339), .ZN(n1304) );
  I_NAND2 U1370 ( .A1(n1305), .B1(n29339), .ZN(n1306) );
  I_NAND2 U1371 ( .A1(n1307), .B1(n29339), .ZN(n1308) );
  I_NAND2 U1372 ( .A1(n1309), .B1(n29339), .ZN(n1310) );
  I_NAND2 U1373 ( .A1(n1311), .B1(n29340), .ZN(n1312) );
  I_NAND2 U1374 ( .A1(n1313), .B1(n29340), .ZN(n1314) );
  I_NAND2 U1375 ( .A1(n1315), .B1(n29340), .ZN(n1316) );
  I_NAND2 U1376 ( .A1(n1317), .B1(n29340), .ZN(n1318) );
  I_NAND2 U1377 ( .A1(n1319), .B1(n29340), .ZN(n1320) );
  I_NAND2 U1378 ( .A1(n1321), .B1(n29340), .ZN(n1322) );
  I_NAND2 U1379 ( .A1(n1323), .B1(n29340), .ZN(n1324) );
  I_NAND2 U1380 ( .A1(n1325), .B1(n29340), .ZN(n1326) );
  I_NAND2 U1381 ( .A1(n1327), .B1(n29340), .ZN(n1328) );
  I_NAND2 U1382 ( .A1(n1329), .B1(n29340), .ZN(n1330) );
  I_NAND2 U1383 ( .A1(n1331), .B1(n29340), .ZN(n1332) );
  I_NAND2 U1384 ( .A1(n1333), .B1(n29340), .ZN(n1334) );
  I_NAND2 U1385 ( .A1(n1335), .B1(n29341), .ZN(n1336) );
  I_NAND2 U1386 ( .A1(n1337), .B1(n29341), .ZN(n1338) );
  I_NAND2 U1387 ( .A1(n1339), .B1(n29341), .ZN(n1340) );
  I_NAND2 U1388 ( .A1(n1341), .B1(n29341), .ZN(n1342) );
  I_NAND2 U1389 ( .A1(n1343), .B1(n29341), .ZN(n1344) );
  I_NAND2 U1390 ( .A1(n1345), .B1(n29341), .ZN(n1346) );
  I_NAND2 U1391 ( .A1(n1347), .B1(n29341), .ZN(n1348) );
  I_NAND2 U1392 ( .A1(n1349), .B1(n29341), .ZN(n1350) );
  I_NAND2 U1393 ( .A1(n1351), .B1(n29341), .ZN(n1352) );
  I_NAND2 U1394 ( .A1(n1353), .B1(n29341), .ZN(n1354) );
  I_NAND2 U1395 ( .A1(n1355), .B1(n29341), .ZN(n1356) );
  I_NAND2 U1396 ( .A1(n1357), .B1(n29341), .ZN(n1358) );
  I_NAND2 U1397 ( .A1(n1359), .B1(n29342), .ZN(n1360) );
  I_NAND2 U1398 ( .A1(n1361), .B1(n29342), .ZN(n1362) );
  I_NAND2 U1399 ( .A1(n1363), .B1(n29342), .ZN(n1364) );
  I_NAND2 U1400 ( .A1(n1365), .B1(n29342), .ZN(n1366) );
  I_NAND2 U1401 ( .A1(n1367), .B1(n29342), .ZN(n1368) );
  I_NAND2 U1402 ( .A1(n1369), .B1(n29342), .ZN(n1370) );
  I_NAND2 U1403 ( .A1(n1371), .B1(n29342), .ZN(n1372) );
  I_NAND2 U1404 ( .A1(n1373), .B1(n29342), .ZN(n1374) );
  I_NAND2 U1405 ( .A1(n1375), .B1(n29342), .ZN(n1376) );
  I_NAND2 U1406 ( .A1(n1377), .B1(n29342), .ZN(n1378) );
  I_NAND2 U1407 ( .A1(n1379), .B1(n29342), .ZN(n1380) );
  I_NAND2 U1408 ( .A1(n1381), .B1(n29342), .ZN(n1382) );
  I_NAND2 U1409 ( .A1(n1383), .B1(n29343), .ZN(n1384) );
  I_NAND2 U1410 ( .A1(n1385), .B1(n29343), .ZN(n1386) );
  I_NAND2 U1411 ( .A1(n1388), .B1(n29343), .ZN(n1389) );
  I_NAND2 U1412 ( .A1(n1390), .B1(n29343), .ZN(n1391) );
  I_NAND2 U1413 ( .A1(n1392), .B1(n29327), .ZN(n1393) );
  I_NAND2 U1414 ( .A1(n1394), .B1(n29322), .ZN(n1395) );
  I_NAND2 U1415 ( .A1(n1396), .B1(n29322), .ZN(n1397) );
  I_NAND2 U1416 ( .A1(n1398), .B1(n29322), .ZN(n1399) );
  I_NAND2 U1417 ( .A1(n1400), .B1(n29322), .ZN(n1401) );
  I_NAND2 U1418 ( .A1(n1402), .B1(n29322), .ZN(n1403) );
  I_NAND2 U1419 ( .A1(n1404), .B1(n29322), .ZN(n1405) );
  I_NAND2 U1420 ( .A1(n1406), .B1(n29322), .ZN(n1407) );
  I_NAND2 U1421 ( .A1(n1408), .B1(n29322), .ZN(n1409) );
  I_NAND2 U1422 ( .A1(n1410), .B1(n29322), .ZN(n1411) );
  I_NAND2 U1423 ( .A1(n1412), .B1(n29322), .ZN(n1413) );
  I_NAND2 U1424 ( .A1(n1414), .B1(n29322), .ZN(n1415) );
  I_NAND2 U1425 ( .A1(n1416), .B1(n29323), .ZN(n1417) );
  I_NAND2 U1426 ( .A1(n1418), .B1(n29323), .ZN(n1419) );
  I_NAND2 U1427 ( .A1(n1420), .B1(n29323), .ZN(n1421) );
  I_NAND2 U1428 ( .A1(n1422), .B1(n29323), .ZN(n1423) );
  I_NAND2 U1429 ( .A1(n1424), .B1(n29323), .ZN(n1425) );
  I_NAND2 U1430 ( .A1(n1426), .B1(n29323), .ZN(n1427) );
  I_NAND2 U1431 ( .A1(n1428), .B1(n29323), .ZN(n1429) );
  I_NAND2 U1432 ( .A1(n1430), .B1(n29323), .ZN(n1431) );
  I_NAND2 U1433 ( .A1(n1432), .B1(n29323), .ZN(n1433) );
  I_NAND2 U1434 ( .A1(n1434), .B1(n29323), .ZN(n1435) );
  I_NAND2 U1435 ( .A1(n1436), .B1(n29323), .ZN(n1437) );
  I_NAND2 U1436 ( .A1(n1438), .B1(n29323), .ZN(n1439) );
  I_NAND2 U1437 ( .A1(n1440), .B1(n29324), .ZN(n1441) );
  I_NAND2 U1438 ( .A1(n1442), .B1(n29324), .ZN(n1443) );
  I_NAND2 U1439 ( .A1(n1444), .B1(n29324), .ZN(n1445) );
  I_NAND2 U1440 ( .A1(n1446), .B1(n29324), .ZN(n1447) );
  I_NAND2 U1441 ( .A1(n1448), .B1(n29324), .ZN(n1449) );
  I_NAND2 U1442 ( .A1(n1450), .B1(n29324), .ZN(n1451) );
  I_NAND2 U1443 ( .A1(n1452), .B1(n29324), .ZN(n1453) );
  I_NAND2 U1444 ( .A1(n1454), .B1(n29324), .ZN(n1455) );
  I_NAND2 U1445 ( .A1(n1456), .B1(n29324), .ZN(n1457) );
  I_NAND2 U1446 ( .A1(n1458), .B1(n29324), .ZN(n1459) );
  I_NAND2 U1447 ( .A1(n1460), .B1(n29324), .ZN(n1461) );
  I_NAND2 U1448 ( .A1(n1462), .B1(n29324), .ZN(n1463) );
  I_NAND2 U1449 ( .A1(n1464), .B1(n29325), .ZN(n1465) );
  I_NAND2 U1450 ( .A1(n1466), .B1(n29325), .ZN(n1467) );
  I_NAND2 U1451 ( .A1(n1468), .B1(n29325), .ZN(n1469) );
  I_NAND2 U1452 ( .A1(n1470), .B1(n29325), .ZN(n1471) );
  I_NAND2 U1453 ( .A1(n1472), .B1(n29325), .ZN(n1473) );
  I_NAND2 U1454 ( .A1(n1474), .B1(n29325), .ZN(n1475) );
  I_NAND2 U1455 ( .A1(n1476), .B1(n29325), .ZN(n1477) );
  I_NAND2 U1456 ( .A1(n1478), .B1(n29325), .ZN(n1479) );
  I_NAND2 U1457 ( .A1(n1480), .B1(n29325), .ZN(n1481) );
  I_NAND2 U1458 ( .A1(n1482), .B1(n29325), .ZN(n1483) );
  I_NAND2 U1459 ( .A1(n1484), .B1(n29325), .ZN(n1485) );
  I_NAND2 U1460 ( .A1(n1486), .B1(n29325), .ZN(n1487) );
  I_NAND2 U1461 ( .A1(n1488), .B1(n29326), .ZN(n1489) );
  I_NAND2 U1462 ( .A1(n1490), .B1(n29326), .ZN(n1491) );
  I_NAND2 U1463 ( .A1(n1492), .B1(n29326), .ZN(n1493) );
  I_NAND2 U1464 ( .A1(n1494), .B1(n29326), .ZN(n1495) );
  I_NAND2 U1465 ( .A1(n1496), .B1(n29326), .ZN(n1497) );
  I_NAND2 U1466 ( .A1(n1498), .B1(n29326), .ZN(n1499) );
  I_NAND2 U1467 ( .A1(n1500), .B1(n29326), .ZN(n1501) );
  I_NAND2 U1468 ( .A1(n1502), .B1(n29326), .ZN(n1503) );
  I_NAND2 U1469 ( .A1(n1504), .B1(n29326), .ZN(n1505) );
  I_NAND2 U1470 ( .A1(n1506), .B1(n29326), .ZN(n1507) );
  I_NAND2 U1471 ( .A1(n1508), .B1(n29326), .ZN(n1509) );
  I_NAND2 U1472 ( .A1(n1510), .B1(n29326), .ZN(n1511) );
  I_NAND2 U1473 ( .A1(n1512), .B1(n29327), .ZN(n1513) );
  I_NAND2 U1474 ( .A1(n1514), .B1(n29327), .ZN(n1515) );
  I_NAND2 U1475 ( .A1(n1517), .B1(n29327), .ZN(n1518) );
  I_NAND2 U1476 ( .A1(n1519), .B1(n29327), .ZN(n1520) );
  I_NAND2 U1477 ( .A1(n1521), .B1(n29327), .ZN(n1522) );
  I_NAND2 U1478 ( .A1(n1523), .B1(n29327), .ZN(n1524) );
  I_NAND2 U1479 ( .A1(n1525), .B1(n29327), .ZN(n1526) );
  I_NAND2 U1480 ( .A1(n1527), .B1(n29327), .ZN(n1528) );
  I_NAND2 U1481 ( .A1(n1529), .B1(n29327), .ZN(n1530) );
  I_NAND2 U1482 ( .A1(n1531), .B1(n29327), .ZN(n1532) );
  I_NAND2 U1483 ( .A1(n1533), .B1(n29327), .ZN(n1534) );
  I_NAND2 U1484 ( .A1(n1535), .B1(n29328), .ZN(n1536) );
  I_NAND2 U1485 ( .A1(n1537), .B1(n29328), .ZN(n1538) );
  I_NAND2 U1486 ( .A1(n1539), .B1(n29328), .ZN(n1540) );
  I_NAND2 U1487 ( .A1(n1541), .B1(n29328), .ZN(n1542) );
  I_NAND2 U1488 ( .A1(n1543), .B1(n29328), .ZN(n1544) );
  I_NAND2 U1489 ( .A1(n1545), .B1(n29328), .ZN(n1546) );
  I_NAND2 U1490 ( .A1(n1547), .B1(n29328), .ZN(n1548) );
  I_NAND2 U1491 ( .A1(n1549), .B1(n29328), .ZN(n1550) );
  I_NAND2 U1492 ( .A1(n1551), .B1(n29328), .ZN(n1552) );
  I_NAND2 U1493 ( .A1(n1553), .B1(n29328), .ZN(n1554) );
  I_NAND2 U1494 ( .A1(n1555), .B1(n29328), .ZN(n1556) );
  I_NAND2 U1495 ( .A1(n1557), .B1(n29328), .ZN(n1558) );
  I_NAND2 U1496 ( .A1(n1559), .B1(n29329), .ZN(n1560) );
  I_NAND2 U1497 ( .A1(n1561), .B1(n29329), .ZN(n1562) );
  I_NAND2 U1498 ( .A1(n1563), .B1(n29329), .ZN(n1564) );
  I_NAND2 U1499 ( .A1(n1565), .B1(n29329), .ZN(n1566) );
  I_NAND2 U1500 ( .A1(n1567), .B1(n29329), .ZN(n1568) );
  I_NAND2 U1501 ( .A1(n1569), .B1(n29329), .ZN(n1570) );
  I_NAND2 U1502 ( .A1(n1571), .B1(n29329), .ZN(n1572) );
  I_NAND2 U1503 ( .A1(n1573), .B1(n29329), .ZN(n1574) );
  I_NAND2 U1504 ( .A1(n1575), .B1(n29329), .ZN(n1576) );
  I_NAND2 U1505 ( .A1(n1577), .B1(n29329), .ZN(n1578) );
  I_NAND2 U1506 ( .A1(n1579), .B1(n29329), .ZN(n1580) );
  I_NAND2 U1507 ( .A1(n1581), .B1(n29329), .ZN(n1582) );
  I_NAND2 U1508 ( .A1(n1583), .B1(n29330), .ZN(n1584) );
  I_NAND2 U1509 ( .A1(n1585), .B1(n29330), .ZN(n1586) );
  I_NAND2 U1510 ( .A1(n1587), .B1(n29330), .ZN(n1588) );
  I_NAND2 U1511 ( .A1(n1589), .B1(n29330), .ZN(n1590) );
  I_NAND2 U1512 ( .A1(n1591), .B1(n29330), .ZN(n1592) );
  I_NAND2 U1513 ( .A1(n1593), .B1(n29330), .ZN(n1594) );
  I_NAND2 U1514 ( .A1(n1595), .B1(n29330), .ZN(n1596) );
  I_NAND2 U1515 ( .A1(n1597), .B1(n29330), .ZN(n1598) );
  I_NAND2 U1516 ( .A1(n1599), .B1(n29330), .ZN(n1600) );
  I_NAND2 U1517 ( .A1(n1601), .B1(n29330), .ZN(n1602) );
  I_NAND2 U1518 ( .A1(n1603), .B1(n29330), .ZN(n1604) );
  I_NAND2 U1519 ( .A1(n1605), .B1(n29330), .ZN(n1606) );
  I_NAND2 U1520 ( .A1(n1607), .B1(n29331), .ZN(n1608) );
  I_NAND2 U1521 ( .A1(n1609), .B1(n29331), .ZN(n1610) );
  I_NAND2 U1522 ( .A1(n1611), .B1(n29331), .ZN(n1612) );
  I_NAND2 U1523 ( .A1(n1613), .B1(n29331), .ZN(n1614) );
  I_NAND2 U1524 ( .A1(n1615), .B1(n29331), .ZN(n1616) );
  I_NAND2 U1525 ( .A1(n1617), .B1(n29331), .ZN(n1618) );
  I_NAND2 U1526 ( .A1(n1619), .B1(n29331), .ZN(n1620) );
  I_NAND2 U1527 ( .A1(n1621), .B1(n29331), .ZN(n1622) );
  I_NAND2 U1528 ( .A1(n1623), .B1(n29331), .ZN(n1624) );
  I_NAND2 U1529 ( .A1(n1625), .B1(n29331), .ZN(n1626) );
  I_NAND2 U1530 ( .A1(n1627), .B1(n29331), .ZN(n1628) );
  I_NAND2 U1531 ( .A1(n1629), .B1(n29331), .ZN(n1630) );
  I_NAND2 U1532 ( .A1(n1631), .B1(n29332), .ZN(n1632) );
  I_NAND2 U1533 ( .A1(n1633), .B1(n29332), .ZN(n1634) );
  I_NAND2 U1534 ( .A1(n1635), .B1(n29332), .ZN(n1636) );
  I_NAND2 U1535 ( .A1(n1637), .B1(n29332), .ZN(n1638) );
  I_NAND2 U1536 ( .A1(n1639), .B1(n29332), .ZN(n1640) );
  I_NAND2 U1537 ( .A1(n1641), .B1(n29332), .ZN(n1642) );
  I_NAND2 U1538 ( .A1(n1643), .B1(n29332), .ZN(n1644) );
  I_NAND2 U1539 ( .A1(n1646), .B1(n29332), .ZN(n1647) );
  I_NAND2 U1540 ( .A1(n1648), .B1(n29332), .ZN(n1649) );
  I_NAND2 U1541 ( .A1(n1650), .B1(n29359), .ZN(n1651) );
  I_NAND2 U1542 ( .A1(n1652), .B1(n29354), .ZN(n1653) );
  I_NAND2 U1543 ( .A1(n1654), .B1(n29354), .ZN(n1655) );
  I_NAND2 U1544 ( .A1(n1656), .B1(n29354), .ZN(n1657) );
  I_NAND2 U1545 ( .A1(n1658), .B1(n29354), .ZN(n1659) );
  I_NAND2 U1546 ( .A1(n1660), .B1(n29354), .ZN(n1661) );
  I_NAND2 U1547 ( .A1(n1662), .B1(n29354), .ZN(n1663) );
  I_NAND2 U1548 ( .A1(n1664), .B1(n29354), .ZN(n1665) );
  I_NAND2 U1549 ( .A1(n1666), .B1(n29354), .ZN(n1667) );
  I_NAND2 U1550 ( .A1(n1668), .B1(n29354), .ZN(n1669) );
  I_NAND2 U1551 ( .A1(n1670), .B1(n29354), .ZN(n1671) );
  I_NAND2 U1552 ( .A1(n1672), .B1(n29354), .ZN(n1673) );
  I_NAND2 U1553 ( .A1(n1674), .B1(n29355), .ZN(n1675) );
  I_NAND2 U1554 ( .A1(n1676), .B1(n29355), .ZN(n1677) );
  I_NAND2 U1555 ( .A1(n1678), .B1(n29355), .ZN(n1679) );
  I_NAND2 U1556 ( .A1(n1680), .B1(n29355), .ZN(n1681) );
  I_NAND2 U1557 ( .A1(n1682), .B1(n29355), .ZN(n1683) );
  I_NAND2 U1558 ( .A1(n1684), .B1(n29355), .ZN(n1685) );
  I_NAND2 U1559 ( .A1(n1686), .B1(n29355), .ZN(n1687) );
  I_NAND2 U1560 ( .A1(n1688), .B1(n29355), .ZN(n1689) );
  I_NAND2 U1561 ( .A1(n1690), .B1(n29355), .ZN(n1691) );
  I_NAND2 U1562 ( .A1(n1692), .B1(n29355), .ZN(n1693) );
  I_NAND2 U1563 ( .A1(n1694), .B1(n29355), .ZN(n1695) );
  I_NAND2 U1564 ( .A1(n1696), .B1(n29355), .ZN(n1697) );
  I_NAND2 U1565 ( .A1(n1698), .B1(n29356), .ZN(n1699) );
  I_NAND2 U1566 ( .A1(n1700), .B1(n29356), .ZN(n1701) );
  I_NAND2 U1567 ( .A1(n1702), .B1(n29356), .ZN(n1703) );
  I_NAND2 U1568 ( .A1(n1704), .B1(n29356), .ZN(n1705) );
  I_NAND2 U1569 ( .A1(n1706), .B1(n29356), .ZN(n1707) );
  I_NAND2 U1570 ( .A1(n1708), .B1(n29356), .ZN(n1709) );
  I_NAND2 U1571 ( .A1(n1710), .B1(n29356), .ZN(n1711) );
  I_NAND2 U1572 ( .A1(n1712), .B1(n29356), .ZN(n1713) );
  I_NAND2 U1573 ( .A1(n1714), .B1(n29356), .ZN(n1715) );
  I_NAND2 U1574 ( .A1(n1716), .B1(n29356), .ZN(n1717) );
  I_NAND2 U1575 ( .A1(n1718), .B1(n29356), .ZN(n1719) );
  I_NAND2 U1576 ( .A1(n1720), .B1(n29356), .ZN(n1721) );
  I_NAND2 U1577 ( .A1(n1722), .B1(n29357), .ZN(n1723) );
  I_NAND2 U1578 ( .A1(n1724), .B1(n29357), .ZN(n1725) );
  I_NAND2 U1579 ( .A1(n1726), .B1(n29357), .ZN(n1727) );
  I_NAND2 U1580 ( .A1(n1728), .B1(n29357), .ZN(n1729) );
  I_NAND2 U1581 ( .A1(n1730), .B1(n29357), .ZN(n1731) );
  I_NAND2 U1582 ( .A1(n1732), .B1(n29357), .ZN(n1733) );
  I_NAND2 U1583 ( .A1(n1734), .B1(n29357), .ZN(n1735) );
  I_NAND2 U1584 ( .A1(n1736), .B1(n29357), .ZN(n1737) );
  I_NAND2 U1585 ( .A1(n1738), .B1(n29357), .ZN(n1739) );
  I_NAND2 U1586 ( .A1(n1740), .B1(n29357), .ZN(n1741) );
  I_NAND2 U1587 ( .A1(n1742), .B1(n29357), .ZN(n1743) );
  I_NAND2 U1588 ( .A1(n1744), .B1(n29357), .ZN(n1745) );
  I_NAND2 U1589 ( .A1(n1746), .B1(n29358), .ZN(n1747) );
  I_NAND2 U1590 ( .A1(n1748), .B1(n29358), .ZN(n1749) );
  I_NAND2 U1591 ( .A1(n1750), .B1(n29358), .ZN(n1751) );
  I_NAND2 U1592 ( .A1(n1752), .B1(n29358), .ZN(n1753) );
  I_NAND2 U1593 ( .A1(n1754), .B1(n29358), .ZN(n1755) );
  I_NAND2 U1594 ( .A1(n1756), .B1(n29358), .ZN(n1757) );
  I_NAND2 U1595 ( .A1(n1758), .B1(n29358), .ZN(n1759) );
  I_NAND2 U1596 ( .A1(n1760), .B1(n29358), .ZN(n1761) );
  I_NAND2 U1597 ( .A1(n1762), .B1(n29358), .ZN(n1763) );
  I_NAND2 U1598 ( .A1(n1764), .B1(n29358), .ZN(n1765) );
  I_NAND2 U1599 ( .A1(n1766), .B1(n29358), .ZN(n1767) );
  I_NAND2 U1600 ( .A1(n1768), .B1(n29358), .ZN(n1769) );
  I_NAND2 U1601 ( .A1(n1770), .B1(n29359), .ZN(n1771) );
  I_NAND2 U1602 ( .A1(n1772), .B1(n29359), .ZN(n1773) );
  I_NAND2 U1603 ( .A1(n1775), .B1(n29359), .ZN(n1776) );
  I_NAND2 U1604 ( .A1(n1777), .B1(n29359), .ZN(n1778) );
  I_NAND2 U1605 ( .A1(n1779), .B1(n29359), .ZN(n1780) );
  I_NAND2 U1606 ( .A1(n1781), .B1(n29359), .ZN(n1782) );
  I_NAND2 U1607 ( .A1(n1783), .B1(n29359), .ZN(n1784) );
  I_NAND2 U1608 ( .A1(n1785), .B1(n29359), .ZN(n1786) );
  I_NAND2 U1609 ( .A1(n1787), .B1(n29359), .ZN(n1788) );
  I_NAND2 U1610 ( .A1(n1789), .B1(n29359), .ZN(n1790) );
  I_NAND2 U1611 ( .A1(n1791), .B1(n29359), .ZN(n1792) );
  I_NAND2 U1612 ( .A1(n1793), .B1(n29360), .ZN(n1794) );
  I_NAND2 U1613 ( .A1(n1795), .B1(n29360), .ZN(n1796) );
  I_NAND2 U1614 ( .A1(n1797), .B1(n29360), .ZN(n1798) );
  I_NAND2 U1615 ( .A1(n1799), .B1(n29360), .ZN(n1800) );
  I_NAND2 U1616 ( .A1(n1801), .B1(n29360), .ZN(n1802) );
  I_NAND2 U1617 ( .A1(n1803), .B1(n29360), .ZN(n1804) );
  I_NAND2 U1618 ( .A1(n1805), .B1(n29360), .ZN(n1806) );
  I_NAND2 U1619 ( .A1(n1807), .B1(n29360), .ZN(n1808) );
  I_NAND2 U1620 ( .A1(n1809), .B1(n29360), .ZN(n1810) );
  I_NAND2 U1621 ( .A1(n1811), .B1(n29360), .ZN(n1812) );
  I_NAND2 U1622 ( .A1(n1813), .B1(n29360), .ZN(n1814) );
  I_NAND2 U1623 ( .A1(n1815), .B1(n29360), .ZN(n1816) );
  I_NAND2 U1624 ( .A1(n1817), .B1(n29361), .ZN(n1818) );
  I_NAND2 U1625 ( .A1(n1819), .B1(n29361), .ZN(n1820) );
  I_NAND2 U1626 ( .A1(n1821), .B1(n29361), .ZN(n1822) );
  I_NAND2 U1627 ( .A1(n1823), .B1(n29361), .ZN(n1824) );
  I_NAND2 U1628 ( .A1(n1825), .B1(n29361), .ZN(n1826) );
  I_NAND2 U1629 ( .A1(n1827), .B1(n29361), .ZN(n1828) );
  I_NAND2 U1630 ( .A1(n1829), .B1(n29361), .ZN(n1830) );
  I_NAND2 U1631 ( .A1(n1831), .B1(n29361), .ZN(n1832) );
  I_NAND2 U1632 ( .A1(n1833), .B1(n29361), .ZN(n1834) );
  I_NAND2 U1633 ( .A1(n1835), .B1(n29361), .ZN(n1836) );
  I_NAND2 U1634 ( .A1(n1837), .B1(n29361), .ZN(n1838) );
  I_NAND2 U1635 ( .A1(n1839), .B1(n29361), .ZN(n1840) );
  I_NAND2 U1636 ( .A1(n1841), .B1(n29362), .ZN(n1842) );
  I_NAND2 U1637 ( .A1(n1843), .B1(n29362), .ZN(n1844) );
  I_NAND2 U1638 ( .A1(n1845), .B1(n29362), .ZN(n1846) );
  I_NAND2 U1639 ( .A1(n1847), .B1(n29362), .ZN(n1848) );
  I_NAND2 U1640 ( .A1(n1849), .B1(n29362), .ZN(n1850) );
  I_NAND2 U1641 ( .A1(n1851), .B1(n29362), .ZN(n1852) );
  I_NAND2 U1642 ( .A1(n1853), .B1(n29362), .ZN(n1854) );
  I_NAND2 U1643 ( .A1(n1855), .B1(n29362), .ZN(n1856) );
  I_NAND2 U1644 ( .A1(n1857), .B1(n29362), .ZN(n1858) );
  I_NAND2 U1645 ( .A1(n1859), .B1(n29362), .ZN(n1860) );
  I_NAND2 U1646 ( .A1(n1861), .B1(n29362), .ZN(n1862) );
  I_NAND2 U1647 ( .A1(n1863), .B1(n29362), .ZN(n1864) );
  I_NAND2 U1648 ( .A1(n1865), .B1(n29363), .ZN(n1866) );
  I_NAND2 U1649 ( .A1(n1867), .B1(n29363), .ZN(n1868) );
  I_NAND2 U1650 ( .A1(n1869), .B1(n29363), .ZN(n1870) );
  I_NAND2 U1651 ( .A1(n1871), .B1(n29363), .ZN(n1872) );
  I_NAND2 U1652 ( .A1(n1873), .B1(n29363), .ZN(n1874) );
  I_NAND2 U1653 ( .A1(n1875), .B1(n29363), .ZN(n1876) );
  I_NAND2 U1654 ( .A1(n1877), .B1(n29363), .ZN(n1878) );
  I_NAND2 U1655 ( .A1(n1879), .B1(n29363), .ZN(n1880) );
  I_NAND2 U1656 ( .A1(n1881), .B1(n29363), .ZN(n1882) );
  I_NAND2 U1657 ( .A1(n1883), .B1(n29363), .ZN(n1884) );
  I_NAND2 U1658 ( .A1(n1885), .B1(n29363), .ZN(n1886) );
  I_NAND2 U1659 ( .A1(n1887), .B1(n29363), .ZN(n1888) );
  I_NAND2 U1660 ( .A1(n1889), .B1(n29364), .ZN(n1890) );
  I_NAND2 U1661 ( .A1(n1891), .B1(n29364), .ZN(n1892) );
  I_NAND2 U1662 ( .A1(n1893), .B1(n29364), .ZN(n1894) );
  I_NAND2 U1663 ( .A1(n1895), .B1(n29364), .ZN(n1896) );
  I_NAND2 U1664 ( .A1(n1897), .B1(n29364), .ZN(n1898) );
  I_NAND2 U1665 ( .A1(n1899), .B1(n29364), .ZN(n1900) );
  I_NAND2 U1666 ( .A1(n1901), .B1(n29364), .ZN(n1902) );
  I_NAND2 U1667 ( .A1(n1904), .B1(n29364), .ZN(n1905) );
  I_NAND2 U1668 ( .A1(n1906), .B1(n29364), .ZN(n1907) );
  I_NAND2 U1669 ( .A1(n1908), .B1(n29348), .ZN(n1909) );
  I_NAND2 U1670 ( .A1(n1910), .B1(n29343), .ZN(n1911) );
  I_NAND2 U1671 ( .A1(n1912), .B1(n29343), .ZN(n1913) );
  I_NAND2 U1672 ( .A1(n1914), .B1(n29343), .ZN(n1915) );
  I_NAND2 U1673 ( .A1(n1916), .B1(n29343), .ZN(n1917) );
  I_NAND2 U1674 ( .A1(n1918), .B1(n29343), .ZN(n1919) );
  I_NAND2 U1675 ( .A1(n1920), .B1(n29343), .ZN(n1921) );
  I_NAND2 U1676 ( .A1(n1922), .B1(n29343), .ZN(n1923) );
  I_NAND2 U1677 ( .A1(n1924), .B1(n29344), .ZN(n1925) );
  I_NAND2 U1678 ( .A1(n1926), .B1(n29344), .ZN(n1927) );
  I_NAND2 U1679 ( .A1(n1928), .B1(n29344), .ZN(n1929) );
  I_NAND2 U1680 ( .A1(n1930), .B1(n29344), .ZN(n1931) );
  I_NAND2 U1681 ( .A1(n1932), .B1(n29344), .ZN(n1933) );
  I_NAND2 U1682 ( .A1(n1934), .B1(n29344), .ZN(n1935) );
  I_NAND2 U1683 ( .A1(n1936), .B1(n29344), .ZN(n1937) );
  I_NAND2 U1684 ( .A1(n1938), .B1(n29344), .ZN(n1939) );
  I_NAND2 U1685 ( .A1(n1940), .B1(n29344), .ZN(n1941) );
  I_NAND2 U1686 ( .A1(n1942), .B1(n29344), .ZN(n1943) );
  I_NAND2 U1687 ( .A1(n1944), .B1(n29344), .ZN(n1945) );
  I_NAND2 U1688 ( .A1(n1946), .B1(n29344), .ZN(n1947) );
  I_NAND2 U1689 ( .A1(n1948), .B1(n29345), .ZN(n1949) );
  I_NAND2 U1690 ( .A1(n1950), .B1(n29345), .ZN(n1951) );
  I_NAND2 U1691 ( .A1(n1952), .B1(n29345), .ZN(n1953) );
  I_NAND2 U1692 ( .A1(n1954), .B1(n29345), .ZN(n1955) );
  I_NAND2 U1693 ( .A1(n1956), .B1(n29345), .ZN(n1957) );
  I_NAND2 U1694 ( .A1(n1958), .B1(n29345), .ZN(n1959) );
  I_NAND2 U1695 ( .A1(n1960), .B1(n29345), .ZN(n1961) );
  I_NAND2 U1696 ( .A1(n1962), .B1(n29345), .ZN(n1963) );
  I_NAND2 U1697 ( .A1(n1964), .B1(n29345), .ZN(n1965) );
  I_NAND2 U1698 ( .A1(n1966), .B1(n29345), .ZN(n1967) );
  I_NAND2 U1699 ( .A1(n1968), .B1(n29345), .ZN(n1969) );
  I_NAND2 U1700 ( .A1(n1970), .B1(n29345), .ZN(n1971) );
  I_NAND2 U1701 ( .A1(n1972), .B1(n29346), .ZN(n1973) );
  I_NAND2 U1702 ( .A1(n1974), .B1(n29346), .ZN(n1975) );
  I_NAND2 U1703 ( .A1(n1976), .B1(n29346), .ZN(n1977) );
  I_NAND2 U1704 ( .A1(n1978), .B1(n29346), .ZN(n1979) );
  I_NAND2 U1705 ( .A1(n1980), .B1(n29346), .ZN(n1981) );
  I_NAND2 U1706 ( .A1(n1982), .B1(n29346), .ZN(n1983) );
  I_NAND2 U1707 ( .A1(n1984), .B1(n29346), .ZN(n1985) );
  I_NAND2 U1708 ( .A1(n1986), .B1(n29346), .ZN(n1987) );
  I_NAND2 U1709 ( .A1(n1988), .B1(n29346), .ZN(n1989) );
  I_NAND2 U1710 ( .A1(n1990), .B1(n29346), .ZN(n1991) );
  I_NAND2 U1711 ( .A1(n1992), .B1(n29346), .ZN(n1993) );
  I_NAND2 U1712 ( .A1(n1994), .B1(n29346), .ZN(n1995) );
  I_NAND2 U1713 ( .A1(n1996), .B1(n29347), .ZN(n1997) );
  I_NAND2 U1714 ( .A1(n1998), .B1(n29347), .ZN(n1999) );
  I_NAND2 U1715 ( .A1(n2000), .B1(n29347), .ZN(n2001) );
  I_NAND2 U1716 ( .A1(n2002), .B1(n29347), .ZN(n2003) );
  I_NAND2 U1717 ( .A1(n2004), .B1(n29347), .ZN(n2005) );
  I_NAND2 U1718 ( .A1(n2006), .B1(n29347), .ZN(n2007) );
  I_NAND2 U1719 ( .A1(n2008), .B1(n29347), .ZN(n2009) );
  I_NAND2 U1720 ( .A1(n2010), .B1(n29347), .ZN(n2011) );
  I_NAND2 U1721 ( .A1(n2012), .B1(n29347), .ZN(n2013) );
  I_NAND2 U1722 ( .A1(n2014), .B1(n29347), .ZN(n2015) );
  I_NAND2 U1723 ( .A1(n2016), .B1(n29347), .ZN(n2017) );
  I_NAND2 U1724 ( .A1(n2018), .B1(n29347), .ZN(n2019) );
  I_NAND2 U1725 ( .A1(n2020), .B1(n29348), .ZN(n2021) );
  I_NAND2 U1726 ( .A1(n2022), .B1(n29348), .ZN(n2023) );
  I_NAND2 U1727 ( .A1(n2024), .B1(n29348), .ZN(n2025) );
  I_NAND2 U1728 ( .A1(n2026), .B1(n29348), .ZN(n2027) );
  I_NAND2 U1729 ( .A1(n2028), .B1(n29348), .ZN(n2029) );
  I_NAND2 U1730 ( .A1(n2030), .B1(n29348), .ZN(n2031) );
  I_NAND2 U1731 ( .A1(n2033), .B1(n29348), .ZN(n2034) );
  I_NAND2 U1732 ( .A1(n2035), .B1(n29348), .ZN(n2036) );
  I_NAND2 U1733 ( .A1(n2037), .B1(n29348), .ZN(n2038) );
  I_NAND2 U1734 ( .A1(n2039), .B1(n29348), .ZN(n2040) );
  I_NAND2 U1735 ( .A1(n2041), .B1(n29348), .ZN(n2042) );
  I_NAND2 U1736 ( .A1(n2043), .B1(n29349), .ZN(n2044) );
  I_NAND2 U1737 ( .A1(n2045), .B1(n29349), .ZN(n2046) );
  I_NAND2 U1738 ( .A1(n2047), .B1(n29349), .ZN(n2048) );
  I_NAND2 U1739 ( .A1(n2049), .B1(n29349), .ZN(n2050) );
  I_NAND2 U1740 ( .A1(n2051), .B1(n29349), .ZN(n2052) );
  I_NAND2 U1741 ( .A1(n2053), .B1(n29349), .ZN(n2054) );
  I_NAND2 U1742 ( .A1(n2055), .B1(n29349), .ZN(n2056) );
  I_NAND2 U1743 ( .A1(n2057), .B1(n29349), .ZN(n2058) );
  I_NAND2 U1744 ( .A1(n2059), .B1(n29349), .ZN(n2060) );
  I_NAND2 U1745 ( .A1(n2061), .B1(n29349), .ZN(n2062) );
  I_NAND2 U1746 ( .A1(n2063), .B1(n29349), .ZN(n2064) );
  I_NAND2 U1747 ( .A1(n2065), .B1(n29349), .ZN(n2066) );
  I_NAND2 U1748 ( .A1(n2067), .B1(n29350), .ZN(n2068) );
  I_NAND2 U1749 ( .A1(n2069), .B1(n29350), .ZN(n2070) );
  I_NAND2 U1750 ( .A1(n2071), .B1(n29350), .ZN(n2072) );
  I_NAND2 U1751 ( .A1(n2073), .B1(n29350), .ZN(n2074) );
  I_NAND2 U1752 ( .A1(n2075), .B1(n29350), .ZN(n2076) );
  I_NAND2 U1753 ( .A1(n2077), .B1(n29350), .ZN(n2078) );
  I_NAND2 U1754 ( .A1(n2079), .B1(n29350), .ZN(n2080) );
  I_NAND2 U1755 ( .A1(n2081), .B1(n29350), .ZN(n2082) );
  I_NAND2 U1756 ( .A1(n2083), .B1(n29350), .ZN(n2084) );
  I_NAND2 U1757 ( .A1(n2085), .B1(n29350), .ZN(n2086) );
  I_NAND2 U1758 ( .A1(n2087), .B1(n29350), .ZN(n2088) );
  I_NAND2 U1759 ( .A1(n2089), .B1(n29350), .ZN(n2090) );
  I_NAND2 U1760 ( .A1(n2091), .B1(n29351), .ZN(n2092) );
  I_NAND2 U1761 ( .A1(n2093), .B1(n29351), .ZN(n2094) );
  I_NAND2 U1762 ( .A1(n2095), .B1(n29351), .ZN(n2096) );
  I_NAND2 U1763 ( .A1(n2097), .B1(n29351), .ZN(n2098) );
  I_NAND2 U1764 ( .A1(n2099), .B1(n29351), .ZN(n2100) );
  I_NAND2 U1765 ( .A1(n2101), .B1(n29351), .ZN(n2102) );
  I_NAND2 U1766 ( .A1(n2103), .B1(n29351), .ZN(n2104) );
  I_NAND2 U1767 ( .A1(n2105), .B1(n29351), .ZN(n2106) );
  I_NAND2 U1768 ( .A1(n2107), .B1(n29351), .ZN(n2108) );
  I_NAND2 U1769 ( .A1(n2109), .B1(n29351), .ZN(n2110) );
  I_NAND2 U1770 ( .A1(n2111), .B1(n29351), .ZN(n2112) );
  I_NAND2 U1771 ( .A1(n2113), .B1(n29351), .ZN(n2114) );
  I_NAND2 U1772 ( .A1(n2115), .B1(n29352), .ZN(n2116) );
  I_NAND2 U1773 ( .A1(n2117), .B1(n29352), .ZN(n2118) );
  I_NAND2 U1774 ( .A1(n2119), .B1(n29352), .ZN(n2120) );
  I_NAND2 U1775 ( .A1(n2121), .B1(n29352), .ZN(n2122) );
  I_NAND2 U1776 ( .A1(n2123), .B1(n29352), .ZN(n2124) );
  I_NAND2 U1777 ( .A1(n2125), .B1(n29352), .ZN(n2126) );
  I_NAND2 U1778 ( .A1(n2127), .B1(n29352), .ZN(n2128) );
  I_NAND2 U1779 ( .A1(n2129), .B1(n29352), .ZN(n2130) );
  I_NAND2 U1780 ( .A1(n2131), .B1(n29352), .ZN(n2132) );
  I_NAND2 U1781 ( .A1(n2133), .B1(n29352), .ZN(n2134) );
  I_NAND2 U1782 ( .A1(n2135), .B1(n29352), .ZN(n2136) );
  I_NAND2 U1783 ( .A1(n2137), .B1(n29352), .ZN(n2138) );
  I_NAND2 U1784 ( .A1(n2139), .B1(n29353), .ZN(n2140) );
  I_NAND2 U1785 ( .A1(n2141), .B1(n29353), .ZN(n2142) );
  I_NAND2 U1786 ( .A1(n2143), .B1(n29353), .ZN(n2144) );
  I_NAND2 U1787 ( .A1(n2145), .B1(n29353), .ZN(n2146) );
  I_NAND2 U1788 ( .A1(n2147), .B1(n29353), .ZN(n2148) );
  I_NAND2 U1789 ( .A1(n2149), .B1(n29353), .ZN(n2150) );
  I_NAND2 U1790 ( .A1(n2151), .B1(n29353), .ZN(n2152) );
  I_NAND2 U1791 ( .A1(n2153), .B1(n29353), .ZN(n2154) );
  I_NAND2 U1792 ( .A1(n2155), .B1(n29353), .ZN(n2156) );
  I_NAND2 U1793 ( .A1(n2159), .B1(n29353), .ZN(n2160) );
  I_NAND2 U1794 ( .A1(n2162), .B1(n29353), .ZN(n2163) );
  I_NAND2 U1795 ( .A1(n2164), .B1(n29354), .ZN(n2165) );
  I_NAND2 U1796 ( .A1(n2166), .B1(n29364), .ZN(n2167) );
  I_NAND2 U1797 ( .A1(n2168), .B1(n29471), .ZN(n2169) );
  I_NAND2 U1798 ( .A1(n2170), .B1(n29466), .ZN(n2171) );
  I_NAND2 U1799 ( .A1(n2172), .B1(n29460), .ZN(n2173) );
  I_NAND2 U1800 ( .A1(n2174), .B1(n29460), .ZN(n2175) );
  I_NAND2 U1801 ( .A1(n2176), .B1(n29460), .ZN(n2177) );
  I_NAND2 U1802 ( .A1(n2178), .B1(n29461), .ZN(n2179) );
  I_NAND2 U1803 ( .A1(n2180), .B1(n29461), .ZN(n2181) );
  I_NAND2 U1804 ( .A1(n2182), .B1(n29461), .ZN(n2183) );
  I_NAND2 U1805 ( .A1(n2184), .B1(n29461), .ZN(n2185) );
  I_NAND2 U1806 ( .A1(n2186), .B1(n29461), .ZN(n2187) );
  I_NAND2 U1807 ( .A1(n2188), .B1(n29461), .ZN(n2189) );
  I_NAND2 U1808 ( .A1(n2190), .B1(n29461), .ZN(n2191) );
  I_NAND2 U1809 ( .A1(n2192), .B1(n29461), .ZN(n2193) );
  I_NAND2 U1810 ( .A1(n2194), .B1(n29461), .ZN(n2195) );
  I_NAND2 U1811 ( .A1(n2196), .B1(n29461), .ZN(n2197) );
  I_NAND2 U1812 ( .A1(n2198), .B1(n29461), .ZN(n2199) );
  I_NAND2 U1813 ( .A1(n2200), .B1(n29461), .ZN(n2201) );
  I_NAND2 U1814 ( .A1(n2202), .B1(n29462), .ZN(n2203) );
  I_NAND2 U1815 ( .A1(n2204), .B1(n29462), .ZN(n2205) );
  I_NAND2 U1816 ( .A1(n2206), .B1(n29462), .ZN(n2207) );
  I_NAND2 U1817 ( .A1(n2208), .B1(n29462), .ZN(n2209) );
  I_NAND2 U1818 ( .A1(n2210), .B1(n29462), .ZN(n2211) );
  I_NAND2 U1819 ( .A1(n2212), .B1(n29462), .ZN(n2213) );
  I_NAND2 U1820 ( .A1(n2214), .B1(n29462), .ZN(n2215) );
  I_NAND2 U1821 ( .A1(n2216), .B1(n29462), .ZN(n2217) );
  I_NAND2 U1822 ( .A1(n2218), .B1(n29462), .ZN(n2219) );
  I_NAND2 U1823 ( .A1(n2220), .B1(n29462), .ZN(n2221) );
  I_NAND2 U1824 ( .A1(n2222), .B1(n29462), .ZN(n2223) );
  I_NAND2 U1825 ( .A1(n2224), .B1(n29462), .ZN(n2225) );
  I_NAND2 U1826 ( .A1(n2226), .B1(n29463), .ZN(n2227) );
  I_NAND2 U1827 ( .A1(n2228), .B1(n29463), .ZN(n2229) );
  I_NAND2 U1828 ( .A1(n2230), .B1(n29463), .ZN(n2231) );
  I_NAND2 U1829 ( .A1(n2232), .B1(n29463), .ZN(n2233) );
  I_NAND2 U1830 ( .A1(n2234), .B1(n29463), .ZN(n2235) );
  I_NAND2 U1831 ( .A1(n2236), .B1(n29463), .ZN(n2237) );
  I_NAND2 U1832 ( .A1(n2238), .B1(n29463), .ZN(n2239) );
  I_NAND2 U1833 ( .A1(n2240), .B1(n29463), .ZN(n2241) );
  I_NAND2 U1834 ( .A1(n2242), .B1(n29463), .ZN(n2243) );
  I_NAND2 U1835 ( .A1(n2244), .B1(n29463), .ZN(n2245) );
  I_NAND2 U1836 ( .A1(n2246), .B1(n29463), .ZN(n2247) );
  I_NAND2 U1837 ( .A1(n2248), .B1(n29463), .ZN(n2249) );
  I_NAND2 U1838 ( .A1(n2250), .B1(n29464), .ZN(n2251) );
  I_NAND2 U1839 ( .A1(n2252), .B1(n29464), .ZN(n2253) );
  I_NAND2 U1840 ( .A1(n2254), .B1(n29464), .ZN(n2255) );
  I_NAND2 U1841 ( .A1(n2256), .B1(n29464), .ZN(n2257) );
  I_NAND2 U1842 ( .A1(n2258), .B1(n29464), .ZN(n2259) );
  I_NAND2 U1843 ( .A1(n2260), .B1(n29464), .ZN(n2261) );
  I_NAND2 U1844 ( .A1(n2262), .B1(n29464), .ZN(n2263) );
  I_NAND2 U1845 ( .A1(n2264), .B1(n29464), .ZN(n2265) );
  I_NAND2 U1846 ( .A1(n2266), .B1(n29464), .ZN(n2267) );
  I_NAND2 U1847 ( .A1(n2268), .B1(n29464), .ZN(n2269) );
  I_NAND2 U1848 ( .A1(n2270), .B1(n29464), .ZN(n2271) );
  I_NAND2 U1849 ( .A1(n2272), .B1(n29464), .ZN(n2273) );
  I_NAND2 U1850 ( .A1(n2274), .B1(n29465), .ZN(n2275) );
  I_NAND2 U1851 ( .A1(n2276), .B1(n29465), .ZN(n2277) );
  I_NAND2 U1852 ( .A1(n2278), .B1(n29465), .ZN(n2279) );
  I_NAND2 U1853 ( .A1(n2280), .B1(n29465), .ZN(n2281) );
  I_NAND2 U1854 ( .A1(n2282), .B1(n29465), .ZN(n2283) );
  I_NAND2 U1855 ( .A1(n2284), .B1(n29465), .ZN(n2285) );
  I_NAND2 U1856 ( .A1(n2286), .B1(n29465), .ZN(n2287) );
  I_NAND2 U1857 ( .A1(n2289), .B1(n29465), .ZN(n2290) );
  I_NAND2 U1858 ( .A1(n2292), .B1(n29465), .ZN(n2293) );
  I_NAND2 U1859 ( .A1(n2294), .B1(n29465), .ZN(n2295) );
  I_NAND2 U1860 ( .A1(n2296), .B1(n29465), .ZN(n2297) );
  I_NAND2 U1861 ( .A1(n2298), .B1(n29465), .ZN(n2299) );
  I_NAND2 U1862 ( .A1(n2300), .B1(n29466), .ZN(n2301) );
  I_NAND2 U1863 ( .A1(n2302), .B1(n29466), .ZN(n2303) );
  I_NAND2 U1864 ( .A1(n2304), .B1(n29466), .ZN(n2305) );
  I_NAND2 U1865 ( .A1(n2306), .B1(n29466), .ZN(n2307) );
  I_NAND2 U1866 ( .A1(n2308), .B1(n29466), .ZN(n2309) );
  I_NAND2 U1867 ( .A1(n2310), .B1(n29466), .ZN(n2311) );
  I_NAND2 U1868 ( .A1(n2312), .B1(n29466), .ZN(n2313) );
  I_NAND2 U1869 ( .A1(n2314), .B1(n29466), .ZN(n2315) );
  I_NAND2 U1870 ( .A1(n2316), .B1(n29466), .ZN(n2317) );
  I_NAND2 U1871 ( .A1(n2318), .B1(n29466), .ZN(n2319) );
  I_NAND2 U1872 ( .A1(n2320), .B1(n29466), .ZN(n2321) );
  I_NAND2 U1873 ( .A1(n2322), .B1(n29467), .ZN(n2323) );
  I_NAND2 U1874 ( .A1(n2324), .B1(n29467), .ZN(n2325) );
  I_NAND2 U1875 ( .A1(n2326), .B1(n29467), .ZN(n2327) );
  I_NAND2 U1876 ( .A1(n2328), .B1(n29467), .ZN(n2329) );
  I_NAND2 U1877 ( .A1(n2330), .B1(n29467), .ZN(n2331) );
  I_NAND2 U1878 ( .A1(n2332), .B1(n29467), .ZN(n2333) );
  I_NAND2 U1879 ( .A1(n2334), .B1(n29467), .ZN(n2335) );
  I_NAND2 U1880 ( .A1(n2336), .B1(n29467), .ZN(n2337) );
  I_NAND2 U1881 ( .A1(n2338), .B1(n29467), .ZN(n2339) );
  I_NAND2 U1882 ( .A1(n2340), .B1(n29467), .ZN(n2341) );
  I_NAND2 U1883 ( .A1(n2342), .B1(n29467), .ZN(n2343) );
  I_NAND2 U1884 ( .A1(n2344), .B1(n29467), .ZN(n2345) );
  I_NAND2 U1885 ( .A1(n2346), .B1(n29468), .ZN(n2347) );
  I_NAND2 U1886 ( .A1(n2348), .B1(n29468), .ZN(n2349) );
  I_NAND2 U1887 ( .A1(n2350), .B1(n29468), .ZN(n2351) );
  I_NAND2 U1888 ( .A1(n2352), .B1(n29468), .ZN(n2353) );
  I_NAND2 U1889 ( .A1(n2354), .B1(n29468), .ZN(n2355) );
  I_NAND2 U1890 ( .A1(n2356), .B1(n29468), .ZN(n2357) );
  I_NAND2 U1891 ( .A1(n2358), .B1(n29468), .ZN(n2359) );
  I_NAND2 U1892 ( .A1(n2360), .B1(n29468), .ZN(n2361) );
  I_NAND2 U1893 ( .A1(n2362), .B1(n29468), .ZN(n2363) );
  I_NAND2 U1894 ( .A1(n2364), .B1(n29468), .ZN(n2365) );
  I_NAND2 U1895 ( .A1(n2366), .B1(n29468), .ZN(n2367) );
  I_NAND2 U1896 ( .A1(n2368), .B1(n29468), .ZN(n2369) );
  I_NAND2 U1897 ( .A1(n2370), .B1(n29469), .ZN(n2371) );
  I_NAND2 U1898 ( .A1(n2372), .B1(n29469), .ZN(n2373) );
  I_NAND2 U1899 ( .A1(n2374), .B1(n29469), .ZN(n2375) );
  I_NAND2 U1900 ( .A1(n2376), .B1(n29469), .ZN(n2377) );
  I_NAND2 U1901 ( .A1(n2378), .B1(n29469), .ZN(n2379) );
  I_NAND2 U1902 ( .A1(n2380), .B1(n29469), .ZN(n2381) );
  I_NAND2 U1903 ( .A1(n2382), .B1(n29469), .ZN(n2383) );
  I_NAND2 U1904 ( .A1(n2384), .B1(n29469), .ZN(n2385) );
  I_NAND2 U1905 ( .A1(n2386), .B1(n29469), .ZN(n2387) );
  I_NAND2 U1906 ( .A1(n2388), .B1(n29469), .ZN(n2389) );
  I_NAND2 U1907 ( .A1(n2390), .B1(n29469), .ZN(n2391) );
  I_NAND2 U1908 ( .A1(n2392), .B1(n29469), .ZN(n2393) );
  I_NAND2 U1909 ( .A1(n2394), .B1(n29470), .ZN(n2395) );
  I_NAND2 U1910 ( .A1(n2396), .B1(n29470), .ZN(n2397) );
  I_NAND2 U1911 ( .A1(n2398), .B1(n29470), .ZN(n2399) );
  I_NAND2 U1912 ( .A1(n2400), .B1(n29470), .ZN(n2401) );
  I_NAND2 U1913 ( .A1(n2402), .B1(n29470), .ZN(n2403) );
  I_NAND2 U1914 ( .A1(n2404), .B1(n29470), .ZN(n2405) );
  I_NAND2 U1915 ( .A1(n2406), .B1(n29470), .ZN(n2407) );
  I_NAND2 U1916 ( .A1(n2408), .B1(n29470), .ZN(n2409) );
  I_NAND2 U1917 ( .A1(n2410), .B1(n29470), .ZN(n2411) );
  I_NAND2 U1918 ( .A1(n2412), .B1(n29470), .ZN(n2413) );
  I_NAND2 U1919 ( .A1(n2414), .B1(n29470), .ZN(n2415) );
  I_NAND2 U1920 ( .A1(n2416), .B1(n29470), .ZN(n2417) );
  I_NAND2 U1921 ( .A1(n2418), .B1(n29471), .ZN(n2419) );
  I_NAND2 U1922 ( .A1(n2421), .B1(n29471), .ZN(n2422) );
  I_NAND2 U1923 ( .A1(n2423), .B1(n29471), .ZN(n2424) );
  I_NAND2 U1924 ( .A1(n2425), .B1(n29471), .ZN(n2426) );
  I_NAND2 U1925 ( .A1(n2427), .B1(n29455), .ZN(n2428) );
  I_NAND2 U1926 ( .A1(n2429), .B1(n29450), .ZN(n2430) );
  I_NAND2 U1927 ( .A1(n2431), .B1(n29450), .ZN(n2432) );
  I_NAND2 U1928 ( .A1(n2433), .B1(n29450), .ZN(n2434) );
  I_NAND2 U1929 ( .A1(n2435), .B1(n29450), .ZN(n2436) );
  I_NAND2 U1930 ( .A1(n2437), .B1(n29450), .ZN(n2438) );
  I_NAND2 U1931 ( .A1(n2439), .B1(n29450), .ZN(n2440) );
  I_NAND2 U1932 ( .A1(n2441), .B1(n29450), .ZN(n2442) );
  I_NAND2 U1933 ( .A1(n2443), .B1(n29450), .ZN(n2444) );
  I_NAND2 U1934 ( .A1(n2445), .B1(n29450), .ZN(n2446) );
  I_NAND2 U1935 ( .A1(n2447), .B1(n29450), .ZN(n2448) );
  I_NAND2 U1936 ( .A1(n2449), .B1(n29451), .ZN(n2450) );
  I_NAND2 U1937 ( .A1(n2451), .B1(n29451), .ZN(n2452) );
  I_NAND2 U1938 ( .A1(n2453), .B1(n29451), .ZN(n2454) );
  I_NAND2 U1939 ( .A1(n2455), .B1(n29451), .ZN(n2456) );
  I_NAND2 U1940 ( .A1(n2457), .B1(n29451), .ZN(n2458) );
  I_NAND2 U1941 ( .A1(n2459), .B1(n29451), .ZN(n2460) );
  I_NAND2 U1942 ( .A1(n2461), .B1(n29451), .ZN(n2462) );
  I_NAND2 U1943 ( .A1(n2463), .B1(n29451), .ZN(n2464) );
  I_NAND2 U1944 ( .A1(n2465), .B1(n29451), .ZN(n2466) );
  I_NAND2 U1945 ( .A1(n2467), .B1(n29451), .ZN(n2468) );
  I_NAND2 U1946 ( .A1(n2469), .B1(n29451), .ZN(n2470) );
  I_NAND2 U1947 ( .A1(n2471), .B1(n29451), .ZN(n2472) );
  I_NAND2 U1948 ( .A1(n2473), .B1(n29452), .ZN(n2474) );
  I_NAND2 U1949 ( .A1(n2475), .B1(n29452), .ZN(n2476) );
  I_NAND2 U1950 ( .A1(n2477), .B1(n29452), .ZN(n2478) );
  I_NAND2 U1951 ( .A1(n2479), .B1(n29452), .ZN(n2480) );
  I_NAND2 U1952 ( .A1(n2481), .B1(n29452), .ZN(n2482) );
  I_NAND2 U1953 ( .A1(n2483), .B1(n29452), .ZN(n2484) );
  I_NAND2 U1954 ( .A1(n2485), .B1(n29452), .ZN(n2486) );
  I_NAND2 U1955 ( .A1(n2487), .B1(n29452), .ZN(n2488) );
  I_NAND2 U1956 ( .A1(n2489), .B1(n29452), .ZN(n2490) );
  I_NAND2 U1957 ( .A1(n2491), .B1(n29452), .ZN(n2492) );
  I_NAND2 U1958 ( .A1(n2493), .B1(n29452), .ZN(n2494) );
  I_NAND2 U1959 ( .A1(n2495), .B1(n29452), .ZN(n2496) );
  I_NAND2 U1960 ( .A1(n2497), .B1(n29453), .ZN(n2498) );
  I_NAND2 U1961 ( .A1(n2499), .B1(n29453), .ZN(n2500) );
  I_NAND2 U1962 ( .A1(n2501), .B1(n29453), .ZN(n2502) );
  I_NAND2 U1963 ( .A1(n2503), .B1(n29453), .ZN(n2504) );
  I_NAND2 U1964 ( .A1(n2505), .B1(n29453), .ZN(n2506) );
  I_NAND2 U1965 ( .A1(n2507), .B1(n29453), .ZN(n2508) );
  I_NAND2 U1966 ( .A1(n2509), .B1(n29453), .ZN(n2510) );
  I_NAND2 U1967 ( .A1(n2511), .B1(n29453), .ZN(n2512) );
  I_NAND2 U1968 ( .A1(n2513), .B1(n29453), .ZN(n2514) );
  I_NAND2 U1969 ( .A1(n2515), .B1(n29453), .ZN(n2516) );
  I_NAND2 U1970 ( .A1(n2517), .B1(n29453), .ZN(n2518) );
  I_NAND2 U1971 ( .A1(n2519), .B1(n29453), .ZN(n2520) );
  I_NAND2 U1972 ( .A1(n2521), .B1(n29454), .ZN(n2522) );
  I_NAND2 U1973 ( .A1(n2523), .B1(n29454), .ZN(n2524) );
  I_NAND2 U1974 ( .A1(n2525), .B1(n29454), .ZN(n2526) );
  I_NAND2 U1975 ( .A1(n2527), .B1(n29454), .ZN(n2528) );
  I_NAND2 U1976 ( .A1(n2529), .B1(n29454), .ZN(n2530) );
  I_NAND2 U1977 ( .A1(n2531), .B1(n29454), .ZN(n2532) );
  I_NAND2 U1978 ( .A1(n2533), .B1(n29454), .ZN(n2534) );
  I_NAND2 U1979 ( .A1(n2535), .B1(n29454), .ZN(n2536) );
  I_NAND2 U1980 ( .A1(n2537), .B1(n29454), .ZN(n2538) );
  I_NAND2 U1981 ( .A1(n2539), .B1(n29454), .ZN(n2540) );
  I_NAND2 U1982 ( .A1(n2541), .B1(n29454), .ZN(n2542) );
  I_NAND2 U1983 ( .A1(n2543), .B1(n29454), .ZN(n2544) );
  I_NAND2 U1984 ( .A1(n2545), .B1(n29455), .ZN(n2546) );
  I_NAND2 U1985 ( .A1(n2547), .B1(n29455), .ZN(n2548) );
  I_NAND2 U1986 ( .A1(n2550), .B1(n29455), .ZN(n2551) );
  I_NAND2 U1987 ( .A1(n2552), .B1(n29455), .ZN(n2553) );
  I_NAND2 U1988 ( .A1(n2554), .B1(n29455), .ZN(n2555) );
  I_NAND2 U1989 ( .A1(n2556), .B1(n29455), .ZN(n2557) );
  I_NAND2 U1990 ( .A1(n2558), .B1(n29455), .ZN(n2559) );
  I_NAND2 U1991 ( .A1(n2560), .B1(n29455), .ZN(n2561) );
  I_NAND2 U1992 ( .A1(n2562), .B1(n29455), .ZN(n2563) );
  I_NAND2 U1993 ( .A1(n2564), .B1(n29455), .ZN(n2565) );
  I_NAND2 U1994 ( .A1(n2566), .B1(n29455), .ZN(n2567) );
  I_NAND2 U1995 ( .A1(n2568), .B1(n29456), .ZN(n2569) );
  I_NAND2 U1996 ( .A1(n2570), .B1(n29456), .ZN(n2571) );
  I_NAND2 U1997 ( .A1(n2572), .B1(n29456), .ZN(n2573) );
  I_NAND2 U1998 ( .A1(n2574), .B1(n29456), .ZN(n2575) );
  I_NAND2 U1999 ( .A1(n2576), .B1(n29456), .ZN(n2577) );
  I_NAND2 U2000 ( .A1(n2578), .B1(n29456), .ZN(n2579) );
  I_NAND2 U2001 ( .A1(n2580), .B1(n29456), .ZN(n2581) );
  I_NAND2 U2002 ( .A1(n2582), .B1(n29456), .ZN(n2583) );
  I_NAND2 U2003 ( .A1(n2584), .B1(n29456), .ZN(n2585) );
  I_NAND2 U2004 ( .A1(n2586), .B1(n29456), .ZN(n2587) );
  I_NAND2 U2005 ( .A1(n2588), .B1(n29456), .ZN(n2589) );
  I_NAND2 U2006 ( .A1(n2590), .B1(n29456), .ZN(n2591) );
  I_NAND2 U2007 ( .A1(n2592), .B1(n29457), .ZN(n2593) );
  I_NAND2 U2008 ( .A1(n2594), .B1(n29457), .ZN(n2595) );
  I_NAND2 U2009 ( .A1(n2596), .B1(n29457), .ZN(n2597) );
  I_NAND2 U2010 ( .A1(n2598), .B1(n29457), .ZN(n2599) );
  I_NAND2 U2011 ( .A1(n2600), .B1(n29457), .ZN(n2601) );
  I_NAND2 U2012 ( .A1(n2602), .B1(n29457), .ZN(n2603) );
  I_NAND2 U2013 ( .A1(n2604), .B1(n29457), .ZN(n2605) );
  I_NAND2 U2014 ( .A1(n2606), .B1(n29457), .ZN(n2607) );
  I_NAND2 U2015 ( .A1(n2608), .B1(n29457), .ZN(n2609) );
  I_NAND2 U2016 ( .A1(n2610), .B1(n29457), .ZN(n2611) );
  I_NAND2 U2017 ( .A1(n2612), .B1(n29457), .ZN(n2613) );
  I_NAND2 U2018 ( .A1(n2614), .B1(n29457), .ZN(n2615) );
  I_NAND2 U2019 ( .A1(n2616), .B1(n29458), .ZN(n2617) );
  I_NAND2 U2020 ( .A1(n2618), .B1(n29458), .ZN(n2619) );
  I_NAND2 U2021 ( .A1(n2620), .B1(n29458), .ZN(n2621) );
  I_NAND2 U2022 ( .A1(n2622), .B1(n29458), .ZN(n2623) );
  I_NAND2 U2023 ( .A1(n2624), .B1(n29458), .ZN(n2625) );
  I_NAND2 U2024 ( .A1(n2626), .B1(n29458), .ZN(n2627) );
  I_NAND2 U2025 ( .A1(n2628), .B1(n29458), .ZN(n2629) );
  I_NAND2 U2026 ( .A1(n2630), .B1(n29458), .ZN(n2631) );
  I_NAND2 U2027 ( .A1(n2632), .B1(n29458), .ZN(n2633) );
  I_NAND2 U2028 ( .A1(n2634), .B1(n29458), .ZN(n2635) );
  I_NAND2 U2029 ( .A1(n2636), .B1(n29458), .ZN(n2637) );
  I_NAND2 U2030 ( .A1(n2638), .B1(n29458), .ZN(n2639) );
  I_NAND2 U2031 ( .A1(n2640), .B1(n29459), .ZN(n2641) );
  I_NAND2 U2032 ( .A1(n2642), .B1(n29459), .ZN(n2643) );
  I_NAND2 U2033 ( .A1(n2644), .B1(n29459), .ZN(n2645) );
  I_NAND2 U2034 ( .A1(n2646), .B1(n29459), .ZN(n2647) );
  I_NAND2 U2035 ( .A1(n2648), .B1(n29459), .ZN(n2649) );
  I_NAND2 U2036 ( .A1(n2650), .B1(n29459), .ZN(n2651) );
  I_NAND2 U2037 ( .A1(n2652), .B1(n29459), .ZN(n2653) );
  I_NAND2 U2038 ( .A1(n2654), .B1(n29459), .ZN(n2655) );
  I_NAND2 U2039 ( .A1(n2656), .B1(n29459), .ZN(n2657) );
  I_NAND2 U2040 ( .A1(n2658), .B1(n29459), .ZN(n2659) );
  I_NAND2 U2041 ( .A1(n2660), .B1(n29459), .ZN(n2661) );
  I_NAND2 U2042 ( .A1(n2662), .B1(n29459), .ZN(n2663) );
  I_NAND2 U2043 ( .A1(n2664), .B1(n29460), .ZN(n2665) );
  I_NAND2 U2044 ( .A1(n2666), .B1(n29460), .ZN(n2667) );
  I_NAND2 U2045 ( .A1(n2668), .B1(n29460), .ZN(n2669) );
  I_NAND2 U2046 ( .A1(n2670), .B1(n29460), .ZN(n2671) );
  I_NAND2 U2047 ( .A1(n2672), .B1(n29460), .ZN(n2673) );
  I_NAND2 U2048 ( .A1(n2674), .B1(n29460), .ZN(n2675) );
  I_NAND2 U2049 ( .A1(n2676), .B1(n29460), .ZN(n2677) );
  I_NAND2 U2050 ( .A1(n2805), .B1(n29487), .ZN(n2806) );
  I_NAND2 U2051 ( .A1(n2934), .B1(n29492), .ZN(n2935) );
  I_NAND2 U2052 ( .A1(n3063), .B1(n29476), .ZN(n3064) );
  I_NAND2 U2053 ( .A1(n3192), .B1(n29481), .ZN(n3193) );
  I_NAND2 U2054 ( .A1(n3322), .B1(n29423), .ZN(n3323) );
  I_NAND2 U2055 ( .A1(n3451), .B1(n29428), .ZN(n3452) );
  I_NAND2 U2056 ( .A1(n3580), .B1(n29412), .ZN(n3581) );
  I_NAND2 U2057 ( .A1(n3709), .B1(n29418), .ZN(n3710) );
  I_NAND2 U2058 ( .A1(n3838), .B1(n29444), .ZN(n3839) );
  I_NAND2 U2059 ( .A1(n3967), .B1(n29450), .ZN(n3968) );
  I_NAND2 U2060 ( .A1(n4096), .B1(n29434), .ZN(n4097) );
  NAND2 U2061 ( .A1(n23), .A2(n27434), .ZN(n13) );
  I_NAND2 U2062 ( .A1(n1123), .B1(n29396), .ZN(n1124) );
  I_NAND2 U2063 ( .A1(n2157), .B1(n29353), .ZN(n2158) );
  BUF U2064 ( .I(n29497), .Z(n29483) );
  BUF U2065 ( .I(n29497), .Z(n29484) );
  BUF U2066 ( .I(n29496), .Z(n29485) );
  BUF U2067 ( .I(n29496), .Z(n29486) );
  BUF U2068 ( .I(n29496), .Z(n29487) );
  BUF U2069 ( .I(n29495), .Z(n29488) );
  BUF U2070 ( .I(n29495), .Z(n29489) );
  BUF U2071 ( .I(n29495), .Z(n29490) );
  BUF U2072 ( .I(n29500), .Z(n29473) );
  BUF U2073 ( .I(n29500), .Z(n29474) );
  BUF U2074 ( .I(n29500), .Z(n29475) );
  BUF U2075 ( .I(n29499), .Z(n29476) );
  BUF U2076 ( .I(n29499), .Z(n29477) );
  BUF U2077 ( .I(n29499), .Z(n29478) );
  BUF U2078 ( .I(n29498), .Z(n29479) );
  BUF U2079 ( .I(n29498), .Z(n29480) );
  BUF U2080 ( .I(n29498), .Z(n29481) );
  BUF U2081 ( .I(n29497), .Z(n29482) );
  BUF U2082 ( .I(n29551), .Z(n29322) );
  BUF U2083 ( .I(n29552), .Z(n29551) );
  BUF U2084 ( .I(n29558), .Z(n29532) );
  BUF U2085 ( .I(n29558), .Z(n29531) );
  BUF U2086 ( .I(n29559), .Z(n29530) );
  BUF U2087 ( .I(n29557), .Z(n29536) );
  BUF U2088 ( .I(n29557), .Z(n29535) );
  BUF U2089 ( .I(n29557), .Z(n29534) );
  BUF U2090 ( .I(n29558), .Z(n29533) );
  BUF U2091 ( .I(n29560), .Z(n29525) );
  BUF U2092 ( .I(n29561), .Z(n29524) );
  BUF U2093 ( .I(n29561), .Z(n29523) );
  BUF U2094 ( .I(n29559), .Z(n29529) );
  BUF U2095 ( .I(n29559), .Z(n29528) );
  BUF U2096 ( .I(n29560), .Z(n29527) );
  BUF U2097 ( .I(n29560), .Z(n29526) );
  BUF U2098 ( .I(n29553), .Z(n29546) );
  BUF U2099 ( .I(n29554), .Z(n29545) );
  BUF U2100 ( .I(n29552), .Z(n29550) );
  BUF U2101 ( .I(n29552), .Z(n29549) );
  BUF U2102 ( .I(n29553), .Z(n29548) );
  BUF U2103 ( .I(n29553), .Z(n29547) );
  BUF U2104 ( .I(n29556), .Z(n29539) );
  BUF U2105 ( .I(n29556), .Z(n29538) );
  BUF U2106 ( .I(n29554), .Z(n29544) );
  BUF U2107 ( .I(n29554), .Z(n29543) );
  BUF U2108 ( .I(n29555), .Z(n29542) );
  BUF U2109 ( .I(n29555), .Z(n29541) );
  BUF U2110 ( .I(n29555), .Z(n29540) );
  BUF U2111 ( .I(n29556), .Z(n29537) );
  BUF U2112 ( .I(n29567), .Z(n29504) );
  BUF U2113 ( .I(n29568), .Z(n29503) );
  BUF U2114 ( .I(n29568), .Z(n29502) );
  BUF U2115 ( .I(n29566), .Z(n29507) );
  BUF U2116 ( .I(n29567), .Z(n29506) );
  BUF U2117 ( .I(n29567), .Z(n29505) );
  BUF U2118 ( .I(n29568), .Z(n29501) );
  BUF U2119 ( .I(n29563), .Z(n29518) );
  BUF U2120 ( .I(n29563), .Z(n29517) );
  BUF U2121 ( .I(n29563), .Z(n29516) );
  BUF U2122 ( .I(n29561), .Z(n29522) );
  BUF U2123 ( .I(n29562), .Z(n29521) );
  BUF U2124 ( .I(n29562), .Z(n29520) );
  BUF U2125 ( .I(n29562), .Z(n29519) );
  BUF U2126 ( .I(n29565), .Z(n29511) );
  BUF U2127 ( .I(n29565), .Z(n29510) );
  BUF U2128 ( .I(n29566), .Z(n29509) );
  BUF U2129 ( .I(n29566), .Z(n29508) );
  BUF U2130 ( .I(n29564), .Z(n29515) );
  BUF U2131 ( .I(n29564), .Z(n29514) );
  BUF U2132 ( .I(n29564), .Z(n29513) );
  BUF U2133 ( .I(n29565), .Z(n29512) );
  BUF U2134 ( .I(n27020), .Z(n27032) );
  BUF U2135 ( .I(n27021), .Z(n27029) );
  BUF U2136 ( .I(n27021), .Z(n27031) );
  BUF U2137 ( .I(n27021), .Z(n27030) );
  BUF U2138 ( .I(n27022), .Z(n27028) );
  BUF U2139 ( .I(n27022), .Z(n27027) );
  BUF U2140 ( .I(n27022), .Z(n27026) );
  BUF U2141 ( .I(n27007), .Z(n27071) );
  BUF U2142 ( .I(n27007), .Z(n27072) );
  BUF U2143 ( .I(n27008), .Z(n27070) );
  BUF U2144 ( .I(n27008), .Z(n27069) );
  BUF U2145 ( .I(n27009), .Z(n27066) );
  BUF U2146 ( .I(n27008), .Z(n27068) );
  BUF U2147 ( .I(n27009), .Z(n27067) );
  BUF U2148 ( .I(n27009), .Z(n27065) );
  BUF U2149 ( .I(n27010), .Z(n27064) );
  BUF U2150 ( .I(n27011), .Z(n27061) );
  BUF U2151 ( .I(n27010), .Z(n27063) );
  BUF U2152 ( .I(n27010), .Z(n27062) );
  BUF U2153 ( .I(n27011), .Z(n27060) );
  BUF U2154 ( .I(n27011), .Z(n27059) );
  BUF U2155 ( .I(n27012), .Z(n27056) );
  BUF U2156 ( .I(n27012), .Z(n27058) );
  BUF U2157 ( .I(n27012), .Z(n27057) );
  BUF U2158 ( .I(n27013), .Z(n27055) );
  BUF U2159 ( .I(n27013), .Z(n27054) );
  BUF U2160 ( .I(n27017), .Z(n27042) );
  BUF U2161 ( .I(n27017), .Z(n27041) );
  BUF U2162 ( .I(n27018), .Z(n27040) );
  BUF U2163 ( .I(n27018), .Z(n27039) );
  BUF U2164 ( .I(n27018), .Z(n27038) );
  BUF U2165 ( .I(n27019), .Z(n27037) );
  BUF U2166 ( .I(n27020), .Z(n27034) );
  BUF U2167 ( .I(n27020), .Z(n27033) );
  BUF U2168 ( .I(n27019), .Z(n27036) );
  BUF U2169 ( .I(n27019), .Z(n27035) );
  BUF U2170 ( .I(n27014), .Z(n27051) );
  BUF U2171 ( .I(n27013), .Z(n27053) );
  BUF U2172 ( .I(n27014), .Z(n27052) );
  BUF U2173 ( .I(n27014), .Z(n27050) );
  BUF U2174 ( .I(n27015), .Z(n27049) );
  BUF U2175 ( .I(n27015), .Z(n27048) );
  BUF U2176 ( .I(n27015), .Z(n27047) );
  BUF U2177 ( .I(n27017), .Z(n27043) );
  BUF U2178 ( .I(n27016), .Z(n27046) );
  BUF U2179 ( .I(n27016), .Z(n27045) );
  BUF U2180 ( .I(n27016), .Z(n27044) );
  BUF U2181 ( .I(n26999), .Z(n27097) );
  BUF U2182 ( .I(n26999), .Z(n27096) );
  BUF U2183 ( .I(n26999), .Z(n27095) );
  BUF U2184 ( .I(n27000), .Z(n27094) );
  BUF U2185 ( .I(n27000), .Z(n27093) );
  BUF U2186 ( .I(n27004), .Z(n27082) );
  BUF U2187 ( .I(n27004), .Z(n27081) );
  BUF U2188 ( .I(n27004), .Z(n27080) );
  BUF U2189 ( .I(n27005), .Z(n27079) );
  BUF U2190 ( .I(n27005), .Z(n27078) );
  BUF U2191 ( .I(n27005), .Z(n27077) );
  BUF U2192 ( .I(n27006), .Z(n27076) );
  BUF U2193 ( .I(n27007), .Z(n27073) );
  BUF U2194 ( .I(n27006), .Z(n27075) );
  BUF U2195 ( .I(n27006), .Z(n27074) );
  BUF U2196 ( .I(n27000), .Z(n27092) );
  BUF U2197 ( .I(n27001), .Z(n27091) );
  BUF U2198 ( .I(n27002), .Z(n27088) );
  BUF U2199 ( .I(n27001), .Z(n27090) );
  BUF U2200 ( .I(n27001), .Z(n27089) );
  BUF U2201 ( .I(n27002), .Z(n27087) );
  BUF U2202 ( .I(n27002), .Z(n27086) );
  BUF U2203 ( .I(n27003), .Z(n27083) );
  BUF U2204 ( .I(n27003), .Z(n27085) );
  BUF U2205 ( .I(n27003), .Z(n27084) );
  BUF U2206 ( .I(n26918), .Z(n27338) );
  BUF U2207 ( .I(n26917), .Z(n26918) );
  BUF U2208 ( .I(n26536), .Z(n26586) );
  BUF U2209 ( .I(n26537), .Z(n26581) );
  BUF U2210 ( .I(n26524), .Z(n26621) );
  BUF U2211 ( .I(n26892), .Z(n26994) );
  BUF U2212 ( .I(n26417), .Z(n26519) );
  BUF U2213 ( .I(n26892), .Z(n26995) );
  BUF U2214 ( .I(n26891), .Z(n26996) );
  BUF U2215 ( .I(n26891), .Z(n26997) );
  BUF U2216 ( .I(n26416), .Z(n26522) );
  BUF U2217 ( .I(n26896), .Z(n26981) );
  BUF U2218 ( .I(n26421), .Z(n26506) );
  BUF U2219 ( .I(n26896), .Z(n26982) );
  BUF U2220 ( .I(n26896), .Z(n26983) );
  BUF U2221 ( .I(n26901), .Z(n26968) );
  BUF U2222 ( .I(n26426), .Z(n26493) );
  BUF U2223 ( .I(n26900), .Z(n26969) );
  BUF U2224 ( .I(n26900), .Z(n26970) );
  BUF U2225 ( .I(n26905), .Z(n26955) );
  BUF U2226 ( .I(n26430), .Z(n26480) );
  BUF U2227 ( .I(n26905), .Z(n26956) );
  BUF U2228 ( .I(n26904), .Z(n26957) );
  BUF U2229 ( .I(n26909), .Z(n26942) );
  BUF U2230 ( .I(n26434), .Z(n26467) );
  BUF U2231 ( .I(n26909), .Z(n26943) );
  BUF U2232 ( .I(n26909), .Z(n26944) );
  BUF U2233 ( .I(n26914), .Z(n26929) );
  BUF U2234 ( .I(n26439), .Z(n26454) );
  BUF U2235 ( .I(n26913), .Z(n26930) );
  BUF U2236 ( .I(n26913), .Z(n26931) );
  BUF U2237 ( .I(n26891), .Z(n26998) );
  BUF U2238 ( .I(n26895), .Z(n26984) );
  BUF U2239 ( .I(n26420), .Z(n26509) );
  BUF U2240 ( .I(n26895), .Z(n26985) );
  BUF U2241 ( .I(n26895), .Z(n26986) );
  BUF U2242 ( .I(n26420), .Z(n26511) );
  BUF U2243 ( .I(n26893), .Z(n26991) );
  BUF U2244 ( .I(n26418), .Z(n26516) );
  BUF U2245 ( .I(n26893), .Z(n26992) );
  BUF U2246 ( .I(n26892), .Z(n26993) );
  BUF U2247 ( .I(n26894), .Z(n26987) );
  BUF U2248 ( .I(n26894), .Z(n26988) );
  BUF U2249 ( .I(n26894), .Z(n26989) );
  BUF U2250 ( .I(n26893), .Z(n26990) );
  BUF U2251 ( .I(n26900), .Z(n26971) );
  BUF U2252 ( .I(n26425), .Z(n26496) );
  BUF U2253 ( .I(n26899), .Z(n26972) );
  BUF U2254 ( .I(n26899), .Z(n26973) );
  BUF U2255 ( .I(n26424), .Z(n26498) );
  BUF U2256 ( .I(n26897), .Z(n26978) );
  BUF U2257 ( .I(n26422), .Z(n26503) );
  BUF U2258 ( .I(n26897), .Z(n26979) );
  BUF U2259 ( .I(n26897), .Z(n26980) );
  BUF U2260 ( .I(n26899), .Z(n26974) );
  BUF U2261 ( .I(n26898), .Z(n26975) );
  BUF U2262 ( .I(n26898), .Z(n26976) );
  BUF U2263 ( .I(n26898), .Z(n26977) );
  BUF U2264 ( .I(n26904), .Z(n26958) );
  BUF U2265 ( .I(n26429), .Z(n26483) );
  BUF U2266 ( .I(n26904), .Z(n26959) );
  BUF U2267 ( .I(n26903), .Z(n26960) );
  BUF U2268 ( .I(n26428), .Z(n26485) );
  BUF U2269 ( .I(n26902), .Z(n26965) );
  BUF U2270 ( .I(n26427), .Z(n26490) );
  BUF U2271 ( .I(n26901), .Z(n26966) );
  BUF U2272 ( .I(n26901), .Z(n26967) );
  BUF U2273 ( .I(n26903), .Z(n26961) );
  BUF U2274 ( .I(n26903), .Z(n26962) );
  BUF U2275 ( .I(n26902), .Z(n26963) );
  BUF U2276 ( .I(n26902), .Z(n26964) );
  BUF U2277 ( .I(n26908), .Z(n26945) );
  BUF U2278 ( .I(n26433), .Z(n26470) );
  BUF U2279 ( .I(n26908), .Z(n26946) );
  BUF U2280 ( .I(n26908), .Z(n26947) );
  BUF U2281 ( .I(n26433), .Z(n26472) );
  BUF U2282 ( .I(n26906), .Z(n26952) );
  BUF U2283 ( .I(n26431), .Z(n26477) );
  BUF U2284 ( .I(n26906), .Z(n26953) );
  BUF U2285 ( .I(n26905), .Z(n26954) );
  BUF U2286 ( .I(n26907), .Z(n26948) );
  BUF U2287 ( .I(n26907), .Z(n26949) );
  BUF U2288 ( .I(n26907), .Z(n26950) );
  BUF U2289 ( .I(n26906), .Z(n26951) );
  BUF U2290 ( .I(n26913), .Z(n26932) );
  BUF U2291 ( .I(n26438), .Z(n26457) );
  BUF U2292 ( .I(n26912), .Z(n26933) );
  BUF U2293 ( .I(n26437), .Z(n26458) );
  BUF U2294 ( .I(n26912), .Z(n26934) );
  BUF U2295 ( .I(n26910), .Z(n26939) );
  BUF U2296 ( .I(n26910), .Z(n26940) );
  BUF U2297 ( .I(n26910), .Z(n26941) );
  BUF U2298 ( .I(n26912), .Z(n26935) );
  BUF U2299 ( .I(n26911), .Z(n26936) );
  BUF U2300 ( .I(n26911), .Z(n26938) );
  BUF U2301 ( .I(n26436), .Z(n26463) );
  BUF U2302 ( .I(n26911), .Z(n26937) );
  BUF U2303 ( .I(n26917), .Z(n26919) );
  BUF U2304 ( .I(n26442), .Z(n26444) );
  BUF U2305 ( .I(n26917), .Z(n26920) );
  BUF U2306 ( .I(n26442), .Z(n26445) );
  BUF U2307 ( .I(n26915), .Z(n26926) );
  BUF U2308 ( .I(n26914), .Z(n26927) );
  BUF U2309 ( .I(n26914), .Z(n26928) );
  BUF U2310 ( .I(n26916), .Z(n26921) );
  BUF U2311 ( .I(n26916), .Z(n26922) );
  BUF U2312 ( .I(n26916), .Z(n26923) );
  BUF U2313 ( .I(n26915), .Z(n26925) );
  BUF U2314 ( .I(n26440), .Z(n26450) );
  BUF U2315 ( .I(n26915), .Z(n26924) );
  BUF U2316 ( .I(n26443), .Z(n26863) );
  BUF U2317 ( .I(n26442), .Z(n26443) );
  BUF U2318 ( .I(n26545), .Z(n26557) );
  BUF U2319 ( .I(n26546), .Z(n26554) );
  BUF U2320 ( .I(n26546), .Z(n26556) );
  BUF U2321 ( .I(n26546), .Z(n26555) );
  BUF U2322 ( .I(n26547), .Z(n26553) );
  BUF U2323 ( .I(n26547), .Z(n26552) );
  BUF U2324 ( .I(n26547), .Z(n26551) );
  BUF U2325 ( .I(n26532), .Z(n26596) );
  BUF U2326 ( .I(n26532), .Z(n26597) );
  BUF U2327 ( .I(n26533), .Z(n26595) );
  BUF U2328 ( .I(n26533), .Z(n26594) );
  BUF U2329 ( .I(n26534), .Z(n26591) );
  BUF U2330 ( .I(n26533), .Z(n26593) );
  BUF U2331 ( .I(n26534), .Z(n26592) );
  BUF U2332 ( .I(n26534), .Z(n26590) );
  BUF U2333 ( .I(n26535), .Z(n26589) );
  BUF U2334 ( .I(n26535), .Z(n26588) );
  BUF U2335 ( .I(n26535), .Z(n26587) );
  BUF U2336 ( .I(n26536), .Z(n26585) );
  BUF U2337 ( .I(n26536), .Z(n26584) );
  BUF U2338 ( .I(n26537), .Z(n26583) );
  BUF U2339 ( .I(n26537), .Z(n26582) );
  BUF U2340 ( .I(n26538), .Z(n26580) );
  BUF U2341 ( .I(n26538), .Z(n26579) );
  BUF U2342 ( .I(n26542), .Z(n26567) );
  BUF U2343 ( .I(n26542), .Z(n26566) );
  BUF U2344 ( .I(n26543), .Z(n26565) );
  BUF U2345 ( .I(n26543), .Z(n26564) );
  BUF U2346 ( .I(n26543), .Z(n26563) );
  BUF U2347 ( .I(n26544), .Z(n26562) );
  BUF U2348 ( .I(n26545), .Z(n26559) );
  BUF U2349 ( .I(n26545), .Z(n26558) );
  BUF U2350 ( .I(n26544), .Z(n26561) );
  BUF U2351 ( .I(n26544), .Z(n26560) );
  BUF U2352 ( .I(n26539), .Z(n26576) );
  BUF U2353 ( .I(n26538), .Z(n26578) );
  BUF U2354 ( .I(n26539), .Z(n26577) );
  BUF U2355 ( .I(n26539), .Z(n26575) );
  BUF U2356 ( .I(n26540), .Z(n26574) );
  BUF U2357 ( .I(n26540), .Z(n26573) );
  BUF U2358 ( .I(n26540), .Z(n26572) );
  BUF U2359 ( .I(n26542), .Z(n26568) );
  BUF U2360 ( .I(n26541), .Z(n26571) );
  BUF U2361 ( .I(n26541), .Z(n26570) );
  BUF U2362 ( .I(n26541), .Z(n26569) );
  BUF U2363 ( .I(n26524), .Z(n26622) );
  BUF U2364 ( .I(n26524), .Z(n26620) );
  BUF U2365 ( .I(n26525), .Z(n26619) );
  BUF U2366 ( .I(n26525), .Z(n26618) );
  BUF U2367 ( .I(n26529), .Z(n26607) );
  BUF U2368 ( .I(n26529), .Z(n26606) );
  BUF U2369 ( .I(n26529), .Z(n26605) );
  BUF U2370 ( .I(n26530), .Z(n26604) );
  BUF U2371 ( .I(n26530), .Z(n26603) );
  BUF U2372 ( .I(n26530), .Z(n26602) );
  BUF U2373 ( .I(n26531), .Z(n26601) );
  BUF U2374 ( .I(n26532), .Z(n26598) );
  BUF U2375 ( .I(n26531), .Z(n26600) );
  BUF U2376 ( .I(n26531), .Z(n26599) );
  BUF U2377 ( .I(n26525), .Z(n26617) );
  BUF U2378 ( .I(n26526), .Z(n26616) );
  BUF U2379 ( .I(n26527), .Z(n26613) );
  BUF U2380 ( .I(n26526), .Z(n26615) );
  BUF U2381 ( .I(n26526), .Z(n26614) );
  BUF U2382 ( .I(n26527), .Z(n26612) );
  BUF U2383 ( .I(n26527), .Z(n26611) );
  BUF U2384 ( .I(n26528), .Z(n26608) );
  BUF U2385 ( .I(n26528), .Z(n26610) );
  BUF U2386 ( .I(n26528), .Z(n26609) );
  BUF U2387 ( .I(n26417), .Z(n26520) );
  BUF U2388 ( .I(n26416), .Z(n26521) );
  BUF U2389 ( .I(n26421), .Z(n26507) );
  BUF U2390 ( .I(n26421), .Z(n26508) );
  BUF U2391 ( .I(n26425), .Z(n26494) );
  BUF U2392 ( .I(n26425), .Z(n26495) );
  BUF U2393 ( .I(n26430), .Z(n26481) );
  BUF U2394 ( .I(n26429), .Z(n26482) );
  BUF U2395 ( .I(n26434), .Z(n26468) );
  BUF U2396 ( .I(n26434), .Z(n26469) );
  BUF U2397 ( .I(n26438), .Z(n26455) );
  BUF U2398 ( .I(n26438), .Z(n26456) );
  BUF U2399 ( .I(n26416), .Z(n26523) );
  BUF U2400 ( .I(n26420), .Z(n26510) );
  BUF U2401 ( .I(n26418), .Z(n26517) );
  BUF U2402 ( .I(n26417), .Z(n26518) );
  BUF U2403 ( .I(n26419), .Z(n26512) );
  BUF U2404 ( .I(n26419), .Z(n26513) );
  BUF U2405 ( .I(n26419), .Z(n26514) );
  BUF U2406 ( .I(n26418), .Z(n26515) );
  BUF U2407 ( .I(n26424), .Z(n26497) );
  BUF U2408 ( .I(n26422), .Z(n26504) );
  BUF U2409 ( .I(n26422), .Z(n26505) );
  BUF U2410 ( .I(n26424), .Z(n26499) );
  BUF U2411 ( .I(n26423), .Z(n26500) );
  BUF U2412 ( .I(n26423), .Z(n26501) );
  BUF U2413 ( .I(n26423), .Z(n26502) );
  BUF U2414 ( .I(n26429), .Z(n26484) );
  BUF U2415 ( .I(n26426), .Z(n26491) );
  BUF U2416 ( .I(n26426), .Z(n26492) );
  BUF U2417 ( .I(n26428), .Z(n26486) );
  BUF U2418 ( .I(n26428), .Z(n26487) );
  BUF U2419 ( .I(n26427), .Z(n26488) );
  BUF U2420 ( .I(n26427), .Z(n26489) );
  BUF U2421 ( .I(n26433), .Z(n26471) );
  BUF U2422 ( .I(n26431), .Z(n26478) );
  BUF U2423 ( .I(n26430), .Z(n26479) );
  BUF U2424 ( .I(n26432), .Z(n26473) );
  BUF U2425 ( .I(n26432), .Z(n26474) );
  BUF U2426 ( .I(n26432), .Z(n26475) );
  BUF U2427 ( .I(n26431), .Z(n26476) );
  BUF U2428 ( .I(n26437), .Z(n26459) );
  BUF U2429 ( .I(n26435), .Z(n26464) );
  BUF U2430 ( .I(n26435), .Z(n26465) );
  BUF U2431 ( .I(n26435), .Z(n26466) );
  BUF U2432 ( .I(n26437), .Z(n26460) );
  BUF U2433 ( .I(n26436), .Z(n26461) );
  BUF U2434 ( .I(n26436), .Z(n26462) );
  BUF U2435 ( .I(n26440), .Z(n26451) );
  BUF U2436 ( .I(n26439), .Z(n26452) );
  BUF U2437 ( .I(n26439), .Z(n26453) );
  BUF U2438 ( .I(n26441), .Z(n26446) );
  BUF U2439 ( .I(n26441), .Z(n26447) );
  BUF U2440 ( .I(n26441), .Z(n26448) );
  BUF U2441 ( .I(n26440), .Z(n26449) );
  INV U2442 ( .I(n198), .ZN(n27434) );
  INV U2443 ( .I(n198), .ZN(n27435) );
  INV U2444 ( .I(n198), .ZN(n27436) );
  I_NAND2 U2445 ( .A1(n2679), .B1(n29460), .ZN(n2680) );
  I_NAND2 U2446 ( .A1(n2681), .B1(n29460), .ZN(n2682) );
  I_NAND2 U2447 ( .A1(n2683), .B1(n29487), .ZN(n2684) );
  I_NAND2 U2448 ( .A1(n2685), .B1(n29482), .ZN(n2686) );
  I_NAND2 U2449 ( .A1(n2687), .B1(n29482), .ZN(n2688) );
  I_NAND2 U2450 ( .A1(n2689), .B1(n29482), .ZN(n2690) );
  I_NAND2 U2451 ( .A1(n2691), .B1(n29482), .ZN(n2692) );
  I_NAND2 U2452 ( .A1(n2693), .B1(n29482), .ZN(n2694) );
  I_NAND2 U2453 ( .A1(n2695), .B1(n29482), .ZN(n2696) );
  I_NAND2 U2454 ( .A1(n2697), .B1(n29482), .ZN(n2698) );
  I_NAND2 U2455 ( .A1(n2699), .B1(n29482), .ZN(n2700) );
  I_NAND2 U2456 ( .A1(n2701), .B1(n29482), .ZN(n2702) );
  I_NAND2 U2457 ( .A1(n2703), .B1(n29482), .ZN(n2704) );
  I_NAND2 U2458 ( .A1(n2705), .B1(n29482), .ZN(n2706) );
  I_NAND2 U2459 ( .A1(n2707), .B1(n29483), .ZN(n2708) );
  I_NAND2 U2460 ( .A1(n2709), .B1(n29483), .ZN(n2710) );
  I_NAND2 U2461 ( .A1(n2711), .B1(n29483), .ZN(n2712) );
  I_NAND2 U2462 ( .A1(n2713), .B1(n29483), .ZN(n2714) );
  I_NAND2 U2463 ( .A1(n2715), .B1(n29483), .ZN(n2716) );
  I_NAND2 U2464 ( .A1(n2717), .B1(n29483), .ZN(n2718) );
  I_NAND2 U2465 ( .A1(n2719), .B1(n29483), .ZN(n2720) );
  I_NAND2 U2466 ( .A1(n2721), .B1(n29483), .ZN(n2722) );
  I_NAND2 U2467 ( .A1(n2723), .B1(n29483), .ZN(n2724) );
  I_NAND2 U2468 ( .A1(n2725), .B1(n29483), .ZN(n2726) );
  I_NAND2 U2469 ( .A1(n2727), .B1(n29483), .ZN(n2728) );
  I_NAND2 U2470 ( .A1(n2729), .B1(n29483), .ZN(n2730) );
  I_NAND2 U2471 ( .A1(n2731), .B1(n29484), .ZN(n2732) );
  I_NAND2 U2472 ( .A1(n2733), .B1(n29484), .ZN(n2734) );
  I_NAND2 U2473 ( .A1(n2735), .B1(n29484), .ZN(n2736) );
  I_NAND2 U2474 ( .A1(n2737), .B1(n29484), .ZN(n2738) );
  I_NAND2 U2475 ( .A1(n2739), .B1(n29484), .ZN(n2740) );
  I_NAND2 U2476 ( .A1(n2741), .B1(n29484), .ZN(n2742) );
  I_NAND2 U2477 ( .A1(n2743), .B1(n29484), .ZN(n2744) );
  I_NAND2 U2478 ( .A1(n2745), .B1(n29484), .ZN(n2746) );
  I_NAND2 U2479 ( .A1(n2747), .B1(n29484), .ZN(n2748) );
  I_NAND2 U2480 ( .A1(n2749), .B1(n29484), .ZN(n2750) );
  I_NAND2 U2481 ( .A1(n2751), .B1(n29484), .ZN(n2752) );
  I_NAND2 U2482 ( .A1(n2753), .B1(n29484), .ZN(n2754) );
  I_NAND2 U2483 ( .A1(n2755), .B1(n29485), .ZN(n2756) );
  I_NAND2 U2484 ( .A1(n2757), .B1(n29485), .ZN(n2758) );
  I_NAND2 U2485 ( .A1(n2759), .B1(n29485), .ZN(n2760) );
  I_NAND2 U2486 ( .A1(n2761), .B1(n29485), .ZN(n2762) );
  I_NAND2 U2487 ( .A1(n2763), .B1(n29485), .ZN(n2764) );
  I_NAND2 U2488 ( .A1(n2765), .B1(n29485), .ZN(n2766) );
  I_NAND2 U2489 ( .A1(n2767), .B1(n29485), .ZN(n2768) );
  I_NAND2 U2490 ( .A1(n2769), .B1(n29485), .ZN(n2770) );
  I_NAND2 U2491 ( .A1(n2771), .B1(n29485), .ZN(n2772) );
  I_NAND2 U2492 ( .A1(n2773), .B1(n29485), .ZN(n2774) );
  I_NAND2 U2493 ( .A1(n2775), .B1(n29485), .ZN(n2776) );
  I_NAND2 U2494 ( .A1(n2777), .B1(n29485), .ZN(n2778) );
  I_NAND2 U2495 ( .A1(n2779), .B1(n29486), .ZN(n2780) );
  I_NAND2 U2496 ( .A1(n2781), .B1(n29486), .ZN(n2782) );
  I_NAND2 U2497 ( .A1(n2783), .B1(n29486), .ZN(n2784) );
  I_NAND2 U2498 ( .A1(n2785), .B1(n29486), .ZN(n2786) );
  I_NAND2 U2499 ( .A1(n2787), .B1(n29486), .ZN(n2788) );
  I_NAND2 U2500 ( .A1(n2789), .B1(n29486), .ZN(n2790) );
  I_NAND2 U2501 ( .A1(n2791), .B1(n29486), .ZN(n2792) );
  I_NAND2 U2502 ( .A1(n2793), .B1(n29486), .ZN(n2794) );
  I_NAND2 U2503 ( .A1(n2795), .B1(n29486), .ZN(n2796) );
  I_NAND2 U2504 ( .A1(n2797), .B1(n29486), .ZN(n2798) );
  I_NAND2 U2505 ( .A1(n2799), .B1(n29486), .ZN(n2800) );
  I_NAND2 U2506 ( .A1(n2801), .B1(n29486), .ZN(n2802) );
  I_NAND2 U2507 ( .A1(n2803), .B1(n29487), .ZN(n2804) );
  I_NAND2 U2508 ( .A1(n2808), .B1(n29487), .ZN(n2809) );
  I_NAND2 U2509 ( .A1(n2810), .B1(n29487), .ZN(n2811) );
  I_NAND2 U2510 ( .A1(n2812), .B1(n29487), .ZN(n2813) );
  I_NAND2 U2511 ( .A1(n2814), .B1(n29487), .ZN(n2815) );
  I_NAND2 U2512 ( .A1(n2816), .B1(n29487), .ZN(n2817) );
  I_NAND2 U2513 ( .A1(n2818), .B1(n29487), .ZN(n2819) );
  I_NAND2 U2514 ( .A1(n2820), .B1(n29487), .ZN(n2821) );
  I_NAND2 U2515 ( .A1(n2822), .B1(n29487), .ZN(n2823) );
  I_NAND2 U2516 ( .A1(n2824), .B1(n29487), .ZN(n2825) );
  I_NAND2 U2517 ( .A1(n2826), .B1(n29488), .ZN(n2827) );
  I_NAND2 U2518 ( .A1(n2828), .B1(n29488), .ZN(n2829) );
  I_NAND2 U2519 ( .A1(n2830), .B1(n29488), .ZN(n2831) );
  I_NAND2 U2520 ( .A1(n2832), .B1(n29488), .ZN(n2833) );
  I_NAND2 U2521 ( .A1(n2834), .B1(n29488), .ZN(n2835) );
  I_NAND2 U2522 ( .A1(n2836), .B1(n29488), .ZN(n2837) );
  I_NAND2 U2523 ( .A1(n2838), .B1(n29488), .ZN(n2839) );
  I_NAND2 U2524 ( .A1(n2840), .B1(n29488), .ZN(n2841) );
  I_NAND2 U2525 ( .A1(n2842), .B1(n29488), .ZN(n2843) );
  I_NAND2 U2526 ( .A1(n2844), .B1(n29488), .ZN(n2845) );
  I_NAND2 U2527 ( .A1(n2846), .B1(n29488), .ZN(n2847) );
  I_NAND2 U2528 ( .A1(n2848), .B1(n29488), .ZN(n2849) );
  I_NAND2 U2529 ( .A1(n2850), .B1(n29489), .ZN(n2851) );
  I_NAND2 U2530 ( .A1(n2852), .B1(n29489), .ZN(n2853) );
  I_NAND2 U2531 ( .A1(n2854), .B1(n29489), .ZN(n2855) );
  I_NAND2 U2532 ( .A1(n2856), .B1(n29489), .ZN(n2857) );
  I_NAND2 U2533 ( .A1(n2858), .B1(n29489), .ZN(n2859) );
  I_NAND2 U2534 ( .A1(n2860), .B1(n29489), .ZN(n2861) );
  I_NAND2 U2535 ( .A1(n2862), .B1(n29489), .ZN(n2863) );
  I_NAND2 U2536 ( .A1(n2864), .B1(n29489), .ZN(n2865) );
  I_NAND2 U2537 ( .A1(n2866), .B1(n29489), .ZN(n2867) );
  I_NAND2 U2538 ( .A1(n2868), .B1(n29489), .ZN(n2869) );
  I_NAND2 U2539 ( .A1(n2870), .B1(n29489), .ZN(n2871) );
  I_NAND2 U2540 ( .A1(n2872), .B1(n29489), .ZN(n2873) );
  I_NAND2 U2541 ( .A1(n2874), .B1(n29490), .ZN(n2875) );
  I_NAND2 U2542 ( .A1(n2876), .B1(n29490), .ZN(n2877) );
  I_NAND2 U2543 ( .A1(n2878), .B1(n29490), .ZN(n2879) );
  I_NAND2 U2544 ( .A1(n2880), .B1(n29490), .ZN(n2881) );
  I_NAND2 U2545 ( .A1(n2882), .B1(n29490), .ZN(n2883) );
  I_NAND2 U2546 ( .A1(n2884), .B1(n29490), .ZN(n2885) );
  I_NAND2 U2547 ( .A1(n2886), .B1(n29490), .ZN(n2887) );
  I_NAND2 U2548 ( .A1(n2888), .B1(n29490), .ZN(n2889) );
  I_NAND2 U2549 ( .A1(n2890), .B1(n29490), .ZN(n2891) );
  I_NAND2 U2550 ( .A1(n2892), .B1(n29490), .ZN(n2893) );
  I_NAND2 U2551 ( .A1(n2894), .B1(n29490), .ZN(n2895) );
  I_NAND2 U2552 ( .A1(n2896), .B1(n29490), .ZN(n2897) );
  I_NAND2 U2553 ( .A1(n2898), .B1(n29491), .ZN(n2899) );
  I_NAND2 U2554 ( .A1(n2900), .B1(n29491), .ZN(n2901) );
  I_NAND2 U2555 ( .A1(n2902), .B1(n29491), .ZN(n2903) );
  I_NAND2 U2556 ( .A1(n2904), .B1(n29491), .ZN(n2905) );
  I_NAND2 U2557 ( .A1(n2906), .B1(n29491), .ZN(n2907) );
  I_NAND2 U2558 ( .A1(n2908), .B1(n29491), .ZN(n2909) );
  I_NAND2 U2559 ( .A1(n2910), .B1(n29491), .ZN(n2911) );
  I_NAND2 U2560 ( .A1(n2912), .B1(n29491), .ZN(n2913) );
  I_NAND2 U2561 ( .A1(n2914), .B1(n29491), .ZN(n2915) );
  I_NAND2 U2562 ( .A1(n2916), .B1(n29491), .ZN(n2917) );
  I_NAND2 U2563 ( .A1(n2918), .B1(n29491), .ZN(n2919) );
  I_NAND2 U2564 ( .A1(n2920), .B1(n29491), .ZN(n2921) );
  I_NAND2 U2565 ( .A1(n2922), .B1(n29492), .ZN(n2923) );
  I_NAND2 U2566 ( .A1(n2924), .B1(n29492), .ZN(n2925) );
  I_NAND2 U2567 ( .A1(n2926), .B1(n29492), .ZN(n2927) );
  I_NAND2 U2568 ( .A1(n2928), .B1(n29492), .ZN(n2929) );
  I_NAND2 U2569 ( .A1(n2930), .B1(n29492), .ZN(n2931) );
  I_NAND2 U2570 ( .A1(n2932), .B1(n29492), .ZN(n2933) );
  I_NAND2 U2571 ( .A1(n2937), .B1(n29492), .ZN(n2938) );
  I_NAND2 U2572 ( .A1(n2939), .B1(n29476), .ZN(n2940) );
  I_NAND2 U2573 ( .A1(n2941), .B1(n29471), .ZN(n2942) );
  I_NAND2 U2574 ( .A1(n2943), .B1(n29471), .ZN(n2944) );
  I_NAND2 U2575 ( .A1(n2945), .B1(n29471), .ZN(n2946) );
  I_NAND2 U2576 ( .A1(n2947), .B1(n29471), .ZN(n2948) );
  I_NAND2 U2577 ( .A1(n2949), .B1(n29471), .ZN(n2950) );
  I_NAND2 U2578 ( .A1(n2951), .B1(n29471), .ZN(n2952) );
  I_NAND2 U2579 ( .A1(n2953), .B1(n29471), .ZN(n2954) );
  I_NAND2 U2580 ( .A1(n2955), .B1(n29472), .ZN(n2956) );
  I_NAND2 U2581 ( .A1(n2957), .B1(n29472), .ZN(n2958) );
  I_NAND2 U2582 ( .A1(n2959), .B1(n29472), .ZN(n2960) );
  I_NAND2 U2583 ( .A1(n2961), .B1(n29472), .ZN(n2962) );
  I_NAND2 U2584 ( .A1(n2963), .B1(n29472), .ZN(n2964) );
  I_NAND2 U2585 ( .A1(n2965), .B1(n29472), .ZN(n2966) );
  I_NAND2 U2586 ( .A1(n2967), .B1(n29472), .ZN(n2968) );
  I_NAND2 U2587 ( .A1(n2969), .B1(n29472), .ZN(n2970) );
  I_NAND2 U2588 ( .A1(n2971), .B1(n29472), .ZN(n2972) );
  I_NAND2 U2589 ( .A1(n2973), .B1(n29472), .ZN(n2974) );
  I_NAND2 U2590 ( .A1(n2975), .B1(n29472), .ZN(n2976) );
  I_NAND2 U2591 ( .A1(n2977), .B1(n29472), .ZN(n2978) );
  I_NAND2 U2592 ( .A1(n2979), .B1(n29473), .ZN(n2980) );
  I_NAND2 U2593 ( .A1(n2981), .B1(n29473), .ZN(n2982) );
  I_NAND2 U2594 ( .A1(n2983), .B1(n29473), .ZN(n2984) );
  I_NAND2 U2595 ( .A1(n2985), .B1(n29473), .ZN(n2986) );
  I_NAND2 U2596 ( .A1(n2987), .B1(n29473), .ZN(n2988) );
  I_NAND2 U2597 ( .A1(n2989), .B1(n29473), .ZN(n2990) );
  I_NAND2 U2598 ( .A1(n2991), .B1(n29473), .ZN(n2992) );
  I_NAND2 U2599 ( .A1(n2993), .B1(n29473), .ZN(n2994) );
  I_NAND2 U2600 ( .A1(n2995), .B1(n29473), .ZN(n2996) );
  I_NAND2 U2601 ( .A1(n2997), .B1(n29473), .ZN(n2998) );
  I_NAND2 U2602 ( .A1(n2999), .B1(n29473), .ZN(n3000) );
  I_NAND2 U2603 ( .A1(n3001), .B1(n29473), .ZN(n3002) );
  I_NAND2 U2604 ( .A1(n3003), .B1(n29474), .ZN(n3004) );
  I_NAND2 U2605 ( .A1(n3005), .B1(n29474), .ZN(n3006) );
  I_NAND2 U2606 ( .A1(n3007), .B1(n29474), .ZN(n3008) );
  I_NAND2 U2607 ( .A1(n3009), .B1(n29474), .ZN(n3010) );
  I_NAND2 U2608 ( .A1(n3011), .B1(n29474), .ZN(n3012) );
  I_NAND2 U2609 ( .A1(n3013), .B1(n29474), .ZN(n3014) );
  I_NAND2 U2610 ( .A1(n3015), .B1(n29474), .ZN(n3016) );
  I_NAND2 U2611 ( .A1(n3017), .B1(n29474), .ZN(n3018) );
  I_NAND2 U2612 ( .A1(n3019), .B1(n29474), .ZN(n3020) );
  I_NAND2 U2613 ( .A1(n3021), .B1(n29474), .ZN(n3022) );
  I_NAND2 U2614 ( .A1(n3023), .B1(n29474), .ZN(n3024) );
  I_NAND2 U2615 ( .A1(n3025), .B1(n29474), .ZN(n3026) );
  I_NAND2 U2616 ( .A1(n3027), .B1(n29475), .ZN(n3028) );
  I_NAND2 U2617 ( .A1(n3029), .B1(n29475), .ZN(n3030) );
  I_NAND2 U2618 ( .A1(n3031), .B1(n29475), .ZN(n3032) );
  I_NAND2 U2619 ( .A1(n3033), .B1(n29475), .ZN(n3034) );
  I_NAND2 U2620 ( .A1(n3035), .B1(n29475), .ZN(n3036) );
  I_NAND2 U2621 ( .A1(n3037), .B1(n29475), .ZN(n3038) );
  I_NAND2 U2622 ( .A1(n3039), .B1(n29475), .ZN(n3040) );
  I_NAND2 U2623 ( .A1(n3041), .B1(n29475), .ZN(n3042) );
  I_NAND2 U2624 ( .A1(n3043), .B1(n29475), .ZN(n3044) );
  I_NAND2 U2625 ( .A1(n3045), .B1(n29475), .ZN(n3046) );
  I_NAND2 U2626 ( .A1(n3047), .B1(n29475), .ZN(n3048) );
  I_NAND2 U2627 ( .A1(n3049), .B1(n29475), .ZN(n3050) );
  I_NAND2 U2628 ( .A1(n3051), .B1(n29476), .ZN(n3052) );
  I_NAND2 U2629 ( .A1(n3053), .B1(n29476), .ZN(n3054) );
  I_NAND2 U2630 ( .A1(n3055), .B1(n29476), .ZN(n3056) );
  I_NAND2 U2631 ( .A1(n3057), .B1(n29476), .ZN(n3058) );
  I_NAND2 U2632 ( .A1(n3059), .B1(n29476), .ZN(n3060) );
  I_NAND2 U2633 ( .A1(n3061), .B1(n29476), .ZN(n3062) );
  I_NAND2 U2634 ( .A1(n3066), .B1(n29476), .ZN(n3067) );
  I_NAND2 U2635 ( .A1(n3068), .B1(n29476), .ZN(n3069) );
  I_NAND2 U2636 ( .A1(n3070), .B1(n29476), .ZN(n3071) );
  I_NAND2 U2637 ( .A1(n3072), .B1(n29476), .ZN(n3073) );
  I_NAND2 U2638 ( .A1(n3074), .B1(n29477), .ZN(n3075) );
  I_NAND2 U2639 ( .A1(n3076), .B1(n29477), .ZN(n3077) );
  I_NAND2 U2640 ( .A1(n3078), .B1(n29477), .ZN(n3079) );
  I_NAND2 U2641 ( .A1(n3080), .B1(n29477), .ZN(n3081) );
  I_NAND2 U2642 ( .A1(n3082), .B1(n29477), .ZN(n3083) );
  I_NAND2 U2643 ( .A1(n3084), .B1(n29477), .ZN(n3085) );
  I_NAND2 U2644 ( .A1(n3086), .B1(n29477), .ZN(n3087) );
  I_NAND2 U2645 ( .A1(n3088), .B1(n29477), .ZN(n3089) );
  I_NAND2 U2646 ( .A1(n3090), .B1(n29477), .ZN(n3091) );
  I_NAND2 U2647 ( .A1(n3092), .B1(n29477), .ZN(n3093) );
  I_NAND2 U2648 ( .A1(n3094), .B1(n29477), .ZN(n3095) );
  I_NAND2 U2649 ( .A1(n3096), .B1(n29477), .ZN(n3097) );
  I_NAND2 U2650 ( .A1(n3098), .B1(n29478), .ZN(n3099) );
  I_NAND2 U2651 ( .A1(n3100), .B1(n29478), .ZN(n3101) );
  I_NAND2 U2652 ( .A1(n3102), .B1(n29478), .ZN(n3103) );
  I_NAND2 U2653 ( .A1(n3104), .B1(n29478), .ZN(n3105) );
  I_NAND2 U2654 ( .A1(n3106), .B1(n29478), .ZN(n3107) );
  I_NAND2 U2655 ( .A1(n3108), .B1(n29478), .ZN(n3109) );
  I_NAND2 U2656 ( .A1(n3110), .B1(n29478), .ZN(n3111) );
  I_NAND2 U2657 ( .A1(n3112), .B1(n29478), .ZN(n3113) );
  I_NAND2 U2658 ( .A1(n3114), .B1(n29478), .ZN(n3115) );
  I_NAND2 U2659 ( .A1(n3116), .B1(n29478), .ZN(n3117) );
  I_NAND2 U2660 ( .A1(n3118), .B1(n29478), .ZN(n3119) );
  I_NAND2 U2661 ( .A1(n3120), .B1(n29478), .ZN(n3121) );
  I_NAND2 U2662 ( .A1(n3122), .B1(n29479), .ZN(n3123) );
  I_NAND2 U2663 ( .A1(n3124), .B1(n29479), .ZN(n3125) );
  I_NAND2 U2664 ( .A1(n3126), .B1(n29479), .ZN(n3127) );
  I_NAND2 U2665 ( .A1(n3128), .B1(n29479), .ZN(n3129) );
  I_NAND2 U2666 ( .A1(n3130), .B1(n29479), .ZN(n3131) );
  I_NAND2 U2667 ( .A1(n3132), .B1(n29479), .ZN(n3133) );
  I_NAND2 U2668 ( .A1(n3134), .B1(n29479), .ZN(n3135) );
  I_NAND2 U2669 ( .A1(n3136), .B1(n29479), .ZN(n3137) );
  I_NAND2 U2670 ( .A1(n3138), .B1(n29479), .ZN(n3139) );
  I_NAND2 U2671 ( .A1(n3140), .B1(n29479), .ZN(n3141) );
  I_NAND2 U2672 ( .A1(n3142), .B1(n29479), .ZN(n3143) );
  I_NAND2 U2673 ( .A1(n3144), .B1(n29479), .ZN(n3145) );
  I_NAND2 U2674 ( .A1(n3146), .B1(n29480), .ZN(n3147) );
  I_NAND2 U2675 ( .A1(n3148), .B1(n29480), .ZN(n3149) );
  I_NAND2 U2676 ( .A1(n3150), .B1(n29480), .ZN(n3151) );
  I_NAND2 U2677 ( .A1(n3152), .B1(n29480), .ZN(n3153) );
  I_NAND2 U2678 ( .A1(n3154), .B1(n29480), .ZN(n3155) );
  I_NAND2 U2679 ( .A1(n3156), .B1(n29480), .ZN(n3157) );
  I_NAND2 U2680 ( .A1(n3158), .B1(n29480), .ZN(n3159) );
  I_NAND2 U2681 ( .A1(n3160), .B1(n29480), .ZN(n3161) );
  I_NAND2 U2682 ( .A1(n3162), .B1(n29480), .ZN(n3163) );
  I_NAND2 U2683 ( .A1(n3164), .B1(n29480), .ZN(n3165) );
  I_NAND2 U2684 ( .A1(n3166), .B1(n29480), .ZN(n3167) );
  I_NAND2 U2685 ( .A1(n3168), .B1(n29480), .ZN(n3169) );
  I_NAND2 U2686 ( .A1(n3170), .B1(n29481), .ZN(n3171) );
  I_NAND2 U2687 ( .A1(n3172), .B1(n29481), .ZN(n3173) );
  I_NAND2 U2688 ( .A1(n3174), .B1(n29481), .ZN(n3175) );
  I_NAND2 U2689 ( .A1(n3176), .B1(n29481), .ZN(n3177) );
  I_NAND2 U2690 ( .A1(n3178), .B1(n29481), .ZN(n3179) );
  I_NAND2 U2691 ( .A1(n3180), .B1(n29481), .ZN(n3181) );
  I_NAND2 U2692 ( .A1(n3182), .B1(n29481), .ZN(n3183) );
  I_NAND2 U2693 ( .A1(n3184), .B1(n29481), .ZN(n3185) );
  I_NAND2 U2694 ( .A1(n3186), .B1(n29481), .ZN(n3187) );
  I_NAND2 U2695 ( .A1(n3188), .B1(n29481), .ZN(n3189) );
  I_NAND2 U2696 ( .A1(n3195), .B1(n29482), .ZN(n3196) );
  I_NAND2 U2697 ( .A1(n3197), .B1(n29428), .ZN(n3198) );
  I_NAND2 U2698 ( .A1(n3199), .B1(n29423), .ZN(n3200) );
  I_NAND2 U2699 ( .A1(n3201), .B1(n29418), .ZN(n3202) );
  I_NAND2 U2700 ( .A1(n3203), .B1(n29418), .ZN(n3204) );
  I_NAND2 U2701 ( .A1(n3205), .B1(n29418), .ZN(n3206) );
  I_NAND2 U2702 ( .A1(n3207), .B1(n29418), .ZN(n3208) );
  I_NAND2 U2703 ( .A1(n3209), .B1(n29418), .ZN(n3210) );
  I_NAND2 U2704 ( .A1(n3211), .B1(n29418), .ZN(n3212) );
  I_NAND2 U2705 ( .A1(n3213), .B1(n29418), .ZN(n3214) );
  I_NAND2 U2706 ( .A1(n3215), .B1(n29418), .ZN(n3216) );
  I_NAND2 U2707 ( .A1(n3217), .B1(n29418), .ZN(n3218) );
  I_NAND2 U2708 ( .A1(n3219), .B1(n29419), .ZN(n3220) );
  I_NAND2 U2709 ( .A1(n3221), .B1(n29419), .ZN(n3222) );
  I_NAND2 U2710 ( .A1(n3223), .B1(n29419), .ZN(n3224) );
  I_NAND2 U2711 ( .A1(n3225), .B1(n29419), .ZN(n3226) );
  I_NAND2 U2712 ( .A1(n3227), .B1(n29419), .ZN(n3228) );
  I_NAND2 U2713 ( .A1(n3229), .B1(n29419), .ZN(n3230) );
  I_NAND2 U2714 ( .A1(n3231), .B1(n29419), .ZN(n3232) );
  I_NAND2 U2715 ( .A1(n3233), .B1(n29419), .ZN(n3234) );
  I_NAND2 U2716 ( .A1(n3235), .B1(n29419), .ZN(n3236) );
  I_NAND2 U2717 ( .A1(n3237), .B1(n29419), .ZN(n3238) );
  I_NAND2 U2718 ( .A1(n3239), .B1(n29419), .ZN(n3240) );
  I_NAND2 U2719 ( .A1(n3241), .B1(n29419), .ZN(n3242) );
  I_NAND2 U2720 ( .A1(n3243), .B1(n29420), .ZN(n3244) );
  I_NAND2 U2721 ( .A1(n3245), .B1(n29420), .ZN(n3246) );
  I_NAND2 U2722 ( .A1(n3247), .B1(n29420), .ZN(n3248) );
  I_NAND2 U2723 ( .A1(n3249), .B1(n29420), .ZN(n3250) );
  I_NAND2 U2724 ( .A1(n3251), .B1(n29420), .ZN(n3252) );
  I_NAND2 U2725 ( .A1(n3253), .B1(n29420), .ZN(n3254) );
  I_NAND2 U2726 ( .A1(n3255), .B1(n29420), .ZN(n3256) );
  I_NAND2 U2727 ( .A1(n3257), .B1(n29420), .ZN(n3258) );
  I_NAND2 U2728 ( .A1(n3259), .B1(n29420), .ZN(n3260) );
  I_NAND2 U2729 ( .A1(n3261), .B1(n29420), .ZN(n3262) );
  I_NAND2 U2730 ( .A1(n3263), .B1(n29420), .ZN(n3264) );
  I_NAND2 U2731 ( .A1(n3265), .B1(n29420), .ZN(n3266) );
  I_NAND2 U2732 ( .A1(n3267), .B1(n29421), .ZN(n3268) );
  I_NAND2 U2733 ( .A1(n3269), .B1(n29421), .ZN(n3270) );
  I_NAND2 U2734 ( .A1(n3271), .B1(n29421), .ZN(n3272) );
  I_NAND2 U2735 ( .A1(n3273), .B1(n29421), .ZN(n3274) );
  I_NAND2 U2736 ( .A1(n3275), .B1(n29421), .ZN(n3276) );
  I_NAND2 U2737 ( .A1(n3277), .B1(n29421), .ZN(n3278) );
  I_NAND2 U2738 ( .A1(n3279), .B1(n29421), .ZN(n3280) );
  I_NAND2 U2739 ( .A1(n3281), .B1(n29421), .ZN(n3282) );
  I_NAND2 U2740 ( .A1(n3283), .B1(n29421), .ZN(n3284) );
  I_NAND2 U2741 ( .A1(n3285), .B1(n29421), .ZN(n3286) );
  I_NAND2 U2742 ( .A1(n3287), .B1(n29421), .ZN(n3288) );
  I_NAND2 U2743 ( .A1(n3289), .B1(n29421), .ZN(n3290) );
  I_NAND2 U2744 ( .A1(n3291), .B1(n29422), .ZN(n3292) );
  I_NAND2 U2745 ( .A1(n3293), .B1(n29422), .ZN(n3294) );
  I_NAND2 U2746 ( .A1(n3295), .B1(n29422), .ZN(n3296) );
  I_NAND2 U2747 ( .A1(n3297), .B1(n29422), .ZN(n3298) );
  I_NAND2 U2748 ( .A1(n3299), .B1(n29422), .ZN(n3300) );
  I_NAND2 U2749 ( .A1(n3301), .B1(n29422), .ZN(n3302) );
  I_NAND2 U2750 ( .A1(n3303), .B1(n29422), .ZN(n3304) );
  I_NAND2 U2751 ( .A1(n3305), .B1(n29422), .ZN(n3306) );
  I_NAND2 U2752 ( .A1(n3307), .B1(n29422), .ZN(n3308) );
  I_NAND2 U2753 ( .A1(n3309), .B1(n29422), .ZN(n3310) );
  I_NAND2 U2754 ( .A1(n3311), .B1(n29422), .ZN(n3312) );
  I_NAND2 U2755 ( .A1(n3313), .B1(n29422), .ZN(n3314) );
  I_NAND2 U2756 ( .A1(n3315), .B1(n29423), .ZN(n3316) );
  I_NAND2 U2757 ( .A1(n3317), .B1(n29423), .ZN(n3318) );
  I_NAND2 U2758 ( .A1(n3319), .B1(n29423), .ZN(n3320) );
  I_NAND2 U2759 ( .A1(n3325), .B1(n29423), .ZN(n3326) );
  I_NAND2 U2760 ( .A1(n3327), .B1(n29423), .ZN(n3328) );
  I_NAND2 U2761 ( .A1(n3329), .B1(n29423), .ZN(n3330) );
  I_NAND2 U2762 ( .A1(n3331), .B1(n29423), .ZN(n3332) );
  I_NAND2 U2763 ( .A1(n3333), .B1(n29423), .ZN(n3334) );
  I_NAND2 U2764 ( .A1(n3335), .B1(n29423), .ZN(n3336) );
  I_NAND2 U2765 ( .A1(n3337), .B1(n29423), .ZN(n3338) );
  I_NAND2 U2766 ( .A1(n3339), .B1(n29424), .ZN(n3340) );
  I_NAND2 U2767 ( .A1(n3341), .B1(n29424), .ZN(n3342) );
  I_NAND2 U2768 ( .A1(n3343), .B1(n29424), .ZN(n3344) );
  I_NAND2 U2769 ( .A1(n3345), .B1(n29424), .ZN(n3346) );
  I_NAND2 U2770 ( .A1(n3347), .B1(n29424), .ZN(n3348) );
  I_NAND2 U2771 ( .A1(n3349), .B1(n29424), .ZN(n3350) );
  I_NAND2 U2772 ( .A1(n3351), .B1(n29424), .ZN(n3352) );
  I_NAND2 U2773 ( .A1(n3353), .B1(n29424), .ZN(n3354) );
  I_NAND2 U2774 ( .A1(n3355), .B1(n29424), .ZN(n3356) );
  I_NAND2 U2775 ( .A1(n3357), .B1(n29424), .ZN(n3358) );
  I_NAND2 U2776 ( .A1(n3359), .B1(n29424), .ZN(n3360) );
  I_NAND2 U2777 ( .A1(n3361), .B1(n29424), .ZN(n3362) );
  I_NAND2 U2778 ( .A1(n3363), .B1(n29425), .ZN(n3364) );
  I_NAND2 U2779 ( .A1(n3365), .B1(n29425), .ZN(n3366) );
  I_NAND2 U2780 ( .A1(n3367), .B1(n29425), .ZN(n3368) );
  I_NAND2 U2781 ( .A1(n3369), .B1(n29425), .ZN(n3370) );
  I_NAND2 U2782 ( .A1(n3371), .B1(n29425), .ZN(n3372) );
  I_NAND2 U2783 ( .A1(n3373), .B1(n29425), .ZN(n3374) );
  I_NAND2 U2784 ( .A1(n3375), .B1(n29425), .ZN(n3376) );
  I_NAND2 U2785 ( .A1(n3377), .B1(n29425), .ZN(n3378) );
  I_NAND2 U2786 ( .A1(n3379), .B1(n29425), .ZN(n3380) );
  I_NAND2 U2787 ( .A1(n3381), .B1(n29425), .ZN(n3382) );
  I_NAND2 U2788 ( .A1(n3383), .B1(n29425), .ZN(n3384) );
  I_NAND2 U2789 ( .A1(n3385), .B1(n29425), .ZN(n3386) );
  I_NAND2 U2790 ( .A1(n3387), .B1(n29426), .ZN(n3388) );
  I_NAND2 U2791 ( .A1(n3389), .B1(n29426), .ZN(n3390) );
  I_NAND2 U2792 ( .A1(n3391), .B1(n29426), .ZN(n3392) );
  I_NAND2 U2793 ( .A1(n3393), .B1(n29426), .ZN(n3394) );
  I_NAND2 U2794 ( .A1(n3395), .B1(n29426), .ZN(n3396) );
  I_NAND2 U2795 ( .A1(n3397), .B1(n29426), .ZN(n3398) );
  I_NAND2 U2796 ( .A1(n3399), .B1(n29426), .ZN(n3400) );
  I_NAND2 U2797 ( .A1(n3401), .B1(n29426), .ZN(n3402) );
  I_NAND2 U2798 ( .A1(n3403), .B1(n29426), .ZN(n3404) );
  I_NAND2 U2799 ( .A1(n3405), .B1(n29426), .ZN(n3406) );
  I_NAND2 U2800 ( .A1(n3407), .B1(n29426), .ZN(n3408) );
  I_NAND2 U2801 ( .A1(n3409), .B1(n29426), .ZN(n3410) );
  I_NAND2 U2802 ( .A1(n3411), .B1(n29427), .ZN(n3412) );
  I_NAND2 U2803 ( .A1(n3413), .B1(n29427), .ZN(n3414) );
  I_NAND2 U2804 ( .A1(n3415), .B1(n29427), .ZN(n3416) );
  I_NAND2 U2805 ( .A1(n3417), .B1(n29427), .ZN(n3418) );
  I_NAND2 U2806 ( .A1(n3419), .B1(n29427), .ZN(n3420) );
  I_NAND2 U2807 ( .A1(n3421), .B1(n29427), .ZN(n3422) );
  I_NAND2 U2808 ( .A1(n3423), .B1(n29427), .ZN(n3424) );
  I_NAND2 U2809 ( .A1(n3425), .B1(n29427), .ZN(n3426) );
  I_NAND2 U2810 ( .A1(n3427), .B1(n29427), .ZN(n3428) );
  I_NAND2 U2811 ( .A1(n3429), .B1(n29427), .ZN(n3430) );
  I_NAND2 U2812 ( .A1(n3431), .B1(n29427), .ZN(n3432) );
  I_NAND2 U2813 ( .A1(n3433), .B1(n29427), .ZN(n3434) );
  I_NAND2 U2814 ( .A1(n3435), .B1(n29428), .ZN(n3436) );
  I_NAND2 U2815 ( .A1(n3437), .B1(n29428), .ZN(n3438) );
  I_NAND2 U2816 ( .A1(n3439), .B1(n29428), .ZN(n3440) );
  I_NAND2 U2817 ( .A1(n3441), .B1(n29428), .ZN(n3442) );
  I_NAND2 U2818 ( .A1(n3443), .B1(n29428), .ZN(n3444) );
  I_NAND2 U2819 ( .A1(n3445), .B1(n29428), .ZN(n3446) );
  I_NAND2 U2820 ( .A1(n3447), .B1(n29428), .ZN(n3448) );
  I_NAND2 U2821 ( .A1(n3449), .B1(n29428), .ZN(n3450) );
  I_NAND2 U2822 ( .A1(n3454), .B1(n29428), .ZN(n3455) );
  I_NAND2 U2823 ( .A1(n3456), .B1(n29412), .ZN(n3457) );
  I_NAND2 U2824 ( .A1(n3458), .B1(n29407), .ZN(n3459) );
  I_NAND2 U2825 ( .A1(n3460), .B1(n29407), .ZN(n3461) );
  I_NAND2 U2826 ( .A1(n3462), .B1(n29407), .ZN(n3463) );
  I_NAND2 U2827 ( .A1(n3464), .B1(n29407), .ZN(n3465) );
  I_NAND2 U2828 ( .A1(n3466), .B1(n29408), .ZN(n3467) );
  I_NAND2 U2829 ( .A1(n3468), .B1(n29408), .ZN(n3469) );
  I_NAND2 U2830 ( .A1(n3470), .B1(n29408), .ZN(n3471) );
  I_NAND2 U2831 ( .A1(n3472), .B1(n29408), .ZN(n3473) );
  I_NAND2 U2832 ( .A1(n3474), .B1(n29408), .ZN(n3475) );
  I_NAND2 U2833 ( .A1(n3476), .B1(n29408), .ZN(n3477) );
  I_NAND2 U2834 ( .A1(n3478), .B1(n29408), .ZN(n3479) );
  I_NAND2 U2835 ( .A1(n3480), .B1(n29408), .ZN(n3481) );
  I_NAND2 U2836 ( .A1(n3482), .B1(n29408), .ZN(n3483) );
  I_NAND2 U2837 ( .A1(n3484), .B1(n29408), .ZN(n3485) );
  I_NAND2 U2838 ( .A1(n3486), .B1(n29408), .ZN(n3487) );
  I_NAND2 U2839 ( .A1(n3488), .B1(n29408), .ZN(n3489) );
  I_NAND2 U2840 ( .A1(n3490), .B1(n29409), .ZN(n3491) );
  I_NAND2 U2841 ( .A1(n3492), .B1(n29409), .ZN(n3493) );
  I_NAND2 U2842 ( .A1(n3494), .B1(n29409), .ZN(n3495) );
  I_NAND2 U2843 ( .A1(n3496), .B1(n29409), .ZN(n3497) );
  I_NAND2 U2844 ( .A1(n3498), .B1(n29409), .ZN(n3499) );
  I_NAND2 U2845 ( .A1(n3500), .B1(n29409), .ZN(n3501) );
  I_NAND2 U2846 ( .A1(n3502), .B1(n29409), .ZN(n3503) );
  I_NAND2 U2847 ( .A1(n3504), .B1(n29409), .ZN(n3505) );
  I_NAND2 U2848 ( .A1(n3506), .B1(n29409), .ZN(n3507) );
  I_NAND2 U2849 ( .A1(n3508), .B1(n29409), .ZN(n3509) );
  I_NAND2 U2850 ( .A1(n3510), .B1(n29409), .ZN(n3511) );
  I_NAND2 U2851 ( .A1(n3512), .B1(n29409), .ZN(n3513) );
  I_NAND2 U2852 ( .A1(n3514), .B1(n29410), .ZN(n3515) );
  I_NAND2 U2853 ( .A1(n3516), .B1(n29410), .ZN(n3517) );
  I_NAND2 U2854 ( .A1(n3518), .B1(n29410), .ZN(n3519) );
  I_NAND2 U2855 ( .A1(n3520), .B1(n29410), .ZN(n3521) );
  I_NAND2 U2856 ( .A1(n3522), .B1(n29410), .ZN(n3523) );
  I_NAND2 U2857 ( .A1(n3524), .B1(n29410), .ZN(n3525) );
  I_NAND2 U2858 ( .A1(n3526), .B1(n29410), .ZN(n3527) );
  I_NAND2 U2859 ( .A1(n3528), .B1(n29410), .ZN(n3529) );
  I_NAND2 U2860 ( .A1(n3530), .B1(n29410), .ZN(n3531) );
  I_NAND2 U2861 ( .A1(n3532), .B1(n29410), .ZN(n3533) );
  I_NAND2 U2862 ( .A1(n3534), .B1(n29410), .ZN(n3535) );
  I_NAND2 U2863 ( .A1(n3536), .B1(n29410), .ZN(n3537) );
  I_NAND2 U2864 ( .A1(n3538), .B1(n29411), .ZN(n3539) );
  I_NAND2 U2865 ( .A1(n3540), .B1(n29411), .ZN(n3541) );
  I_NAND2 U2866 ( .A1(n3542), .B1(n29411), .ZN(n3543) );
  I_NAND2 U2867 ( .A1(n3544), .B1(n29411), .ZN(n3545) );
  I_NAND2 U2868 ( .A1(n3546), .B1(n29411), .ZN(n3547) );
  I_NAND2 U2869 ( .A1(n3548), .B1(n29411), .ZN(n3549) );
  I_NAND2 U2870 ( .A1(n3550), .B1(n29411), .ZN(n3551) );
  I_NAND2 U2871 ( .A1(n3552), .B1(n29411), .ZN(n3553) );
  I_NAND2 U2872 ( .A1(n3554), .B1(n29411), .ZN(n3555) );
  I_NAND2 U2873 ( .A1(n3556), .B1(n29411), .ZN(n3557) );
  I_NAND2 U2874 ( .A1(n3558), .B1(n29411), .ZN(n3559) );
  I_NAND2 U2875 ( .A1(n3560), .B1(n29411), .ZN(n3561) );
  I_NAND2 U2876 ( .A1(n3562), .B1(n29412), .ZN(n3563) );
  I_NAND2 U2877 ( .A1(n3564), .B1(n29412), .ZN(n3565) );
  I_NAND2 U2878 ( .A1(n3566), .B1(n29412), .ZN(n3567) );
  I_NAND2 U2879 ( .A1(n3568), .B1(n29412), .ZN(n3569) );
  I_NAND2 U2880 ( .A1(n3570), .B1(n29412), .ZN(n3571) );
  I_NAND2 U2881 ( .A1(n3572), .B1(n29412), .ZN(n3573) );
  I_NAND2 U2882 ( .A1(n3574), .B1(n29412), .ZN(n3575) );
  I_NAND2 U2883 ( .A1(n3576), .B1(n29412), .ZN(n3577) );
  I_NAND2 U2884 ( .A1(n3578), .B1(n29412), .ZN(n3579) );
  I_NAND2 U2885 ( .A1(n3583), .B1(n29412), .ZN(n3584) );
  I_NAND2 U2886 ( .A1(n3585), .B1(n29413), .ZN(n3586) );
  I_NAND2 U2887 ( .A1(n3587), .B1(n29413), .ZN(n3588) );
  I_NAND2 U2888 ( .A1(n3589), .B1(n29413), .ZN(n3590) );
  I_NAND2 U2889 ( .A1(n3591), .B1(n29413), .ZN(n3592) );
  I_NAND2 U2890 ( .A1(n3593), .B1(n29413), .ZN(n3594) );
  I_NAND2 U2891 ( .A1(n3595), .B1(n29413), .ZN(n3596) );
  I_NAND2 U2892 ( .A1(n3597), .B1(n29413), .ZN(n3598) );
  I_NAND2 U2893 ( .A1(n3599), .B1(n29413), .ZN(n3600) );
  I_NAND2 U2894 ( .A1(n3601), .B1(n29413), .ZN(n3602) );
  I_NAND2 U2895 ( .A1(n3603), .B1(n29413), .ZN(n3604) );
  I_NAND2 U2896 ( .A1(n3605), .B1(n29413), .ZN(n3606) );
  I_NAND2 U2897 ( .A1(n3607), .B1(n29413), .ZN(n3608) );
  I_NAND2 U2898 ( .A1(n3609), .B1(n29414), .ZN(n3610) );
  I_NAND2 U2899 ( .A1(n3611), .B1(n29414), .ZN(n3612) );
  I_NAND2 U2900 ( .A1(n3613), .B1(n29414), .ZN(n3614) );
  I_NAND2 U2901 ( .A1(n3615), .B1(n29414), .ZN(n3616) );
  I_NAND2 U2902 ( .A1(n3617), .B1(n29414), .ZN(n3618) );
  I_NAND2 U2903 ( .A1(n3619), .B1(n29414), .ZN(n3620) );
  I_NAND2 U2904 ( .A1(n3621), .B1(n29414), .ZN(n3622) );
  I_NAND2 U2905 ( .A1(n3623), .B1(n29414), .ZN(n3624) );
  I_NAND2 U2906 ( .A1(n3625), .B1(n29414), .ZN(n3626) );
  I_NAND2 U2907 ( .A1(n3627), .B1(n29414), .ZN(n3628) );
  I_NAND2 U2908 ( .A1(n3629), .B1(n29414), .ZN(n3630) );
  I_NAND2 U2909 ( .A1(n3631), .B1(n29414), .ZN(n3632) );
  I_NAND2 U2910 ( .A1(n3633), .B1(n29415), .ZN(n3634) );
  I_NAND2 U2911 ( .A1(n3635), .B1(n29415), .ZN(n3636) );
  I_NAND2 U2912 ( .A1(n3637), .B1(n29415), .ZN(n3638) );
  I_NAND2 U2913 ( .A1(n3639), .B1(n29415), .ZN(n3640) );
  I_NAND2 U2914 ( .A1(n3641), .B1(n29415), .ZN(n3642) );
  I_NAND2 U2915 ( .A1(n3643), .B1(n29415), .ZN(n3644) );
  I_NAND2 U2916 ( .A1(n3645), .B1(n29415), .ZN(n3646) );
  I_NAND2 U2917 ( .A1(n3647), .B1(n29415), .ZN(n3648) );
  I_NAND2 U2918 ( .A1(n3649), .B1(n29415), .ZN(n3650) );
  I_NAND2 U2919 ( .A1(n3651), .B1(n29415), .ZN(n3652) );
  I_NAND2 U2920 ( .A1(n3653), .B1(n29415), .ZN(n3654) );
  I_NAND2 U2921 ( .A1(n3655), .B1(n29415), .ZN(n3656) );
  I_NAND2 U2922 ( .A1(n3657), .B1(n29416), .ZN(n3658) );
  I_NAND2 U2923 ( .A1(n3659), .B1(n29416), .ZN(n3660) );
  I_NAND2 U2924 ( .A1(n3661), .B1(n29416), .ZN(n3662) );
  I_NAND2 U2925 ( .A1(n3663), .B1(n29416), .ZN(n3664) );
  I_NAND2 U2926 ( .A1(n3665), .B1(n29416), .ZN(n3666) );
  I_NAND2 U2927 ( .A1(n3667), .B1(n29416), .ZN(n3668) );
  I_NAND2 U2928 ( .A1(n3669), .B1(n29416), .ZN(n3670) );
  I_NAND2 U2929 ( .A1(n3671), .B1(n29416), .ZN(n3672) );
  I_NAND2 U2930 ( .A1(n3673), .B1(n29416), .ZN(n3674) );
  I_NAND2 U2931 ( .A1(n3675), .B1(n29416), .ZN(n3676) );
  I_NAND2 U2932 ( .A1(n3677), .B1(n29416), .ZN(n3678) );
  I_NAND2 U2933 ( .A1(n3679), .B1(n29416), .ZN(n3680) );
  I_NAND2 U2934 ( .A1(n3681), .B1(n29417), .ZN(n3682) );
  I_NAND2 U2935 ( .A1(n3683), .B1(n29417), .ZN(n3684) );
  I_NAND2 U2936 ( .A1(n3685), .B1(n29417), .ZN(n3686) );
  I_NAND2 U2937 ( .A1(n3687), .B1(n29417), .ZN(n3688) );
  I_NAND2 U2938 ( .A1(n3689), .B1(n29417), .ZN(n3690) );
  I_NAND2 U2939 ( .A1(n3691), .B1(n29417), .ZN(n3692) );
  I_NAND2 U2940 ( .A1(n3693), .B1(n29417), .ZN(n3694) );
  I_NAND2 U2941 ( .A1(n3695), .B1(n29417), .ZN(n3696) );
  I_NAND2 U2942 ( .A1(n3697), .B1(n29417), .ZN(n3698) );
  I_NAND2 U2943 ( .A1(n3699), .B1(n29417), .ZN(n3700) );
  I_NAND2 U2944 ( .A1(n3701), .B1(n29417), .ZN(n3702) );
  I_NAND2 U2945 ( .A1(n3703), .B1(n29417), .ZN(n3704) );
  I_NAND2 U2946 ( .A1(n3705), .B1(n29418), .ZN(n3706) );
  I_NAND2 U2947 ( .A1(n3707), .B1(n29418), .ZN(n3708) );
  I_NAND2 U2948 ( .A1(n3712), .B1(n29444), .ZN(n3713) );
  I_NAND2 U2949 ( .A1(n3714), .B1(n29439), .ZN(n3715) );
  I_NAND2 U2950 ( .A1(n3716), .B1(n29439), .ZN(n3717) );
  I_NAND2 U2951 ( .A1(n3718), .B1(n29439), .ZN(n3719) );
  I_NAND2 U2952 ( .A1(n3720), .B1(n29439), .ZN(n3721) );
  I_NAND2 U2953 ( .A1(n3722), .B1(n29439), .ZN(n3723) );
  I_NAND2 U2954 ( .A1(n3724), .B1(n29450), .ZN(n3725) );
  I_NAND2 U2955 ( .A1(n3726), .B1(n29439), .ZN(n3727) );
  I_NAND2 U2956 ( .A1(n3728), .B1(n29440), .ZN(n3729) );
  I_NAND2 U2957 ( .A1(n3730), .B1(n29440), .ZN(n3731) );
  I_NAND2 U2958 ( .A1(n3732), .B1(n29440), .ZN(n3733) );
  I_NAND2 U2959 ( .A1(n3734), .B1(n29440), .ZN(n3735) );
  I_NAND2 U2960 ( .A1(n3736), .B1(n29440), .ZN(n3737) );
  I_NAND2 U2961 ( .A1(n3738), .B1(n29440), .ZN(n3739) );
  I_NAND2 U2962 ( .A1(n3740), .B1(n29440), .ZN(n3741) );
  I_NAND2 U2963 ( .A1(n3742), .B1(n29440), .ZN(n3743) );
  I_NAND2 U2964 ( .A1(n3744), .B1(n29440), .ZN(n3745) );
  I_NAND2 U2965 ( .A1(n3746), .B1(n29440), .ZN(n3747) );
  I_NAND2 U2966 ( .A1(n3748), .B1(n29440), .ZN(n3749) );
  I_NAND2 U2967 ( .A1(n3750), .B1(n29440), .ZN(n3751) );
  I_NAND2 U2968 ( .A1(n3752), .B1(n29441), .ZN(n3753) );
  I_NAND2 U2969 ( .A1(n3754), .B1(n29441), .ZN(n3755) );
  I_NAND2 U2970 ( .A1(n3756), .B1(n29441), .ZN(n3757) );
  I_NAND2 U2971 ( .A1(n3758), .B1(n29441), .ZN(n3759) );
  I_NAND2 U2972 ( .A1(n3760), .B1(n29441), .ZN(n3761) );
  I_NAND2 U2973 ( .A1(n3762), .B1(n29441), .ZN(n3763) );
  I_NAND2 U2974 ( .A1(n3764), .B1(n29441), .ZN(n3765) );
  I_NAND2 U2975 ( .A1(n3766), .B1(n29441), .ZN(n3767) );
  I_NAND2 U2976 ( .A1(n3768), .B1(n29441), .ZN(n3769) );
  I_NAND2 U2977 ( .A1(n3770), .B1(n29441), .ZN(n3771) );
  I_NAND2 U2978 ( .A1(n3772), .B1(n29441), .ZN(n3773) );
  I_NAND2 U2979 ( .A1(n3774), .B1(n29441), .ZN(n3775) );
  I_NAND2 U2980 ( .A1(n3776), .B1(n29442), .ZN(n3777) );
  I_NAND2 U2981 ( .A1(n3778), .B1(n29442), .ZN(n3779) );
  I_NAND2 U2982 ( .A1(n3780), .B1(n29442), .ZN(n3781) );
  I_NAND2 U2983 ( .A1(n3782), .B1(n29442), .ZN(n3783) );
  I_NAND2 U2984 ( .A1(n3784), .B1(n29442), .ZN(n3785) );
  I_NAND2 U2985 ( .A1(n3786), .B1(n29442), .ZN(n3787) );
  I_NAND2 U2986 ( .A1(n3788), .B1(n29442), .ZN(n3789) );
  I_NAND2 U2987 ( .A1(n3790), .B1(n29442), .ZN(n3791) );
  I_NAND2 U2988 ( .A1(n3792), .B1(n29442), .ZN(n3793) );
  I_NAND2 U2989 ( .A1(n3794), .B1(n29442), .ZN(n3795) );
  I_NAND2 U2990 ( .A1(n3796), .B1(n29442), .ZN(n3797) );
  I_NAND2 U2991 ( .A1(n3798), .B1(n29442), .ZN(n3799) );
  I_NAND2 U2992 ( .A1(n3800), .B1(n29443), .ZN(n3801) );
  I_NAND2 U2993 ( .A1(n3802), .B1(n29443), .ZN(n3803) );
  I_NAND2 U2994 ( .A1(n3804), .B1(n29443), .ZN(n3805) );
  I_NAND2 U2995 ( .A1(n3806), .B1(n29443), .ZN(n3807) );
  I_NAND2 U2996 ( .A1(n3808), .B1(n29443), .ZN(n3809) );
  I_NAND2 U2997 ( .A1(n3810), .B1(n29443), .ZN(n3811) );
  I_NAND2 U2998 ( .A1(n3812), .B1(n29443), .ZN(n3813) );
  I_NAND2 U2999 ( .A1(n3814), .B1(n29443), .ZN(n3815) );
  I_NAND2 U3000 ( .A1(n3816), .B1(n29443), .ZN(n3817) );
  I_NAND2 U3001 ( .A1(n3818), .B1(n29443), .ZN(n3819) );
  I_NAND2 U3002 ( .A1(n3820), .B1(n29443), .ZN(n3821) );
  I_NAND2 U3003 ( .A1(n3822), .B1(n29443), .ZN(n3823) );
  I_NAND2 U3004 ( .A1(n3824), .B1(n29444), .ZN(n3825) );
  I_NAND2 U3005 ( .A1(n3826), .B1(n29444), .ZN(n3827) );
  I_NAND2 U3006 ( .A1(n3828), .B1(n29444), .ZN(n3829) );
  I_NAND2 U3007 ( .A1(n3830), .B1(n29444), .ZN(n3831) );
  I_NAND2 U3008 ( .A1(n3832), .B1(n29444), .ZN(n3833) );
  I_NAND2 U3009 ( .A1(n3834), .B1(n29444), .ZN(n3835) );
  I_NAND2 U3010 ( .A1(n3836), .B1(n29444), .ZN(n3837) );
  I_NAND2 U3011 ( .A1(n3841), .B1(n29444), .ZN(n3842) );
  I_NAND2 U3012 ( .A1(n3843), .B1(n29444), .ZN(n3844) );
  I_NAND2 U3013 ( .A1(n3845), .B1(n29444), .ZN(n3846) );
  I_NAND2 U3014 ( .A1(n3847), .B1(n29445), .ZN(n3848) );
  I_NAND2 U3015 ( .A1(n3849), .B1(n29445), .ZN(n3850) );
  I_NAND2 U3016 ( .A1(n3851), .B1(n29445), .ZN(n3852) );
  I_NAND2 U3017 ( .A1(n3853), .B1(n29445), .ZN(n3854) );
  I_NAND2 U3018 ( .A1(n3855), .B1(n29445), .ZN(n3856) );
  I_NAND2 U3019 ( .A1(n3857), .B1(n29445), .ZN(n3858) );
  I_NAND2 U3020 ( .A1(n3859), .B1(n29445), .ZN(n3860) );
  I_NAND2 U3021 ( .A1(n3861), .B1(n29445), .ZN(n3862) );
  I_NAND2 U3022 ( .A1(n3863), .B1(n29445), .ZN(n3864) );
  I_NAND2 U3023 ( .A1(n3865), .B1(n29445), .ZN(n3866) );
  I_NAND2 U3024 ( .A1(n3867), .B1(n29445), .ZN(n3868) );
  I_NAND2 U3025 ( .A1(n3869), .B1(n29445), .ZN(n3870) );
  I_NAND2 U3026 ( .A1(n3871), .B1(n29446), .ZN(n3872) );
  I_NAND2 U3027 ( .A1(n3873), .B1(n29446), .ZN(n3874) );
  I_NAND2 U3028 ( .A1(n3875), .B1(n29446), .ZN(n3876) );
  I_NAND2 U3029 ( .A1(n3877), .B1(n29446), .ZN(n3878) );
  I_NAND2 U3030 ( .A1(n3879), .B1(n29446), .ZN(n3880) );
  I_NAND2 U3031 ( .A1(n3881), .B1(n29446), .ZN(n3882) );
  I_NAND2 U3032 ( .A1(n3883), .B1(n29446), .ZN(n3884) );
  I_NAND2 U3033 ( .A1(n3885), .B1(n29446), .ZN(n3886) );
  I_NAND2 U3034 ( .A1(n3887), .B1(n29446), .ZN(n3888) );
  I_NAND2 U3035 ( .A1(n3889), .B1(n29446), .ZN(n3890) );
  I_NAND2 U3036 ( .A1(n3891), .B1(n29446), .ZN(n3892) );
  I_NAND2 U3037 ( .A1(n3893), .B1(n29446), .ZN(n3894) );
  I_NAND2 U3038 ( .A1(n3895), .B1(n29447), .ZN(n3896) );
  I_NAND2 U3039 ( .A1(n3897), .B1(n29447), .ZN(n3898) );
  I_NAND2 U3040 ( .A1(n3899), .B1(n29447), .ZN(n3900) );
  I_NAND2 U3041 ( .A1(n3901), .B1(n29447), .ZN(n3902) );
  I_NAND2 U3042 ( .A1(n3903), .B1(n29447), .ZN(n3904) );
  I_NAND2 U3043 ( .A1(n3905), .B1(n29447), .ZN(n3906) );
  I_NAND2 U3044 ( .A1(n3907), .B1(n29447), .ZN(n3908) );
  I_NAND2 U3045 ( .A1(n3909), .B1(n29447), .ZN(n3910) );
  I_NAND2 U3046 ( .A1(n3911), .B1(n29447), .ZN(n3912) );
  I_NAND2 U3047 ( .A1(n3913), .B1(n29447), .ZN(n3914) );
  I_NAND2 U3048 ( .A1(n3915), .B1(n29447), .ZN(n3916) );
  I_NAND2 U3049 ( .A1(n3917), .B1(n29447), .ZN(n3918) );
  I_NAND2 U3050 ( .A1(n3919), .B1(n29448), .ZN(n3920) );
  I_NAND2 U3051 ( .A1(n3921), .B1(n29448), .ZN(n3922) );
  I_NAND2 U3052 ( .A1(n3923), .B1(n29448), .ZN(n3924) );
  I_NAND2 U3053 ( .A1(n3925), .B1(n29448), .ZN(n3926) );
  I_NAND2 U3054 ( .A1(n3927), .B1(n29448), .ZN(n3928) );
  I_NAND2 U3055 ( .A1(n3929), .B1(n29448), .ZN(n3930) );
  I_NAND2 U3056 ( .A1(n3931), .B1(n29448), .ZN(n3932) );
  I_NAND2 U3057 ( .A1(n3933), .B1(n29448), .ZN(n3934) );
  I_NAND2 U3058 ( .A1(n3935), .B1(n29448), .ZN(n3936) );
  I_NAND2 U3059 ( .A1(n3937), .B1(n29448), .ZN(n3938) );
  I_NAND2 U3060 ( .A1(n3939), .B1(n29448), .ZN(n3940) );
  I_NAND2 U3061 ( .A1(n3941), .B1(n29448), .ZN(n3942) );
  I_NAND2 U3062 ( .A1(n3943), .B1(n29449), .ZN(n3944) );
  I_NAND2 U3063 ( .A1(n3945), .B1(n29449), .ZN(n3946) );
  I_NAND2 U3064 ( .A1(n3947), .B1(n29449), .ZN(n3948) );
  I_NAND2 U3065 ( .A1(n3949), .B1(n29449), .ZN(n3950) );
  I_NAND2 U3066 ( .A1(n3951), .B1(n29449), .ZN(n3952) );
  I_NAND2 U3067 ( .A1(n3953), .B1(n29449), .ZN(n3954) );
  I_NAND2 U3068 ( .A1(n3955), .B1(n29449), .ZN(n3956) );
  I_NAND2 U3069 ( .A1(n3957), .B1(n29449), .ZN(n3958) );
  I_NAND2 U3070 ( .A1(n3959), .B1(n29449), .ZN(n3960) );
  I_NAND2 U3071 ( .A1(n3961), .B1(n29449), .ZN(n3962) );
  I_NAND2 U3072 ( .A1(n3963), .B1(n29449), .ZN(n3964) );
  I_NAND2 U3073 ( .A1(n3965), .B1(n29449), .ZN(n3966) );
  I_NAND2 U3074 ( .A1(n3970), .B1(n29434), .ZN(n3971) );
  I_NAND2 U3075 ( .A1(n3972), .B1(n29428), .ZN(n3973) );
  I_NAND2 U3076 ( .A1(n3974), .B1(n29429), .ZN(n3975) );
  I_NAND2 U3077 ( .A1(n3976), .B1(n29429), .ZN(n3977) );
  I_NAND2 U3078 ( .A1(n3978), .B1(n29429), .ZN(n3979) );
  I_NAND2 U3079 ( .A1(n3980), .B1(n29429), .ZN(n3981) );
  I_NAND2 U3080 ( .A1(n3982), .B1(n29429), .ZN(n3983) );
  I_NAND2 U3081 ( .A1(n3984), .B1(n29429), .ZN(n3985) );
  I_NAND2 U3082 ( .A1(n3986), .B1(n29429), .ZN(n3987) );
  I_NAND2 U3083 ( .A1(n3988), .B1(n29429), .ZN(n3989) );
  I_NAND2 U3084 ( .A1(n3990), .B1(n29429), .ZN(n3991) );
  I_NAND2 U3085 ( .A1(n3992), .B1(n29429), .ZN(n3993) );
  I_NAND2 U3086 ( .A1(n3994), .B1(n29429), .ZN(n3995) );
  I_NAND2 U3087 ( .A1(n3996), .B1(n29429), .ZN(n3997) );
  I_NAND2 U3088 ( .A1(n3998), .B1(n29430), .ZN(n3999) );
  I_NAND2 U3089 ( .A1(n4000), .B1(n29430), .ZN(n4001) );
  I_NAND2 U3090 ( .A1(n4002), .B1(n29430), .ZN(n4003) );
  I_NAND2 U3091 ( .A1(n4004), .B1(n29430), .ZN(n4005) );
  I_NAND2 U3092 ( .A1(n4006), .B1(n29430), .ZN(n4007) );
  I_NAND2 U3093 ( .A1(n4008), .B1(n29430), .ZN(n4009) );
  I_NAND2 U3094 ( .A1(n4010), .B1(n29430), .ZN(n4011) );
  I_NAND2 U3095 ( .A1(n4012), .B1(n29430), .ZN(n4013) );
  I_NAND2 U3096 ( .A1(n4014), .B1(n29430), .ZN(n4015) );
  I_NAND2 U3097 ( .A1(n4016), .B1(n29430), .ZN(n4017) );
  I_NAND2 U3098 ( .A1(n4018), .B1(n29430), .ZN(n4019) );
  I_NAND2 U3099 ( .A1(n4020), .B1(n29430), .ZN(n4021) );
  I_NAND2 U3100 ( .A1(n4022), .B1(n29431), .ZN(n4023) );
  I_NAND2 U3101 ( .A1(n4024), .B1(n29431), .ZN(n4025) );
  I_NAND2 U3102 ( .A1(n4026), .B1(n29431), .ZN(n4027) );
  I_NAND2 U3103 ( .A1(n4028), .B1(n29431), .ZN(n4029) );
  I_NAND2 U3104 ( .A1(n4030), .B1(n29431), .ZN(n4031) );
  I_NAND2 U3105 ( .A1(n4032), .B1(n29431), .ZN(n4033) );
  I_NAND2 U3106 ( .A1(n4034), .B1(n29431), .ZN(n4035) );
  I_NAND2 U3107 ( .A1(n4036), .B1(n29431), .ZN(n4037) );
  I_NAND2 U3108 ( .A1(n4038), .B1(n29431), .ZN(n4039) );
  I_NAND2 U3109 ( .A1(n4040), .B1(n29431), .ZN(n4041) );
  I_NAND2 U3110 ( .A1(n4042), .B1(n29431), .ZN(n4043) );
  I_NAND2 U3111 ( .A1(n4044), .B1(n29431), .ZN(n4045) );
  I_NAND2 U3112 ( .A1(n4046), .B1(n29432), .ZN(n4047) );
  I_NAND2 U3113 ( .A1(n4048), .B1(n29432), .ZN(n4049) );
  I_NAND2 U3114 ( .A1(n4050), .B1(n29432), .ZN(n4051) );
  I_NAND2 U3115 ( .A1(n4052), .B1(n29432), .ZN(n4053) );
  I_NAND2 U3116 ( .A1(n4054), .B1(n29432), .ZN(n4055) );
  I_NAND2 U3117 ( .A1(n4056), .B1(n29432), .ZN(n4057) );
  I_NAND2 U3118 ( .A1(n4058), .B1(n29432), .ZN(n4059) );
  I_NAND2 U3119 ( .A1(n4060), .B1(n29432), .ZN(n4061) );
  I_NAND2 U3120 ( .A1(n4062), .B1(n29432), .ZN(n4063) );
  I_NAND2 U3121 ( .A1(n4064), .B1(n29432), .ZN(n4065) );
  I_NAND2 U3122 ( .A1(n4066), .B1(n29432), .ZN(n4067) );
  I_NAND2 U3123 ( .A1(n4068), .B1(n29432), .ZN(n4069) );
  I_NAND2 U3124 ( .A1(n4070), .B1(n29433), .ZN(n4071) );
  I_NAND2 U3125 ( .A1(n4072), .B1(n29433), .ZN(n4073) );
  I_NAND2 U3126 ( .A1(n4074), .B1(n29433), .ZN(n4075) );
  I_NAND2 U3127 ( .A1(n4076), .B1(n29433), .ZN(n4077) );
  I_NAND2 U3128 ( .A1(n4078), .B1(n29433), .ZN(n4079) );
  I_NAND2 U3129 ( .A1(n4080), .B1(n29433), .ZN(n4081) );
  I_NAND2 U3130 ( .A1(n4082), .B1(n29433), .ZN(n4083) );
  I_NAND2 U3131 ( .A1(n4084), .B1(n29433), .ZN(n4085) );
  I_NAND2 U3132 ( .A1(n4086), .B1(n29433), .ZN(n4087) );
  I_NAND2 U3133 ( .A1(n4088), .B1(n29433), .ZN(n4089) );
  I_NAND2 U3134 ( .A1(n4090), .B1(n29433), .ZN(n4091) );
  I_NAND2 U3135 ( .A1(n4092), .B1(n29433), .ZN(n4093) );
  I_NAND2 U3136 ( .A1(n4094), .B1(n29434), .ZN(n4095) );
  I_NAND2 U3137 ( .A1(n4101), .B1(n29434), .ZN(n4102) );
  I_NAND2 U3138 ( .A1(n4104), .B1(n29434), .ZN(n4105) );
  I_NAND2 U3139 ( .A1(n4107), .B1(n29434), .ZN(n4108) );
  I_NAND2 U3140 ( .A1(n4110), .B1(n29434), .ZN(n4111) );
  I_NAND2 U3141 ( .A1(n4113), .B1(n29434), .ZN(n4114) );
  I_NAND2 U3142 ( .A1(n4116), .B1(n29434), .ZN(n4117) );
  I_NAND2 U3143 ( .A1(n4119), .B1(n29434), .ZN(n4120) );
  I_NAND2 U3144 ( .A1(n4122), .B1(n29434), .ZN(n4123) );
  I_NAND2 U3145 ( .A1(n4125), .B1(n29434), .ZN(n4126) );
  I_NAND2 U3146 ( .A1(n4127), .B1(n29435), .ZN(n4128) );
  I_NAND2 U3147 ( .A1(n4129), .B1(n29435), .ZN(n4130) );
  I_NAND2 U3148 ( .A1(n4131), .B1(n29435), .ZN(n4132) );
  I_NAND2 U3149 ( .A1(n4133), .B1(n29435), .ZN(n4134) );
  I_NAND2 U3150 ( .A1(n4135), .B1(n29435), .ZN(n4136) );
  I_NAND2 U3151 ( .A1(n4137), .B1(n29435), .ZN(n4138) );
  I_NAND2 U3152 ( .A1(n4139), .B1(n29435), .ZN(n4140) );
  I_NAND2 U3153 ( .A1(n4142), .B1(n29435), .ZN(n4143) );
  I_NAND2 U3154 ( .A1(n4144), .B1(n29435), .ZN(n4145) );
  I_NAND2 U3155 ( .A1(n4146), .B1(n29435), .ZN(n4147) );
  I_NAND2 U3156 ( .A1(n4148), .B1(n29435), .ZN(n4149) );
  I_NAND2 U3157 ( .A1(n4150), .B1(n29435), .ZN(n4151) );
  I_NAND2 U3158 ( .A1(n4152), .B1(n29436), .ZN(n4153) );
  I_NAND2 U3159 ( .A1(n4154), .B1(n29436), .ZN(n4155) );
  I_NAND2 U3160 ( .A1(n4156), .B1(n29436), .ZN(n4157) );
  I_NAND2 U3161 ( .A1(n4159), .B1(n29436), .ZN(n4160) );
  I_NAND2 U3162 ( .A1(n4161), .B1(n29436), .ZN(n4162) );
  I_NAND2 U3163 ( .A1(n4163), .B1(n29436), .ZN(n4164) );
  I_NAND2 U3164 ( .A1(n4165), .B1(n29436), .ZN(n4166) );
  I_NAND2 U3165 ( .A1(n4167), .B1(n29436), .ZN(n4168) );
  I_NAND2 U3166 ( .A1(n4169), .B1(n29436), .ZN(n4170) );
  I_NAND2 U3167 ( .A1(n4171), .B1(n29436), .ZN(n4172) );
  I_NAND2 U3168 ( .A1(n4173), .B1(n29436), .ZN(n4174) );
  I_NAND2 U3169 ( .A1(n4176), .B1(n29436), .ZN(n4177) );
  I_NAND2 U3170 ( .A1(n4178), .B1(n29437), .ZN(n4179) );
  I_NAND2 U3171 ( .A1(n4180), .B1(n29437), .ZN(n4181) );
  I_NAND2 U3172 ( .A1(n4182), .B1(n29437), .ZN(n4183) );
  I_NAND2 U3173 ( .A1(n4184), .B1(n29437), .ZN(n4185) );
  I_NAND2 U3174 ( .A1(n4186), .B1(n29437), .ZN(n4187) );
  I_NAND2 U3175 ( .A1(n4188), .B1(n29437), .ZN(n4189) );
  I_NAND2 U3176 ( .A1(n4190), .B1(n29437), .ZN(n4191) );
  I_NAND2 U3177 ( .A1(n4193), .B1(n29437), .ZN(n4194) );
  I_NAND2 U3178 ( .A1(n4195), .B1(n29437), .ZN(n4196) );
  I_NAND2 U3179 ( .A1(n4197), .B1(n29437), .ZN(n4198) );
  I_NAND2 U3180 ( .A1(n4199), .B1(n29437), .ZN(n4200) );
  I_NAND2 U3181 ( .A1(n4201), .B1(n29437), .ZN(n4202) );
  I_NAND2 U3182 ( .A1(n4203), .B1(n29438), .ZN(n4204) );
  I_NAND2 U3183 ( .A1(n4205), .B1(n29438), .ZN(n4206) );
  I_NAND2 U3184 ( .A1(n4207), .B1(n29438), .ZN(n4208) );
  I_NAND2 U3185 ( .A1(n4210), .B1(n29438), .ZN(n4211) );
  I_NAND2 U3186 ( .A1(n4212), .B1(n29438), .ZN(n4213) );
  I_NAND2 U3187 ( .A1(n4214), .B1(n29438), .ZN(n4215) );
  I_NAND2 U3188 ( .A1(n4216), .B1(n29438), .ZN(n4217) );
  I_NAND2 U3189 ( .A1(n4218), .B1(n29438), .ZN(n4219) );
  I_NAND2 U3190 ( .A1(n4220), .B1(n29438), .ZN(n4221) );
  I_NAND2 U3191 ( .A1(n4222), .B1(n29438), .ZN(n4223) );
  I_NAND2 U3192 ( .A1(n4224), .B1(n29438), .ZN(n4225) );
  I_NAND2 U3193 ( .A1(n4227), .B1(n29438), .ZN(n4228) );
  I_NAND2 U3194 ( .A1(n4229), .B1(n29439), .ZN(n4230) );
  I_NAND2 U3195 ( .A1(n4231), .B1(n29439), .ZN(n4232) );
  I_NAND2 U3196 ( .A1(n4233), .B1(n29439), .ZN(n4234) );
  I_NAND2 U3197 ( .A1(n4235), .B1(n29439), .ZN(n4236) );
  I_NAND2 U3198 ( .A1(n4237), .B1(n29439), .ZN(n4238) );
  NAND2 U3199 ( .A1(n27431), .A2(n23), .ZN(n216) );
  NAND2 U3200 ( .A1(n27431), .A2(n5), .ZN(n219) );
  NAND2 U3201 ( .A1(n27431), .A2(n6), .ZN(n221) );
  NAND2 U3202 ( .A1(n27431), .A2(n7), .ZN(n223) );
  NAND2 U3203 ( .A1(n27431), .A2(n8), .ZN(n225) );
  NAND2 U3204 ( .A1(n27431), .A2(n9), .ZN(n227) );
  NAND2 U3205 ( .A1(n27431), .A2(n42), .ZN(n229) );
  NAND2 U3206 ( .A1(n27431), .A2(n45), .ZN(n231) );
  NAND2 U3207 ( .A1(n27431), .A2(n48), .ZN(n233) );
  NAND2 U3208 ( .A1(n27431), .A2(n51), .ZN(n235) );
  NAND2 U3209 ( .A1(n27431), .A2(n54), .ZN(n237) );
  NAND2 U3210 ( .A1(n27431), .A2(n57), .ZN(n239) );
  NAND2 U3211 ( .A1(n27432), .A2(n60), .ZN(n241) );
  NAND2 U3212 ( .A1(n27432), .A2(n63), .ZN(n243) );
  NAND2 U3213 ( .A1(n27433), .A2(n66), .ZN(n245) );
  NAND2 U3214 ( .A1(n27431), .A2(n69), .ZN(n247) );
  NAND2 U3215 ( .A1(n27433), .A2(n72), .ZN(n249) );
  NAND2 U3216 ( .A1(n27432), .A2(n75), .ZN(n251) );
  NAND2 U3217 ( .A1(n27433), .A2(n78), .ZN(n253) );
  NAND2 U3218 ( .A1(n27431), .A2(n81), .ZN(n255) );
  NAND2 U3219 ( .A1(n27431), .A2(n84), .ZN(n257) );
  NAND2 U3220 ( .A1(n27432), .A2(n87), .ZN(n259) );
  NAND2 U3221 ( .A1(n27433), .A2(n90), .ZN(n261) );
  NAND2 U3222 ( .A1(n27431), .A2(n93), .ZN(n263) );
  NAND2 U3223 ( .A1(n27432), .A2(n96), .ZN(n265) );
  NAND2 U3224 ( .A1(n27432), .A2(n99), .ZN(n267) );
  NAND2 U3225 ( .A1(n27432), .A2(n102), .ZN(n269) );
  NAND2 U3226 ( .A1(n27432), .A2(n105), .ZN(n271) );
  NAND2 U3227 ( .A1(n27432), .A2(n108), .ZN(n273) );
  NAND2 U3228 ( .A1(n27432), .A2(n111), .ZN(n275) );
  NAND2 U3229 ( .A1(n27432), .A2(n114), .ZN(n277) );
  NAND2 U3230 ( .A1(n27432), .A2(n117), .ZN(n279) );
  NAND2 U3231 ( .A1(n27432), .A2(n120), .ZN(n281) );
  NAND2 U3232 ( .A1(n27432), .A2(n123), .ZN(n283) );
  NAND2 U3233 ( .A1(n27432), .A2(n126), .ZN(n285) );
  NAND2 U3234 ( .A1(n27432), .A2(n129), .ZN(n287) );
  NAND2 U3235 ( .A1(n27433), .A2(n132), .ZN(n289) );
  NAND2 U3236 ( .A1(n27433), .A2(n135), .ZN(n291) );
  NAND2 U3237 ( .A1(n27433), .A2(n138), .ZN(n293) );
  NAND2 U3238 ( .A1(n27433), .A2(n141), .ZN(n295) );
  NAND2 U3239 ( .A1(n27433), .A2(n144), .ZN(n297) );
  NAND2 U3240 ( .A1(n27433), .A2(n147), .ZN(n299) );
  NAND2 U3241 ( .A1(n27433), .A2(n150), .ZN(n301) );
  NAND2 U3242 ( .A1(n27433), .A2(n153), .ZN(n303) );
  NAND2 U3243 ( .A1(n27433), .A2(n156), .ZN(n305) );
  NAND2 U3244 ( .A1(n27433), .A2(n159), .ZN(n307) );
  NAND2 U3245 ( .A1(n27433), .A2(n162), .ZN(n309) );
  NAND2 U3246 ( .A1(n27433), .A2(n165), .ZN(n311) );
  NAND2 U3247 ( .A1(n27433), .A2(n10), .ZN(n313) );
  NAND2 U3248 ( .A1(n27431), .A2(n11), .ZN(n315) );
  NAND2 U3249 ( .A1(n27432), .A2(n12), .ZN(n317) );
  NAND2 U3250 ( .A1(n27433), .A2(n24), .ZN(n319) );
  NAND2 U3251 ( .A1(n27431), .A2(n27), .ZN(n321) );
  NAND2 U3252 ( .A1(n27432), .A2(n30), .ZN(n323) );
  NAND2 U3253 ( .A1(n27433), .A2(n33), .ZN(n325) );
  NAND2 U3254 ( .A1(n27431), .A2(n36), .ZN(n327) );
  NAND2 U3255 ( .A1(n27432), .A2(n39), .ZN(n329) );
  NAND2 U3256 ( .A1(n27433), .A2(n168), .ZN(n331) );
  NAND2 U3257 ( .A1(n27431), .A2(n171), .ZN(n333) );
  NAND2 U3258 ( .A1(n27432), .A2(n174), .ZN(n335) );
  NAND2 U3259 ( .A1(n27428), .A2(n23), .ZN(n346) );
  NAND2 U3260 ( .A1(n27428), .A2(n5), .ZN(n349) );
  NAND2 U3261 ( .A1(n27428), .A2(n6), .ZN(n351) );
  NAND2 U3262 ( .A1(n27428), .A2(n7), .ZN(n353) );
  NAND2 U3263 ( .A1(n27428), .A2(n8), .ZN(n355) );
  NAND2 U3264 ( .A1(n27428), .A2(n9), .ZN(n357) );
  NAND2 U3265 ( .A1(n27428), .A2(n42), .ZN(n359) );
  NAND2 U3266 ( .A1(n27428), .A2(n45), .ZN(n361) );
  NAND2 U3267 ( .A1(n27428), .A2(n48), .ZN(n363) );
  NAND2 U3268 ( .A1(n27428), .A2(n51), .ZN(n365) );
  NAND2 U3269 ( .A1(n27428), .A2(n54), .ZN(n367) );
  NAND2 U3270 ( .A1(n27428), .A2(n57), .ZN(n369) );
  NAND2 U3271 ( .A1(n27429), .A2(n60), .ZN(n371) );
  NAND2 U3272 ( .A1(n27429), .A2(n63), .ZN(n373) );
  NAND2 U3273 ( .A1(n27430), .A2(n66), .ZN(n375) );
  NAND2 U3274 ( .A1(n27428), .A2(n69), .ZN(n377) );
  NAND2 U3275 ( .A1(n27430), .A2(n72), .ZN(n379) );
  NAND2 U3276 ( .A1(n27429), .A2(n75), .ZN(n381) );
  NAND2 U3277 ( .A1(n27430), .A2(n78), .ZN(n383) );
  NAND2 U3278 ( .A1(n27428), .A2(n81), .ZN(n385) );
  NAND2 U3279 ( .A1(n27428), .A2(n84), .ZN(n387) );
  NAND2 U3280 ( .A1(n27429), .A2(n87), .ZN(n389) );
  NAND2 U3281 ( .A1(n27430), .A2(n90), .ZN(n391) );
  NAND2 U3282 ( .A1(n27428), .A2(n93), .ZN(n393) );
  NAND2 U3283 ( .A1(n27429), .A2(n96), .ZN(n395) );
  NAND2 U3284 ( .A1(n27429), .A2(n99), .ZN(n397) );
  NAND2 U3285 ( .A1(n27429), .A2(n102), .ZN(n399) );
  NAND2 U3286 ( .A1(n27429), .A2(n105), .ZN(n401) );
  NAND2 U3287 ( .A1(n27429), .A2(n108), .ZN(n403) );
  NAND2 U3288 ( .A1(n27429), .A2(n111), .ZN(n405) );
  NAND2 U3289 ( .A1(n27429), .A2(n114), .ZN(n407) );
  NAND2 U3290 ( .A1(n27429), .A2(n117), .ZN(n409) );
  NAND2 U3291 ( .A1(n27429), .A2(n120), .ZN(n411) );
  NAND2 U3292 ( .A1(n27429), .A2(n123), .ZN(n413) );
  NAND2 U3293 ( .A1(n27429), .A2(n126), .ZN(n415) );
  NAND2 U3294 ( .A1(n27429), .A2(n129), .ZN(n417) );
  NAND2 U3295 ( .A1(n27430), .A2(n132), .ZN(n419) );
  NAND2 U3296 ( .A1(n27430), .A2(n135), .ZN(n421) );
  NAND2 U3297 ( .A1(n27430), .A2(n138), .ZN(n423) );
  NAND2 U3298 ( .A1(n27430), .A2(n141), .ZN(n425) );
  NAND2 U3299 ( .A1(n27430), .A2(n144), .ZN(n427) );
  NAND2 U3300 ( .A1(n27430), .A2(n147), .ZN(n429) );
  NAND2 U3301 ( .A1(n27430), .A2(n150), .ZN(n431) );
  NAND2 U3302 ( .A1(n27430), .A2(n153), .ZN(n433) );
  NAND2 U3303 ( .A1(n27430), .A2(n156), .ZN(n435) );
  NAND2 U3304 ( .A1(n27430), .A2(n159), .ZN(n437) );
  NAND2 U3305 ( .A1(n27430), .A2(n162), .ZN(n439) );
  NAND2 U3306 ( .A1(n27430), .A2(n165), .ZN(n441) );
  NAND2 U3307 ( .A1(n27430), .A2(n10), .ZN(n443) );
  NAND2 U3308 ( .A1(n27428), .A2(n11), .ZN(n445) );
  NAND2 U3309 ( .A1(n27429), .A2(n12), .ZN(n447) );
  NAND2 U3310 ( .A1(n27430), .A2(n24), .ZN(n449) );
  NAND2 U3311 ( .A1(n27428), .A2(n27), .ZN(n451) );
  NAND2 U3312 ( .A1(n27429), .A2(n30), .ZN(n453) );
  NAND2 U3313 ( .A1(n27430), .A2(n33), .ZN(n455) );
  NAND2 U3314 ( .A1(n27428), .A2(n36), .ZN(n457) );
  NAND2 U3315 ( .A1(n27429), .A2(n39), .ZN(n459) );
  NAND2 U3316 ( .A1(n27430), .A2(n168), .ZN(n461) );
  NAND2 U3317 ( .A1(n27428), .A2(n171), .ZN(n463) );
  NAND2 U3318 ( .A1(n27429), .A2(n174), .ZN(n465) );
  NAND2 U3319 ( .A1(n27425), .A2(n23), .ZN(n476) );
  NAND2 U3320 ( .A1(n27425), .A2(n5), .ZN(n479) );
  NAND2 U3321 ( .A1(n27425), .A2(n6), .ZN(n481) );
  NAND2 U3322 ( .A1(n27425), .A2(n7), .ZN(n483) );
  NAND2 U3323 ( .A1(n27425), .A2(n8), .ZN(n485) );
  NAND2 U3324 ( .A1(n27425), .A2(n9), .ZN(n487) );
  NAND2 U3325 ( .A1(n27425), .A2(n42), .ZN(n489) );
  NAND2 U3326 ( .A1(n27425), .A2(n45), .ZN(n491) );
  NAND2 U3327 ( .A1(n27425), .A2(n48), .ZN(n493) );
  NAND2 U3328 ( .A1(n27425), .A2(n51), .ZN(n495) );
  NAND2 U3329 ( .A1(n27425), .A2(n54), .ZN(n497) );
  NAND2 U3330 ( .A1(n27425), .A2(n57), .ZN(n499) );
  NAND2 U3331 ( .A1(n27426), .A2(n60), .ZN(n501) );
  NAND2 U3332 ( .A1(n27426), .A2(n63), .ZN(n503) );
  NAND2 U3333 ( .A1(n27427), .A2(n66), .ZN(n505) );
  NAND2 U3334 ( .A1(n27425), .A2(n69), .ZN(n507) );
  NAND2 U3335 ( .A1(n27427), .A2(n72), .ZN(n509) );
  NAND2 U3336 ( .A1(n27426), .A2(n75), .ZN(n511) );
  NAND2 U3337 ( .A1(n27427), .A2(n78), .ZN(n513) );
  NAND2 U3338 ( .A1(n27425), .A2(n81), .ZN(n515) );
  NAND2 U3339 ( .A1(n27425), .A2(n84), .ZN(n517) );
  NAND2 U3340 ( .A1(n27426), .A2(n87), .ZN(n519) );
  NAND2 U3341 ( .A1(n27427), .A2(n90), .ZN(n521) );
  NAND2 U3342 ( .A1(n27425), .A2(n93), .ZN(n523) );
  NAND2 U3343 ( .A1(n27426), .A2(n96), .ZN(n525) );
  NAND2 U3344 ( .A1(n27426), .A2(n99), .ZN(n527) );
  NAND2 U3345 ( .A1(n27426), .A2(n102), .ZN(n529) );
  NAND2 U3346 ( .A1(n27426), .A2(n105), .ZN(n531) );
  NAND2 U3347 ( .A1(n27426), .A2(n108), .ZN(n533) );
  NAND2 U3348 ( .A1(n27426), .A2(n111), .ZN(n535) );
  NAND2 U3349 ( .A1(n27426), .A2(n114), .ZN(n537) );
  NAND2 U3350 ( .A1(n27426), .A2(n117), .ZN(n539) );
  NAND2 U3351 ( .A1(n27426), .A2(n120), .ZN(n541) );
  NAND2 U3352 ( .A1(n27426), .A2(n123), .ZN(n543) );
  NAND2 U3353 ( .A1(n27426), .A2(n126), .ZN(n545) );
  NAND2 U3354 ( .A1(n27426), .A2(n129), .ZN(n547) );
  NAND2 U3355 ( .A1(n27427), .A2(n132), .ZN(n549) );
  NAND2 U3356 ( .A1(n27427), .A2(n135), .ZN(n551) );
  NAND2 U3357 ( .A1(n27427), .A2(n138), .ZN(n553) );
  NAND2 U3358 ( .A1(n27427), .A2(n141), .ZN(n555) );
  NAND2 U3359 ( .A1(n27427), .A2(n144), .ZN(n557) );
  NAND2 U3360 ( .A1(n27427), .A2(n147), .ZN(n559) );
  NAND2 U3361 ( .A1(n27427), .A2(n150), .ZN(n561) );
  NAND2 U3362 ( .A1(n27427), .A2(n153), .ZN(n563) );
  NAND2 U3363 ( .A1(n27427), .A2(n156), .ZN(n565) );
  NAND2 U3364 ( .A1(n27427), .A2(n159), .ZN(n567) );
  NAND2 U3365 ( .A1(n27427), .A2(n162), .ZN(n569) );
  NAND2 U3366 ( .A1(n27427), .A2(n165), .ZN(n571) );
  NAND2 U3367 ( .A1(n27427), .A2(n10), .ZN(n573) );
  NAND2 U3368 ( .A1(n27425), .A2(n11), .ZN(n575) );
  NAND2 U3369 ( .A1(n27426), .A2(n12), .ZN(n577) );
  NAND2 U3370 ( .A1(n27427), .A2(n24), .ZN(n579) );
  NAND2 U3371 ( .A1(n27425), .A2(n27), .ZN(n581) );
  NAND2 U3372 ( .A1(n27426), .A2(n30), .ZN(n583) );
  NAND2 U3373 ( .A1(n27427), .A2(n33), .ZN(n585) );
  NAND2 U3374 ( .A1(n27425), .A2(n36), .ZN(n587) );
  NAND2 U3375 ( .A1(n27426), .A2(n39), .ZN(n589) );
  NAND2 U3376 ( .A1(n27427), .A2(n168), .ZN(n591) );
  NAND2 U3377 ( .A1(n27425), .A2(n171), .ZN(n593) );
  NAND2 U3378 ( .A1(n27426), .A2(n174), .ZN(n595) );
  NAND2 U3379 ( .A1(n27422), .A2(n23), .ZN(n606) );
  NAND2 U3380 ( .A1(n27422), .A2(n5), .ZN(n609) );
  NAND2 U3381 ( .A1(n27422), .A2(n6), .ZN(n611) );
  NAND2 U3382 ( .A1(n27422), .A2(n7), .ZN(n613) );
  NAND2 U3383 ( .A1(n27422), .A2(n8), .ZN(n615) );
  NAND2 U3384 ( .A1(n27422), .A2(n9), .ZN(n617) );
  NAND2 U3385 ( .A1(n27422), .A2(n42), .ZN(n619) );
  NAND2 U3386 ( .A1(n27422), .A2(n45), .ZN(n621) );
  NAND2 U3387 ( .A1(n27422), .A2(n48), .ZN(n623) );
  NAND2 U3388 ( .A1(n27422), .A2(n51), .ZN(n625) );
  NAND2 U3389 ( .A1(n27422), .A2(n54), .ZN(n627) );
  NAND2 U3390 ( .A1(n27422), .A2(n57), .ZN(n629) );
  NAND2 U3391 ( .A1(n27423), .A2(n60), .ZN(n631) );
  NAND2 U3392 ( .A1(n27423), .A2(n63), .ZN(n633) );
  NAND2 U3393 ( .A1(n27424), .A2(n66), .ZN(n635) );
  NAND2 U3394 ( .A1(n27422), .A2(n69), .ZN(n637) );
  NAND2 U3395 ( .A1(n27424), .A2(n72), .ZN(n639) );
  NAND2 U3396 ( .A1(n27423), .A2(n75), .ZN(n641) );
  NAND2 U3397 ( .A1(n27424), .A2(n78), .ZN(n643) );
  NAND2 U3398 ( .A1(n27422), .A2(n81), .ZN(n645) );
  NAND2 U3399 ( .A1(n27422), .A2(n84), .ZN(n647) );
  NAND2 U3400 ( .A1(n27423), .A2(n87), .ZN(n649) );
  NAND2 U3401 ( .A1(n27424), .A2(n90), .ZN(n651) );
  NAND2 U3402 ( .A1(n27422), .A2(n93), .ZN(n653) );
  NAND2 U3403 ( .A1(n27423), .A2(n96), .ZN(n655) );
  NAND2 U3404 ( .A1(n27423), .A2(n99), .ZN(n657) );
  NAND2 U3405 ( .A1(n27423), .A2(n102), .ZN(n659) );
  NAND2 U3406 ( .A1(n27423), .A2(n105), .ZN(n661) );
  NAND2 U3407 ( .A1(n27423), .A2(n108), .ZN(n663) );
  NAND2 U3408 ( .A1(n27423), .A2(n111), .ZN(n665) );
  NAND2 U3409 ( .A1(n27423), .A2(n114), .ZN(n667) );
  NAND2 U3410 ( .A1(n27423), .A2(n117), .ZN(n669) );
  NAND2 U3411 ( .A1(n27423), .A2(n120), .ZN(n671) );
  NAND2 U3412 ( .A1(n27423), .A2(n123), .ZN(n673) );
  NAND2 U3413 ( .A1(n27423), .A2(n126), .ZN(n675) );
  NAND2 U3414 ( .A1(n27423), .A2(n129), .ZN(n677) );
  NAND2 U3415 ( .A1(n27424), .A2(n132), .ZN(n679) );
  NAND2 U3416 ( .A1(n27424), .A2(n135), .ZN(n681) );
  NAND2 U3417 ( .A1(n27424), .A2(n138), .ZN(n683) );
  NAND2 U3418 ( .A1(n27424), .A2(n141), .ZN(n685) );
  NAND2 U3419 ( .A1(n27424), .A2(n144), .ZN(n687) );
  NAND2 U3420 ( .A1(n27424), .A2(n147), .ZN(n689) );
  NAND2 U3421 ( .A1(n27424), .A2(n150), .ZN(n691) );
  NAND2 U3422 ( .A1(n27424), .A2(n153), .ZN(n693) );
  NAND2 U3423 ( .A1(n27424), .A2(n156), .ZN(n695) );
  NAND2 U3424 ( .A1(n27424), .A2(n159), .ZN(n697) );
  NAND2 U3425 ( .A1(n27424), .A2(n162), .ZN(n699) );
  NAND2 U3426 ( .A1(n27424), .A2(n165), .ZN(n701) );
  NAND2 U3427 ( .A1(n27424), .A2(n10), .ZN(n703) );
  NAND2 U3428 ( .A1(n27422), .A2(n11), .ZN(n705) );
  NAND2 U3429 ( .A1(n27423), .A2(n12), .ZN(n707) );
  NAND2 U3430 ( .A1(n27424), .A2(n24), .ZN(n709) );
  NAND2 U3431 ( .A1(n27422), .A2(n27), .ZN(n711) );
  NAND2 U3432 ( .A1(n27423), .A2(n30), .ZN(n713) );
  NAND2 U3433 ( .A1(n27424), .A2(n33), .ZN(n715) );
  NAND2 U3434 ( .A1(n27422), .A2(n36), .ZN(n717) );
  NAND2 U3435 ( .A1(n27423), .A2(n39), .ZN(n719) );
  NAND2 U3436 ( .A1(n27424), .A2(n168), .ZN(n721) );
  NAND2 U3437 ( .A1(n27422), .A2(n171), .ZN(n723) );
  NAND2 U3438 ( .A1(n27423), .A2(n174), .ZN(n725) );
  NAND2 U3439 ( .A1(n27419), .A2(n23), .ZN(n736) );
  NAND2 U3440 ( .A1(n27419), .A2(n5), .ZN(n739) );
  NAND2 U3441 ( .A1(n27419), .A2(n6), .ZN(n741) );
  NAND2 U3442 ( .A1(n27419), .A2(n7), .ZN(n743) );
  NAND2 U3443 ( .A1(n27419), .A2(n8), .ZN(n745) );
  NAND2 U3444 ( .A1(n27419), .A2(n9), .ZN(n747) );
  NAND2 U3445 ( .A1(n27419), .A2(n42), .ZN(n749) );
  NAND2 U3446 ( .A1(n27419), .A2(n45), .ZN(n751) );
  NAND2 U3447 ( .A1(n27419), .A2(n48), .ZN(n753) );
  NAND2 U3448 ( .A1(n27419), .A2(n51), .ZN(n755) );
  NAND2 U3449 ( .A1(n27419), .A2(n54), .ZN(n757) );
  NAND2 U3450 ( .A1(n27419), .A2(n57), .ZN(n759) );
  NAND2 U3451 ( .A1(n27420), .A2(n60), .ZN(n761) );
  NAND2 U3452 ( .A1(n27420), .A2(n63), .ZN(n763) );
  NAND2 U3453 ( .A1(n27421), .A2(n66), .ZN(n765) );
  NAND2 U3454 ( .A1(n27419), .A2(n69), .ZN(n767) );
  NAND2 U3455 ( .A1(n27421), .A2(n72), .ZN(n769) );
  NAND2 U3456 ( .A1(n27420), .A2(n75), .ZN(n771) );
  NAND2 U3457 ( .A1(n27421), .A2(n78), .ZN(n773) );
  NAND2 U3458 ( .A1(n27419), .A2(n81), .ZN(n775) );
  NAND2 U3459 ( .A1(n27419), .A2(n84), .ZN(n777) );
  NAND2 U3460 ( .A1(n27420), .A2(n87), .ZN(n779) );
  NAND2 U3461 ( .A1(n27421), .A2(n90), .ZN(n781) );
  NAND2 U3462 ( .A1(n27419), .A2(n93), .ZN(n783) );
  NAND2 U3463 ( .A1(n27420), .A2(n96), .ZN(n785) );
  NAND2 U3464 ( .A1(n27420), .A2(n99), .ZN(n787) );
  NAND2 U3465 ( .A1(n27420), .A2(n102), .ZN(n789) );
  NAND2 U3466 ( .A1(n27420), .A2(n105), .ZN(n791) );
  NAND2 U3467 ( .A1(n27420), .A2(n108), .ZN(n793) );
  NAND2 U3468 ( .A1(n27420), .A2(n111), .ZN(n795) );
  NAND2 U3469 ( .A1(n27420), .A2(n114), .ZN(n797) );
  NAND2 U3470 ( .A1(n27420), .A2(n117), .ZN(n799) );
  NAND2 U3471 ( .A1(n27420), .A2(n120), .ZN(n801) );
  NAND2 U3472 ( .A1(n27420), .A2(n123), .ZN(n803) );
  NAND2 U3473 ( .A1(n27420), .A2(n126), .ZN(n805) );
  NAND2 U3474 ( .A1(n27420), .A2(n129), .ZN(n807) );
  NAND2 U3475 ( .A1(n27421), .A2(n132), .ZN(n809) );
  NAND2 U3476 ( .A1(n27421), .A2(n135), .ZN(n811) );
  NAND2 U3477 ( .A1(n27421), .A2(n138), .ZN(n813) );
  NAND2 U3478 ( .A1(n27421), .A2(n141), .ZN(n815) );
  NAND2 U3479 ( .A1(n27421), .A2(n144), .ZN(n817) );
  NAND2 U3480 ( .A1(n27421), .A2(n147), .ZN(n819) );
  NAND2 U3481 ( .A1(n27421), .A2(n150), .ZN(n821) );
  NAND2 U3482 ( .A1(n27421), .A2(n153), .ZN(n823) );
  NAND2 U3483 ( .A1(n27421), .A2(n156), .ZN(n825) );
  NAND2 U3484 ( .A1(n27421), .A2(n159), .ZN(n827) );
  NAND2 U3485 ( .A1(n27421), .A2(n162), .ZN(n829) );
  NAND2 U3486 ( .A1(n27421), .A2(n165), .ZN(n831) );
  NAND2 U3487 ( .A1(n27421), .A2(n10), .ZN(n833) );
  NAND2 U3488 ( .A1(n27419), .A2(n11), .ZN(n835) );
  NAND2 U3489 ( .A1(n27420), .A2(n12), .ZN(n837) );
  NAND2 U3490 ( .A1(n27421), .A2(n24), .ZN(n839) );
  NAND2 U3491 ( .A1(n27419), .A2(n27), .ZN(n841) );
  NAND2 U3492 ( .A1(n27420), .A2(n30), .ZN(n843) );
  NAND2 U3493 ( .A1(n27421), .A2(n33), .ZN(n845) );
  NAND2 U3494 ( .A1(n27419), .A2(n36), .ZN(n847) );
  NAND2 U3495 ( .A1(n27420), .A2(n39), .ZN(n849) );
  NAND2 U3496 ( .A1(n27421), .A2(n168), .ZN(n851) );
  NAND2 U3497 ( .A1(n27419), .A2(n171), .ZN(n853) );
  NAND2 U3498 ( .A1(n27420), .A2(n174), .ZN(n855) );
  NAND2 U3499 ( .A1(n27416), .A2(n23), .ZN(n866) );
  NAND2 U3500 ( .A1(n27416), .A2(n5), .ZN(n869) );
  NAND2 U3501 ( .A1(n27416), .A2(n6), .ZN(n871) );
  NAND2 U3502 ( .A1(n27416), .A2(n7), .ZN(n873) );
  NAND2 U3503 ( .A1(n27416), .A2(n8), .ZN(n875) );
  NAND2 U3504 ( .A1(n27416), .A2(n9), .ZN(n877) );
  NAND2 U3505 ( .A1(n27416), .A2(n42), .ZN(n879) );
  NAND2 U3506 ( .A1(n27416), .A2(n45), .ZN(n881) );
  NAND2 U3507 ( .A1(n27416), .A2(n48), .ZN(n883) );
  NAND2 U3508 ( .A1(n27416), .A2(n51), .ZN(n885) );
  NAND2 U3509 ( .A1(n27416), .A2(n54), .ZN(n887) );
  NAND2 U3510 ( .A1(n27416), .A2(n57), .ZN(n889) );
  NAND2 U3511 ( .A1(n27417), .A2(n60), .ZN(n891) );
  NAND2 U3512 ( .A1(n27417), .A2(n63), .ZN(n893) );
  NAND2 U3513 ( .A1(n27418), .A2(n66), .ZN(n895) );
  NAND2 U3514 ( .A1(n27416), .A2(n69), .ZN(n897) );
  NAND2 U3515 ( .A1(n27418), .A2(n72), .ZN(n899) );
  NAND2 U3516 ( .A1(n27417), .A2(n75), .ZN(n901) );
  NAND2 U3517 ( .A1(n27418), .A2(n78), .ZN(n903) );
  NAND2 U3518 ( .A1(n27416), .A2(n81), .ZN(n905) );
  NAND2 U3519 ( .A1(n27416), .A2(n84), .ZN(n907) );
  NAND2 U3520 ( .A1(n27417), .A2(n87), .ZN(n909) );
  NAND2 U3521 ( .A1(n27418), .A2(n90), .ZN(n911) );
  NAND2 U3522 ( .A1(n27416), .A2(n93), .ZN(n913) );
  NAND2 U3523 ( .A1(n27417), .A2(n96), .ZN(n915) );
  NAND2 U3524 ( .A1(n27417), .A2(n99), .ZN(n917) );
  NAND2 U3525 ( .A1(n27417), .A2(n102), .ZN(n919) );
  NAND2 U3526 ( .A1(n27417), .A2(n105), .ZN(n921) );
  NAND2 U3527 ( .A1(n27417), .A2(n108), .ZN(n923) );
  NAND2 U3528 ( .A1(n27417), .A2(n111), .ZN(n925) );
  NAND2 U3529 ( .A1(n27417), .A2(n114), .ZN(n927) );
  NAND2 U3530 ( .A1(n27417), .A2(n117), .ZN(n929) );
  NAND2 U3531 ( .A1(n27417), .A2(n120), .ZN(n931) );
  NAND2 U3532 ( .A1(n27417), .A2(n123), .ZN(n933) );
  NAND2 U3533 ( .A1(n27417), .A2(n126), .ZN(n935) );
  NAND2 U3534 ( .A1(n27417), .A2(n129), .ZN(n937) );
  NAND2 U3535 ( .A1(n27418), .A2(n132), .ZN(n939) );
  NAND2 U3536 ( .A1(n27418), .A2(n135), .ZN(n941) );
  NAND2 U3537 ( .A1(n27418), .A2(n138), .ZN(n943) );
  NAND2 U3538 ( .A1(n27418), .A2(n141), .ZN(n945) );
  NAND2 U3539 ( .A1(n27418), .A2(n144), .ZN(n947) );
  NAND2 U3540 ( .A1(n27418), .A2(n147), .ZN(n949) );
  NAND2 U3541 ( .A1(n27418), .A2(n150), .ZN(n951) );
  NAND2 U3542 ( .A1(n27418), .A2(n153), .ZN(n953) );
  NAND2 U3543 ( .A1(n27418), .A2(n156), .ZN(n955) );
  NAND2 U3544 ( .A1(n27418), .A2(n159), .ZN(n957) );
  NAND2 U3545 ( .A1(n27418), .A2(n162), .ZN(n959) );
  NAND2 U3546 ( .A1(n27418), .A2(n165), .ZN(n961) );
  NAND2 U3547 ( .A1(n27418), .A2(n10), .ZN(n963) );
  NAND2 U3548 ( .A1(n27416), .A2(n11), .ZN(n965) );
  NAND2 U3549 ( .A1(n27417), .A2(n12), .ZN(n967) );
  NAND2 U3550 ( .A1(n27418), .A2(n24), .ZN(n969) );
  NAND2 U3551 ( .A1(n27416), .A2(n27), .ZN(n971) );
  NAND2 U3552 ( .A1(n27417), .A2(n30), .ZN(n973) );
  NAND2 U3553 ( .A1(n27418), .A2(n33), .ZN(n975) );
  NAND2 U3554 ( .A1(n27416), .A2(n36), .ZN(n977) );
  NAND2 U3555 ( .A1(n27417), .A2(n39), .ZN(n979) );
  NAND2 U3556 ( .A1(n27418), .A2(n168), .ZN(n981) );
  NAND2 U3557 ( .A1(n27416), .A2(n171), .ZN(n983) );
  NAND2 U3558 ( .A1(n27417), .A2(n174), .ZN(n985) );
  NAND2 U3559 ( .A1(n27413), .A2(n23), .ZN(n996) );
  NAND2 U3560 ( .A1(n27413), .A2(n5), .ZN(n999) );
  NAND2 U3561 ( .A1(n27413), .A2(n6), .ZN(n1001) );
  NAND2 U3562 ( .A1(n27413), .A2(n7), .ZN(n1003) );
  NAND2 U3563 ( .A1(n27413), .A2(n8), .ZN(n1005) );
  NAND2 U3564 ( .A1(n27413), .A2(n9), .ZN(n1007) );
  NAND2 U3565 ( .A1(n27413), .A2(n42), .ZN(n1009) );
  NAND2 U3566 ( .A1(n27413), .A2(n45), .ZN(n1011) );
  NAND2 U3567 ( .A1(n27413), .A2(n48), .ZN(n1013) );
  NAND2 U3568 ( .A1(n27413), .A2(n51), .ZN(n1015) );
  NAND2 U3569 ( .A1(n27413), .A2(n54), .ZN(n1017) );
  NAND2 U3570 ( .A1(n27413), .A2(n57), .ZN(n1019) );
  NAND2 U3571 ( .A1(n27414), .A2(n60), .ZN(n1021) );
  NAND2 U3572 ( .A1(n27414), .A2(n63), .ZN(n1023) );
  NAND2 U3573 ( .A1(n27415), .A2(n66), .ZN(n1025) );
  NAND2 U3574 ( .A1(n27413), .A2(n69), .ZN(n1027) );
  NAND2 U3575 ( .A1(n27415), .A2(n72), .ZN(n1029) );
  NAND2 U3576 ( .A1(n27414), .A2(n75), .ZN(n1031) );
  NAND2 U3577 ( .A1(n27415), .A2(n78), .ZN(n1033) );
  NAND2 U3578 ( .A1(n27413), .A2(n81), .ZN(n1035) );
  NAND2 U3579 ( .A1(n27413), .A2(n84), .ZN(n1037) );
  NAND2 U3580 ( .A1(n27414), .A2(n87), .ZN(n1039) );
  NAND2 U3581 ( .A1(n27415), .A2(n90), .ZN(n1041) );
  NAND2 U3582 ( .A1(n27413), .A2(n93), .ZN(n1043) );
  NAND2 U3583 ( .A1(n27414), .A2(n96), .ZN(n1045) );
  NAND2 U3584 ( .A1(n27414), .A2(n99), .ZN(n1047) );
  NAND2 U3585 ( .A1(n27414), .A2(n102), .ZN(n1049) );
  NAND2 U3586 ( .A1(n27414), .A2(n105), .ZN(n1051) );
  NAND2 U3587 ( .A1(n27414), .A2(n108), .ZN(n1053) );
  NAND2 U3588 ( .A1(n27414), .A2(n111), .ZN(n1055) );
  NAND2 U3589 ( .A1(n27414), .A2(n114), .ZN(n1057) );
  NAND2 U3590 ( .A1(n27414), .A2(n117), .ZN(n1059) );
  NAND2 U3591 ( .A1(n27414), .A2(n120), .ZN(n1061) );
  NAND2 U3592 ( .A1(n27414), .A2(n123), .ZN(n1063) );
  NAND2 U3593 ( .A1(n27414), .A2(n126), .ZN(n1065) );
  NAND2 U3594 ( .A1(n27414), .A2(n129), .ZN(n1067) );
  NAND2 U3595 ( .A1(n27415), .A2(n132), .ZN(n1069) );
  NAND2 U3596 ( .A1(n27415), .A2(n135), .ZN(n1071) );
  NAND2 U3597 ( .A1(n27415), .A2(n138), .ZN(n1073) );
  NAND2 U3598 ( .A1(n27415), .A2(n141), .ZN(n1075) );
  NAND2 U3599 ( .A1(n27415), .A2(n144), .ZN(n1077) );
  NAND2 U3600 ( .A1(n27415), .A2(n147), .ZN(n1079) );
  NAND2 U3601 ( .A1(n27415), .A2(n150), .ZN(n1081) );
  NAND2 U3602 ( .A1(n27415), .A2(n153), .ZN(n1083) );
  NAND2 U3603 ( .A1(n27415), .A2(n156), .ZN(n1085) );
  NAND2 U3604 ( .A1(n27415), .A2(n159), .ZN(n1087) );
  NAND2 U3605 ( .A1(n27415), .A2(n162), .ZN(n1089) );
  NAND2 U3606 ( .A1(n27415), .A2(n165), .ZN(n1091) );
  NAND2 U3607 ( .A1(n27415), .A2(n10), .ZN(n1093) );
  NAND2 U3608 ( .A1(n27413), .A2(n11), .ZN(n1095) );
  NAND2 U3609 ( .A1(n27414), .A2(n12), .ZN(n1097) );
  NAND2 U3610 ( .A1(n27415), .A2(n24), .ZN(n1099) );
  NAND2 U3611 ( .A1(n27413), .A2(n27), .ZN(n1101) );
  NAND2 U3612 ( .A1(n27414), .A2(n30), .ZN(n1103) );
  NAND2 U3613 ( .A1(n27415), .A2(n33), .ZN(n1105) );
  NAND2 U3614 ( .A1(n27413), .A2(n36), .ZN(n1107) );
  NAND2 U3615 ( .A1(n27414), .A2(n39), .ZN(n1109) );
  NAND2 U3616 ( .A1(n27415), .A2(n168), .ZN(n1111) );
  NAND2 U3617 ( .A1(n27413), .A2(n171), .ZN(n1113) );
  NAND2 U3618 ( .A1(n27414), .A2(n174), .ZN(n1115) );
  NAND2 U3619 ( .A1(n27410), .A2(n23), .ZN(n1126) );
  NAND2 U3620 ( .A1(n27410), .A2(n5), .ZN(n1129) );
  NAND2 U3621 ( .A1(n27410), .A2(n6), .ZN(n1131) );
  NAND2 U3622 ( .A1(n27410), .A2(n7), .ZN(n1133) );
  NAND2 U3623 ( .A1(n27410), .A2(n8), .ZN(n1135) );
  NAND2 U3624 ( .A1(n27410), .A2(n9), .ZN(n1137) );
  NAND2 U3625 ( .A1(n27410), .A2(n42), .ZN(n1139) );
  NAND2 U3626 ( .A1(n27410), .A2(n45), .ZN(n1141) );
  NAND2 U3627 ( .A1(n27410), .A2(n48), .ZN(n1143) );
  NAND2 U3628 ( .A1(n27410), .A2(n51), .ZN(n1145) );
  NAND2 U3629 ( .A1(n27410), .A2(n54), .ZN(n1147) );
  NAND2 U3630 ( .A1(n27410), .A2(n57), .ZN(n1149) );
  NAND2 U3631 ( .A1(n27411), .A2(n60), .ZN(n1151) );
  NAND2 U3632 ( .A1(n27411), .A2(n63), .ZN(n1153) );
  NAND2 U3633 ( .A1(n27411), .A2(n66), .ZN(n1155) );
  NAND2 U3634 ( .A1(n27411), .A2(n69), .ZN(n1157) );
  NAND2 U3635 ( .A1(n27411), .A2(n72), .ZN(n1159) );
  NAND2 U3636 ( .A1(n27411), .A2(n75), .ZN(n1161) );
  NAND2 U3637 ( .A1(n27411), .A2(n78), .ZN(n1163) );
  NAND2 U3638 ( .A1(n27411), .A2(n81), .ZN(n1165) );
  NAND2 U3639 ( .A1(n27411), .A2(n84), .ZN(n1167) );
  NAND2 U3640 ( .A1(n27411), .A2(n87), .ZN(n1169) );
  NAND2 U3641 ( .A1(n27411), .A2(n90), .ZN(n1171) );
  NAND2 U3642 ( .A1(n27411), .A2(n93), .ZN(n1173) );
  NAND2 U3643 ( .A1(n27412), .A2(n96), .ZN(n1175) );
  NAND2 U3644 ( .A1(n27412), .A2(n99), .ZN(n1177) );
  NAND2 U3645 ( .A1(n27412), .A2(n102), .ZN(n1179) );
  NAND2 U3646 ( .A1(n27412), .A2(n105), .ZN(n1181) );
  NAND2 U3647 ( .A1(n27412), .A2(n108), .ZN(n1183) );
  NAND2 U3648 ( .A1(n27412), .A2(n111), .ZN(n1185) );
  NAND2 U3649 ( .A1(n27412), .A2(n114), .ZN(n1187) );
  NAND2 U3650 ( .A1(n27412), .A2(n117), .ZN(n1189) );
  NAND2 U3651 ( .A1(n27412), .A2(n120), .ZN(n1191) );
  NAND2 U3652 ( .A1(n27412), .A2(n123), .ZN(n1193) );
  NAND2 U3653 ( .A1(n27412), .A2(n126), .ZN(n1195) );
  NAND2 U3654 ( .A1(n27412), .A2(n129), .ZN(n1197) );
  NAND2 U3655 ( .A1(n27411), .A2(n132), .ZN(n1199) );
  NAND2 U3656 ( .A1(n27412), .A2(n135), .ZN(n1201) );
  NAND2 U3657 ( .A1(n27410), .A2(n138), .ZN(n1203) );
  NAND2 U3658 ( .A1(n27411), .A2(n141), .ZN(n1205) );
  NAND2 U3659 ( .A1(n27412), .A2(n144), .ZN(n1207) );
  NAND2 U3660 ( .A1(n27410), .A2(n147), .ZN(n1209) );
  NAND2 U3661 ( .A1(n27411), .A2(n150), .ZN(n1211) );
  NAND2 U3662 ( .A1(n27412), .A2(n153), .ZN(n1213) );
  NAND2 U3663 ( .A1(n27410), .A2(n156), .ZN(n1215) );
  NAND2 U3664 ( .A1(n27411), .A2(n159), .ZN(n1217) );
  NAND2 U3665 ( .A1(n27412), .A2(n162), .ZN(n1219) );
  NAND2 U3666 ( .A1(n27410), .A2(n165), .ZN(n1221) );
  NAND2 U3667 ( .A1(n27412), .A2(n10), .ZN(n1223) );
  NAND2 U3668 ( .A1(n27410), .A2(n11), .ZN(n1225) );
  NAND2 U3669 ( .A1(n27410), .A2(n12), .ZN(n1227) );
  NAND2 U3670 ( .A1(n27411), .A2(n24), .ZN(n1229) );
  NAND2 U3671 ( .A1(n27412), .A2(n27), .ZN(n1231) );
  NAND2 U3672 ( .A1(n27411), .A2(n30), .ZN(n1233) );
  NAND2 U3673 ( .A1(n27410), .A2(n33), .ZN(n1235) );
  NAND2 U3674 ( .A1(n27411), .A2(n36), .ZN(n1237) );
  NAND2 U3675 ( .A1(n27412), .A2(n39), .ZN(n1239) );
  NAND2 U3676 ( .A1(n27412), .A2(n168), .ZN(n1241) );
  NAND2 U3677 ( .A1(n27410), .A2(n171), .ZN(n1243) );
  NAND2 U3678 ( .A1(n27411), .A2(n174), .ZN(n1245) );
  NAND2 U3679 ( .A1(n27407), .A2(n23), .ZN(n1256) );
  NAND2 U3680 ( .A1(n27407), .A2(n5), .ZN(n1259) );
  NAND2 U3681 ( .A1(n27407), .A2(n6), .ZN(n1261) );
  NAND2 U3682 ( .A1(n27407), .A2(n7), .ZN(n1263) );
  NAND2 U3683 ( .A1(n27407), .A2(n8), .ZN(n1265) );
  NAND2 U3684 ( .A1(n27407), .A2(n9), .ZN(n1267) );
  NAND2 U3685 ( .A1(n27407), .A2(n42), .ZN(n1269) );
  NAND2 U3686 ( .A1(n27407), .A2(n45), .ZN(n1271) );
  NAND2 U3687 ( .A1(n27407), .A2(n48), .ZN(n1273) );
  NAND2 U3688 ( .A1(n27407), .A2(n51), .ZN(n1275) );
  NAND2 U3689 ( .A1(n27407), .A2(n54), .ZN(n1277) );
  NAND2 U3690 ( .A1(n27407), .A2(n57), .ZN(n1279) );
  NAND2 U3691 ( .A1(n27408), .A2(n60), .ZN(n1281) );
  NAND2 U3692 ( .A1(n27408), .A2(n63), .ZN(n1283) );
  NAND2 U3693 ( .A1(n27408), .A2(n66), .ZN(n1285) );
  NAND2 U3694 ( .A1(n27408), .A2(n69), .ZN(n1287) );
  NAND2 U3695 ( .A1(n27408), .A2(n72), .ZN(n1289) );
  NAND2 U3696 ( .A1(n27408), .A2(n75), .ZN(n1291) );
  NAND2 U3697 ( .A1(n27408), .A2(n78), .ZN(n1293) );
  NAND2 U3698 ( .A1(n27408), .A2(n81), .ZN(n1295) );
  NAND2 U3699 ( .A1(n27408), .A2(n84), .ZN(n1297) );
  NAND2 U3700 ( .A1(n27408), .A2(n87), .ZN(n1299) );
  NAND2 U3701 ( .A1(n27408), .A2(n90), .ZN(n1301) );
  NAND2 U3702 ( .A1(n27408), .A2(n93), .ZN(n1303) );
  NAND2 U3703 ( .A1(n27409), .A2(n96), .ZN(n1305) );
  NAND2 U3704 ( .A1(n27409), .A2(n99), .ZN(n1307) );
  NAND2 U3705 ( .A1(n27409), .A2(n102), .ZN(n1309) );
  NAND2 U3706 ( .A1(n27409), .A2(n105), .ZN(n1311) );
  NAND2 U3707 ( .A1(n27409), .A2(n108), .ZN(n1313) );
  NAND2 U3708 ( .A1(n27409), .A2(n111), .ZN(n1315) );
  NAND2 U3709 ( .A1(n27409), .A2(n114), .ZN(n1317) );
  NAND2 U3710 ( .A1(n27409), .A2(n117), .ZN(n1319) );
  NAND2 U3711 ( .A1(n27409), .A2(n120), .ZN(n1321) );
  NAND2 U3712 ( .A1(n27409), .A2(n123), .ZN(n1323) );
  NAND2 U3713 ( .A1(n27409), .A2(n126), .ZN(n1325) );
  NAND2 U3714 ( .A1(n27409), .A2(n129), .ZN(n1327) );
  NAND2 U3715 ( .A1(n27408), .A2(n132), .ZN(n1329) );
  NAND2 U3716 ( .A1(n27409), .A2(n135), .ZN(n1331) );
  NAND2 U3717 ( .A1(n27407), .A2(n138), .ZN(n1333) );
  NAND2 U3718 ( .A1(n27408), .A2(n141), .ZN(n1335) );
  NAND2 U3719 ( .A1(n27409), .A2(n144), .ZN(n1337) );
  NAND2 U3720 ( .A1(n27407), .A2(n147), .ZN(n1339) );
  NAND2 U3721 ( .A1(n27408), .A2(n150), .ZN(n1341) );
  NAND2 U3722 ( .A1(n27409), .A2(n153), .ZN(n1343) );
  NAND2 U3723 ( .A1(n27407), .A2(n156), .ZN(n1345) );
  NAND2 U3724 ( .A1(n27408), .A2(n159), .ZN(n1347) );
  NAND2 U3725 ( .A1(n27409), .A2(n162), .ZN(n1349) );
  NAND2 U3726 ( .A1(n27407), .A2(n165), .ZN(n1351) );
  NAND2 U3727 ( .A1(n27409), .A2(n10), .ZN(n1353) );
  NAND2 U3728 ( .A1(n27407), .A2(n11), .ZN(n1355) );
  NAND2 U3729 ( .A1(n27407), .A2(n12), .ZN(n1357) );
  NAND2 U3730 ( .A1(n27408), .A2(n24), .ZN(n1359) );
  NAND2 U3731 ( .A1(n27409), .A2(n27), .ZN(n1361) );
  NAND2 U3732 ( .A1(n27408), .A2(n30), .ZN(n1363) );
  NAND2 U3733 ( .A1(n27407), .A2(n33), .ZN(n1365) );
  NAND2 U3734 ( .A1(n27408), .A2(n36), .ZN(n1367) );
  NAND2 U3735 ( .A1(n27409), .A2(n39), .ZN(n1369) );
  NAND2 U3736 ( .A1(n27409), .A2(n168), .ZN(n1371) );
  NAND2 U3737 ( .A1(n27407), .A2(n171), .ZN(n1373) );
  NAND2 U3738 ( .A1(n27408), .A2(n174), .ZN(n1375) );
  NAND2 U3739 ( .A1(n27404), .A2(n23), .ZN(n1385) );
  NAND2 U3740 ( .A1(n27404), .A2(n5), .ZN(n1388) );
  NAND2 U3741 ( .A1(n27404), .A2(n6), .ZN(n1390) );
  NAND2 U3742 ( .A1(n27404), .A2(n7), .ZN(n1392) );
  NAND2 U3743 ( .A1(n27404), .A2(n8), .ZN(n1394) );
  NAND2 U3744 ( .A1(n27404), .A2(n9), .ZN(n1396) );
  NAND2 U3745 ( .A1(n27404), .A2(n42), .ZN(n1398) );
  NAND2 U3746 ( .A1(n27404), .A2(n45), .ZN(n1400) );
  NAND2 U3747 ( .A1(n27404), .A2(n48), .ZN(n1402) );
  NAND2 U3748 ( .A1(n27404), .A2(n51), .ZN(n1404) );
  NAND2 U3749 ( .A1(n27404), .A2(n54), .ZN(n1406) );
  NAND2 U3750 ( .A1(n27404), .A2(n57), .ZN(n1408) );
  NAND2 U3751 ( .A1(n27405), .A2(n60), .ZN(n1410) );
  NAND2 U3752 ( .A1(n27405), .A2(n63), .ZN(n1412) );
  NAND2 U3753 ( .A1(n27405), .A2(n66), .ZN(n1414) );
  NAND2 U3754 ( .A1(n27405), .A2(n69), .ZN(n1416) );
  NAND2 U3755 ( .A1(n27405), .A2(n72), .ZN(n1418) );
  NAND2 U3756 ( .A1(n27405), .A2(n75), .ZN(n1420) );
  NAND2 U3757 ( .A1(n27405), .A2(n78), .ZN(n1422) );
  NAND2 U3758 ( .A1(n27405), .A2(n81), .ZN(n1424) );
  NAND2 U3759 ( .A1(n27405), .A2(n84), .ZN(n1426) );
  NAND2 U3760 ( .A1(n27405), .A2(n87), .ZN(n1428) );
  NAND2 U3761 ( .A1(n27405), .A2(n90), .ZN(n1430) );
  NAND2 U3762 ( .A1(n27405), .A2(n93), .ZN(n1432) );
  NAND2 U3763 ( .A1(n27406), .A2(n96), .ZN(n1434) );
  NAND2 U3764 ( .A1(n27406), .A2(n99), .ZN(n1436) );
  NAND2 U3765 ( .A1(n27406), .A2(n102), .ZN(n1438) );
  NAND2 U3766 ( .A1(n27406), .A2(n105), .ZN(n1440) );
  NAND2 U3767 ( .A1(n27406), .A2(n108), .ZN(n1442) );
  NAND2 U3768 ( .A1(n27406), .A2(n111), .ZN(n1444) );
  NAND2 U3769 ( .A1(n27406), .A2(n114), .ZN(n1446) );
  NAND2 U3770 ( .A1(n27406), .A2(n117), .ZN(n1448) );
  NAND2 U3771 ( .A1(n27406), .A2(n120), .ZN(n1450) );
  NAND2 U3772 ( .A1(n27406), .A2(n123), .ZN(n1452) );
  NAND2 U3773 ( .A1(n27406), .A2(n126), .ZN(n1454) );
  NAND2 U3774 ( .A1(n27406), .A2(n129), .ZN(n1456) );
  NAND2 U3775 ( .A1(n27405), .A2(n132), .ZN(n1458) );
  NAND2 U3776 ( .A1(n27406), .A2(n135), .ZN(n1460) );
  NAND2 U3777 ( .A1(n27404), .A2(n138), .ZN(n1462) );
  NAND2 U3778 ( .A1(n27405), .A2(n141), .ZN(n1464) );
  NAND2 U3779 ( .A1(n27406), .A2(n144), .ZN(n1466) );
  NAND2 U3780 ( .A1(n27404), .A2(n147), .ZN(n1468) );
  NAND2 U3781 ( .A1(n27405), .A2(n150), .ZN(n1470) );
  NAND2 U3782 ( .A1(n27406), .A2(n153), .ZN(n1472) );
  NAND2 U3783 ( .A1(n27404), .A2(n156), .ZN(n1474) );
  NAND2 U3784 ( .A1(n27405), .A2(n159), .ZN(n1476) );
  NAND2 U3785 ( .A1(n27406), .A2(n162), .ZN(n1478) );
  NAND2 U3786 ( .A1(n27404), .A2(n165), .ZN(n1480) );
  NAND2 U3787 ( .A1(n27406), .A2(n10), .ZN(n1482) );
  NAND2 U3788 ( .A1(n27404), .A2(n11), .ZN(n1484) );
  NAND2 U3789 ( .A1(n27404), .A2(n12), .ZN(n1486) );
  NAND2 U3790 ( .A1(n27405), .A2(n24), .ZN(n1488) );
  NAND2 U3791 ( .A1(n27406), .A2(n27), .ZN(n1490) );
  NAND2 U3792 ( .A1(n27405), .A2(n30), .ZN(n1492) );
  NAND2 U3793 ( .A1(n27404), .A2(n33), .ZN(n1494) );
  NAND2 U3794 ( .A1(n27405), .A2(n36), .ZN(n1496) );
  NAND2 U3795 ( .A1(n27406), .A2(n39), .ZN(n1498) );
  NAND2 U3796 ( .A1(n27406), .A2(n168), .ZN(n1500) );
  NAND2 U3797 ( .A1(n27404), .A2(n171), .ZN(n1502) );
  NAND2 U3798 ( .A1(n27405), .A2(n174), .ZN(n1504) );
  NAND2 U3799 ( .A1(n27401), .A2(n23), .ZN(n1514) );
  NAND2 U3800 ( .A1(n27401), .A2(n5), .ZN(n1517) );
  NAND2 U3801 ( .A1(n27401), .A2(n6), .ZN(n1519) );
  NAND2 U3802 ( .A1(n27401), .A2(n7), .ZN(n1521) );
  NAND2 U3803 ( .A1(n27401), .A2(n8), .ZN(n1523) );
  NAND2 U3804 ( .A1(n27401), .A2(n9), .ZN(n1525) );
  NAND2 U3805 ( .A1(n27401), .A2(n42), .ZN(n1527) );
  NAND2 U3806 ( .A1(n27401), .A2(n45), .ZN(n1529) );
  NAND2 U3807 ( .A1(n27401), .A2(n48), .ZN(n1531) );
  NAND2 U3808 ( .A1(n27401), .A2(n51), .ZN(n1533) );
  NAND2 U3809 ( .A1(n27401), .A2(n54), .ZN(n1535) );
  NAND2 U3810 ( .A1(n27401), .A2(n57), .ZN(n1537) );
  NAND2 U3811 ( .A1(n27402), .A2(n60), .ZN(n1539) );
  NAND2 U3812 ( .A1(n27402), .A2(n63), .ZN(n1541) );
  NAND2 U3813 ( .A1(n27402), .A2(n66), .ZN(n1543) );
  NAND2 U3814 ( .A1(n27402), .A2(n69), .ZN(n1545) );
  NAND2 U3815 ( .A1(n27402), .A2(n72), .ZN(n1547) );
  NAND2 U3816 ( .A1(n27402), .A2(n75), .ZN(n1549) );
  NAND2 U3817 ( .A1(n27402), .A2(n78), .ZN(n1551) );
  NAND2 U3818 ( .A1(n27402), .A2(n81), .ZN(n1553) );
  NAND2 U3819 ( .A1(n27402), .A2(n84), .ZN(n1555) );
  NAND2 U3820 ( .A1(n27402), .A2(n87), .ZN(n1557) );
  NAND2 U3821 ( .A1(n27402), .A2(n90), .ZN(n1559) );
  NAND2 U3822 ( .A1(n27402), .A2(n93), .ZN(n1561) );
  NAND2 U3823 ( .A1(n27403), .A2(n96), .ZN(n1563) );
  NAND2 U3824 ( .A1(n27403), .A2(n99), .ZN(n1565) );
  NAND2 U3825 ( .A1(n27403), .A2(n102), .ZN(n1567) );
  NAND2 U3826 ( .A1(n27403), .A2(n105), .ZN(n1569) );
  NAND2 U3827 ( .A1(n27403), .A2(n108), .ZN(n1571) );
  NAND2 U3828 ( .A1(n27403), .A2(n111), .ZN(n1573) );
  NAND2 U3829 ( .A1(n27403), .A2(n114), .ZN(n1575) );
  NAND2 U3830 ( .A1(n27403), .A2(n117), .ZN(n1577) );
  NAND2 U3831 ( .A1(n27403), .A2(n120), .ZN(n1579) );
  NAND2 U3832 ( .A1(n27403), .A2(n123), .ZN(n1581) );
  NAND2 U3833 ( .A1(n27403), .A2(n126), .ZN(n1583) );
  NAND2 U3834 ( .A1(n27403), .A2(n129), .ZN(n1585) );
  NAND2 U3835 ( .A1(n27402), .A2(n132), .ZN(n1587) );
  NAND2 U3836 ( .A1(n27403), .A2(n135), .ZN(n1589) );
  NAND2 U3837 ( .A1(n27401), .A2(n138), .ZN(n1591) );
  NAND2 U3838 ( .A1(n27402), .A2(n141), .ZN(n1593) );
  NAND2 U3839 ( .A1(n27403), .A2(n144), .ZN(n1595) );
  NAND2 U3840 ( .A1(n27401), .A2(n147), .ZN(n1597) );
  NAND2 U3841 ( .A1(n27402), .A2(n150), .ZN(n1599) );
  NAND2 U3842 ( .A1(n27403), .A2(n153), .ZN(n1601) );
  NAND2 U3843 ( .A1(n27401), .A2(n156), .ZN(n1603) );
  NAND2 U3844 ( .A1(n27402), .A2(n159), .ZN(n1605) );
  NAND2 U3845 ( .A1(n27403), .A2(n162), .ZN(n1607) );
  NAND2 U3846 ( .A1(n27401), .A2(n165), .ZN(n1609) );
  NAND2 U3847 ( .A1(n27403), .A2(n10), .ZN(n1611) );
  NAND2 U3848 ( .A1(n27401), .A2(n11), .ZN(n1613) );
  NAND2 U3849 ( .A1(n27401), .A2(n12), .ZN(n1615) );
  NAND2 U3850 ( .A1(n27402), .A2(n24), .ZN(n1617) );
  NAND2 U3851 ( .A1(n27403), .A2(n27), .ZN(n1619) );
  NAND2 U3852 ( .A1(n27402), .A2(n30), .ZN(n1621) );
  NAND2 U3853 ( .A1(n27401), .A2(n33), .ZN(n1623) );
  NAND2 U3854 ( .A1(n27402), .A2(n36), .ZN(n1625) );
  NAND2 U3855 ( .A1(n27403), .A2(n39), .ZN(n1627) );
  NAND2 U3856 ( .A1(n27403), .A2(n168), .ZN(n1629) );
  NAND2 U3857 ( .A1(n27401), .A2(n171), .ZN(n1631) );
  NAND2 U3858 ( .A1(n27402), .A2(n174), .ZN(n1633) );
  NAND2 U3859 ( .A1(n27398), .A2(n23), .ZN(n1643) );
  NAND2 U3860 ( .A1(n27398), .A2(n5), .ZN(n1646) );
  NAND2 U3861 ( .A1(n27398), .A2(n6), .ZN(n1648) );
  NAND2 U3862 ( .A1(n27398), .A2(n7), .ZN(n1650) );
  NAND2 U3863 ( .A1(n27398), .A2(n8), .ZN(n1652) );
  NAND2 U3864 ( .A1(n27398), .A2(n9), .ZN(n1654) );
  NAND2 U3865 ( .A1(n27398), .A2(n42), .ZN(n1656) );
  NAND2 U3866 ( .A1(n27398), .A2(n45), .ZN(n1658) );
  NAND2 U3867 ( .A1(n27398), .A2(n48), .ZN(n1660) );
  NAND2 U3868 ( .A1(n27398), .A2(n51), .ZN(n1662) );
  NAND2 U3869 ( .A1(n27398), .A2(n54), .ZN(n1664) );
  NAND2 U3870 ( .A1(n27398), .A2(n57), .ZN(n1666) );
  NAND2 U3871 ( .A1(n27399), .A2(n60), .ZN(n1668) );
  NAND2 U3872 ( .A1(n27399), .A2(n63), .ZN(n1670) );
  NAND2 U3873 ( .A1(n27399), .A2(n66), .ZN(n1672) );
  NAND2 U3874 ( .A1(n27399), .A2(n69), .ZN(n1674) );
  NAND2 U3875 ( .A1(n27399), .A2(n72), .ZN(n1676) );
  NAND2 U3876 ( .A1(n27399), .A2(n75), .ZN(n1678) );
  NAND2 U3877 ( .A1(n27399), .A2(n78), .ZN(n1680) );
  NAND2 U3878 ( .A1(n27399), .A2(n81), .ZN(n1682) );
  NAND2 U3879 ( .A1(n27399), .A2(n84), .ZN(n1684) );
  NAND2 U3880 ( .A1(n27399), .A2(n87), .ZN(n1686) );
  NAND2 U3881 ( .A1(n27399), .A2(n90), .ZN(n1688) );
  NAND2 U3882 ( .A1(n27399), .A2(n93), .ZN(n1690) );
  NAND2 U3883 ( .A1(n27400), .A2(n96), .ZN(n1692) );
  NAND2 U3884 ( .A1(n27400), .A2(n99), .ZN(n1694) );
  NAND2 U3885 ( .A1(n27400), .A2(n102), .ZN(n1696) );
  NAND2 U3886 ( .A1(n27400), .A2(n105), .ZN(n1698) );
  NAND2 U3887 ( .A1(n27400), .A2(n108), .ZN(n1700) );
  NAND2 U3888 ( .A1(n27400), .A2(n111), .ZN(n1702) );
  NAND2 U3889 ( .A1(n27400), .A2(n114), .ZN(n1704) );
  NAND2 U3890 ( .A1(n27400), .A2(n117), .ZN(n1706) );
  NAND2 U3891 ( .A1(n27400), .A2(n120), .ZN(n1708) );
  NAND2 U3892 ( .A1(n27400), .A2(n123), .ZN(n1710) );
  NAND2 U3893 ( .A1(n27400), .A2(n126), .ZN(n1712) );
  NAND2 U3894 ( .A1(n27400), .A2(n129), .ZN(n1714) );
  NAND2 U3895 ( .A1(n27399), .A2(n132), .ZN(n1716) );
  NAND2 U3896 ( .A1(n27400), .A2(n135), .ZN(n1718) );
  NAND2 U3897 ( .A1(n27398), .A2(n138), .ZN(n1720) );
  NAND2 U3898 ( .A1(n27399), .A2(n141), .ZN(n1722) );
  NAND2 U3899 ( .A1(n27400), .A2(n144), .ZN(n1724) );
  NAND2 U3900 ( .A1(n27398), .A2(n147), .ZN(n1726) );
  NAND2 U3901 ( .A1(n27399), .A2(n150), .ZN(n1728) );
  NAND2 U3902 ( .A1(n27400), .A2(n153), .ZN(n1730) );
  NAND2 U3903 ( .A1(n27398), .A2(n156), .ZN(n1732) );
  NAND2 U3904 ( .A1(n27399), .A2(n159), .ZN(n1734) );
  NAND2 U3905 ( .A1(n27400), .A2(n162), .ZN(n1736) );
  NAND2 U3906 ( .A1(n27398), .A2(n165), .ZN(n1738) );
  NAND2 U3907 ( .A1(n27400), .A2(n10), .ZN(n1740) );
  NAND2 U3908 ( .A1(n27398), .A2(n11), .ZN(n1742) );
  NAND2 U3909 ( .A1(n27398), .A2(n12), .ZN(n1744) );
  NAND2 U3910 ( .A1(n27399), .A2(n24), .ZN(n1746) );
  NAND2 U3911 ( .A1(n27400), .A2(n27), .ZN(n1748) );
  NAND2 U3912 ( .A1(n27399), .A2(n30), .ZN(n1750) );
  NAND2 U3913 ( .A1(n27398), .A2(n33), .ZN(n1752) );
  NAND2 U3914 ( .A1(n27399), .A2(n36), .ZN(n1754) );
  NAND2 U3915 ( .A1(n27400), .A2(n39), .ZN(n1756) );
  NAND2 U3916 ( .A1(n27400), .A2(n168), .ZN(n1758) );
  NAND2 U3917 ( .A1(n27398), .A2(n171), .ZN(n1760) );
  NAND2 U3918 ( .A1(n27399), .A2(n174), .ZN(n1762) );
  NAND2 U3919 ( .A1(n27395), .A2(n23), .ZN(n1772) );
  NAND2 U3920 ( .A1(n27395), .A2(n5), .ZN(n1775) );
  NAND2 U3921 ( .A1(n27395), .A2(n6), .ZN(n1777) );
  NAND2 U3922 ( .A1(n27395), .A2(n7), .ZN(n1779) );
  NAND2 U3923 ( .A1(n27395), .A2(n8), .ZN(n1781) );
  NAND2 U3924 ( .A1(n27395), .A2(n9), .ZN(n1783) );
  NAND2 U3925 ( .A1(n27395), .A2(n42), .ZN(n1785) );
  NAND2 U3926 ( .A1(n27395), .A2(n45), .ZN(n1787) );
  NAND2 U3927 ( .A1(n27395), .A2(n48), .ZN(n1789) );
  NAND2 U3928 ( .A1(n27395), .A2(n51), .ZN(n1791) );
  NAND2 U3929 ( .A1(n27395), .A2(n54), .ZN(n1793) );
  NAND2 U3930 ( .A1(n27395), .A2(n57), .ZN(n1795) );
  NAND2 U3931 ( .A1(n27396), .A2(n60), .ZN(n1797) );
  NAND2 U3932 ( .A1(n27396), .A2(n63), .ZN(n1799) );
  NAND2 U3933 ( .A1(n27396), .A2(n66), .ZN(n1801) );
  NAND2 U3934 ( .A1(n27396), .A2(n69), .ZN(n1803) );
  NAND2 U3935 ( .A1(n27396), .A2(n72), .ZN(n1805) );
  NAND2 U3936 ( .A1(n27396), .A2(n75), .ZN(n1807) );
  NAND2 U3937 ( .A1(n27396), .A2(n78), .ZN(n1809) );
  NAND2 U3938 ( .A1(n27396), .A2(n81), .ZN(n1811) );
  NAND2 U3939 ( .A1(n27396), .A2(n84), .ZN(n1813) );
  NAND2 U3940 ( .A1(n27396), .A2(n87), .ZN(n1815) );
  NAND2 U3941 ( .A1(n27396), .A2(n90), .ZN(n1817) );
  NAND2 U3942 ( .A1(n27396), .A2(n93), .ZN(n1819) );
  NAND2 U3943 ( .A1(n27397), .A2(n96), .ZN(n1821) );
  NAND2 U3944 ( .A1(n27397), .A2(n99), .ZN(n1823) );
  NAND2 U3945 ( .A1(n27397), .A2(n102), .ZN(n1825) );
  NAND2 U3946 ( .A1(n27397), .A2(n105), .ZN(n1827) );
  NAND2 U3947 ( .A1(n27397), .A2(n108), .ZN(n1829) );
  NAND2 U3948 ( .A1(n27397), .A2(n111), .ZN(n1831) );
  NAND2 U3949 ( .A1(n27397), .A2(n114), .ZN(n1833) );
  NAND2 U3950 ( .A1(n27397), .A2(n117), .ZN(n1835) );
  NAND2 U3951 ( .A1(n27397), .A2(n120), .ZN(n1837) );
  NAND2 U3952 ( .A1(n27397), .A2(n123), .ZN(n1839) );
  NAND2 U3953 ( .A1(n27397), .A2(n126), .ZN(n1841) );
  NAND2 U3954 ( .A1(n27397), .A2(n129), .ZN(n1843) );
  NAND2 U3955 ( .A1(n27396), .A2(n132), .ZN(n1845) );
  NAND2 U3956 ( .A1(n27397), .A2(n135), .ZN(n1847) );
  NAND2 U3957 ( .A1(n27395), .A2(n138), .ZN(n1849) );
  NAND2 U3958 ( .A1(n27396), .A2(n141), .ZN(n1851) );
  NAND2 U3959 ( .A1(n27397), .A2(n144), .ZN(n1853) );
  NAND2 U3960 ( .A1(n27395), .A2(n147), .ZN(n1855) );
  NAND2 U3961 ( .A1(n27396), .A2(n150), .ZN(n1857) );
  NAND2 U3962 ( .A1(n27397), .A2(n153), .ZN(n1859) );
  NAND2 U3963 ( .A1(n27395), .A2(n156), .ZN(n1861) );
  NAND2 U3964 ( .A1(n27396), .A2(n159), .ZN(n1863) );
  NAND2 U3965 ( .A1(n27397), .A2(n162), .ZN(n1865) );
  NAND2 U3966 ( .A1(n27395), .A2(n165), .ZN(n1867) );
  NAND2 U3967 ( .A1(n27397), .A2(n10), .ZN(n1869) );
  NAND2 U3968 ( .A1(n27395), .A2(n11), .ZN(n1871) );
  NAND2 U3969 ( .A1(n27395), .A2(n12), .ZN(n1873) );
  NAND2 U3970 ( .A1(n27396), .A2(n24), .ZN(n1875) );
  NAND2 U3971 ( .A1(n27397), .A2(n27), .ZN(n1877) );
  NAND2 U3972 ( .A1(n27396), .A2(n30), .ZN(n1879) );
  NAND2 U3973 ( .A1(n27395), .A2(n33), .ZN(n1881) );
  NAND2 U3974 ( .A1(n27396), .A2(n36), .ZN(n1883) );
  NAND2 U3975 ( .A1(n27397), .A2(n39), .ZN(n1885) );
  NAND2 U3976 ( .A1(n27397), .A2(n168), .ZN(n1887) );
  NAND2 U3977 ( .A1(n27395), .A2(n171), .ZN(n1889) );
  NAND2 U3978 ( .A1(n27396), .A2(n174), .ZN(n1891) );
  NAND2 U3979 ( .A1(n27392), .A2(n23), .ZN(n1901) );
  NAND2 U3980 ( .A1(n27392), .A2(n5), .ZN(n1904) );
  NAND2 U3981 ( .A1(n27392), .A2(n6), .ZN(n1906) );
  NAND2 U3982 ( .A1(n27392), .A2(n7), .ZN(n1908) );
  NAND2 U3983 ( .A1(n27392), .A2(n8), .ZN(n1910) );
  NAND2 U3984 ( .A1(n27392), .A2(n9), .ZN(n1912) );
  NAND2 U3985 ( .A1(n27392), .A2(n42), .ZN(n1914) );
  NAND2 U3986 ( .A1(n27392), .A2(n45), .ZN(n1916) );
  NAND2 U3987 ( .A1(n27392), .A2(n48), .ZN(n1918) );
  NAND2 U3988 ( .A1(n27392), .A2(n51), .ZN(n1920) );
  NAND2 U3989 ( .A1(n27392), .A2(n54), .ZN(n1922) );
  NAND2 U3990 ( .A1(n27392), .A2(n57), .ZN(n1924) );
  NAND2 U3991 ( .A1(n27393), .A2(n60), .ZN(n1926) );
  NAND2 U3992 ( .A1(n27393), .A2(n63), .ZN(n1928) );
  NAND2 U3993 ( .A1(n27393), .A2(n66), .ZN(n1930) );
  NAND2 U3994 ( .A1(n27393), .A2(n69), .ZN(n1932) );
  NAND2 U3995 ( .A1(n27393), .A2(n72), .ZN(n1934) );
  NAND2 U3996 ( .A1(n27393), .A2(n75), .ZN(n1936) );
  NAND2 U3997 ( .A1(n27393), .A2(n78), .ZN(n1938) );
  NAND2 U3998 ( .A1(n27393), .A2(n81), .ZN(n1940) );
  NAND2 U3999 ( .A1(n27393), .A2(n84), .ZN(n1942) );
  NAND2 U4000 ( .A1(n27393), .A2(n87), .ZN(n1944) );
  NAND2 U4001 ( .A1(n27393), .A2(n90), .ZN(n1946) );
  NAND2 U4002 ( .A1(n27393), .A2(n93), .ZN(n1948) );
  NAND2 U4003 ( .A1(n27394), .A2(n96), .ZN(n1950) );
  NAND2 U4004 ( .A1(n27394), .A2(n99), .ZN(n1952) );
  NAND2 U4005 ( .A1(n27394), .A2(n102), .ZN(n1954) );
  NAND2 U4006 ( .A1(n27394), .A2(n105), .ZN(n1956) );
  NAND2 U4007 ( .A1(n27394), .A2(n108), .ZN(n1958) );
  NAND2 U4008 ( .A1(n27394), .A2(n111), .ZN(n1960) );
  NAND2 U4009 ( .A1(n27394), .A2(n114), .ZN(n1962) );
  NAND2 U4010 ( .A1(n27394), .A2(n117), .ZN(n1964) );
  NAND2 U4011 ( .A1(n27394), .A2(n120), .ZN(n1966) );
  NAND2 U4012 ( .A1(n27394), .A2(n123), .ZN(n1968) );
  NAND2 U4013 ( .A1(n27394), .A2(n126), .ZN(n1970) );
  NAND2 U4014 ( .A1(n27394), .A2(n129), .ZN(n1972) );
  NAND2 U4015 ( .A1(n27393), .A2(n132), .ZN(n1974) );
  NAND2 U4016 ( .A1(n27394), .A2(n135), .ZN(n1976) );
  NAND2 U4017 ( .A1(n27392), .A2(n138), .ZN(n1978) );
  NAND2 U4018 ( .A1(n27393), .A2(n141), .ZN(n1980) );
  NAND2 U4019 ( .A1(n27394), .A2(n144), .ZN(n1982) );
  NAND2 U4020 ( .A1(n27392), .A2(n147), .ZN(n1984) );
  NAND2 U4021 ( .A1(n27393), .A2(n150), .ZN(n1986) );
  NAND2 U4022 ( .A1(n27394), .A2(n153), .ZN(n1988) );
  NAND2 U4023 ( .A1(n27392), .A2(n156), .ZN(n1990) );
  NAND2 U4024 ( .A1(n27393), .A2(n159), .ZN(n1992) );
  NAND2 U4025 ( .A1(n27394), .A2(n162), .ZN(n1994) );
  NAND2 U4026 ( .A1(n27392), .A2(n165), .ZN(n1996) );
  NAND2 U4027 ( .A1(n27394), .A2(n10), .ZN(n1998) );
  NAND2 U4028 ( .A1(n27392), .A2(n11), .ZN(n2000) );
  NAND2 U4029 ( .A1(n27392), .A2(n12), .ZN(n2002) );
  NAND2 U4030 ( .A1(n27393), .A2(n24), .ZN(n2004) );
  NAND2 U4031 ( .A1(n27394), .A2(n27), .ZN(n2006) );
  NAND2 U4032 ( .A1(n27393), .A2(n30), .ZN(n2008) );
  NAND2 U4033 ( .A1(n27392), .A2(n33), .ZN(n2010) );
  NAND2 U4034 ( .A1(n27393), .A2(n36), .ZN(n2012) );
  NAND2 U4035 ( .A1(n27394), .A2(n39), .ZN(n2014) );
  NAND2 U4036 ( .A1(n27394), .A2(n168), .ZN(n2016) );
  NAND2 U4037 ( .A1(n27392), .A2(n171), .ZN(n2018) );
  NAND2 U4038 ( .A1(n27393), .A2(n174), .ZN(n2020) );
  NAND2 U4039 ( .A1(n27389), .A2(n23), .ZN(n2030) );
  NAND2 U4040 ( .A1(n27389), .A2(n5), .ZN(n2033) );
  NAND2 U4041 ( .A1(n27389), .A2(n6), .ZN(n2035) );
  NAND2 U4042 ( .A1(n27389), .A2(n7), .ZN(n2037) );
  NAND2 U4043 ( .A1(n27389), .A2(n8), .ZN(n2039) );
  NAND2 U4044 ( .A1(n27389), .A2(n9), .ZN(n2041) );
  NAND2 U4045 ( .A1(n27389), .A2(n42), .ZN(n2043) );
  NAND2 U4046 ( .A1(n27389), .A2(n45), .ZN(n2045) );
  NAND2 U4047 ( .A1(n27389), .A2(n48), .ZN(n2047) );
  NAND2 U4048 ( .A1(n27389), .A2(n51), .ZN(n2049) );
  NAND2 U4049 ( .A1(n27389), .A2(n54), .ZN(n2051) );
  NAND2 U4050 ( .A1(n27389), .A2(n57), .ZN(n2053) );
  NAND2 U4051 ( .A1(n27390), .A2(n60), .ZN(n2055) );
  NAND2 U4052 ( .A1(n27390), .A2(n63), .ZN(n2057) );
  NAND2 U4053 ( .A1(n27390), .A2(n66), .ZN(n2059) );
  NAND2 U4054 ( .A1(n27390), .A2(n69), .ZN(n2061) );
  NAND2 U4055 ( .A1(n27390), .A2(n72), .ZN(n2063) );
  NAND2 U4056 ( .A1(n27390), .A2(n75), .ZN(n2065) );
  NAND2 U4057 ( .A1(n27390), .A2(n78), .ZN(n2067) );
  NAND2 U4058 ( .A1(n27390), .A2(n81), .ZN(n2069) );
  NAND2 U4059 ( .A1(n27390), .A2(n84), .ZN(n2071) );
  NAND2 U4060 ( .A1(n27390), .A2(n87), .ZN(n2073) );
  NAND2 U4061 ( .A1(n27390), .A2(n90), .ZN(n2075) );
  NAND2 U4062 ( .A1(n27390), .A2(n93), .ZN(n2077) );
  NAND2 U4063 ( .A1(n27391), .A2(n96), .ZN(n2079) );
  NAND2 U4064 ( .A1(n27391), .A2(n99), .ZN(n2081) );
  NAND2 U4065 ( .A1(n27391), .A2(n102), .ZN(n2083) );
  NAND2 U4066 ( .A1(n27391), .A2(n105), .ZN(n2085) );
  NAND2 U4067 ( .A1(n27391), .A2(n108), .ZN(n2087) );
  NAND2 U4068 ( .A1(n27391), .A2(n111), .ZN(n2089) );
  NAND2 U4069 ( .A1(n27391), .A2(n114), .ZN(n2091) );
  NAND2 U4070 ( .A1(n27391), .A2(n117), .ZN(n2093) );
  NAND2 U4071 ( .A1(n27391), .A2(n120), .ZN(n2095) );
  NAND2 U4072 ( .A1(n27391), .A2(n123), .ZN(n2097) );
  NAND2 U4073 ( .A1(n27391), .A2(n126), .ZN(n2099) );
  NAND2 U4074 ( .A1(n27391), .A2(n129), .ZN(n2101) );
  NAND2 U4075 ( .A1(n27390), .A2(n132), .ZN(n2103) );
  NAND2 U4076 ( .A1(n27391), .A2(n135), .ZN(n2105) );
  NAND2 U4077 ( .A1(n27389), .A2(n138), .ZN(n2107) );
  NAND2 U4078 ( .A1(n27390), .A2(n141), .ZN(n2109) );
  NAND2 U4079 ( .A1(n27391), .A2(n144), .ZN(n2111) );
  NAND2 U4080 ( .A1(n27389), .A2(n147), .ZN(n2113) );
  NAND2 U4081 ( .A1(n27390), .A2(n150), .ZN(n2115) );
  NAND2 U4082 ( .A1(n27391), .A2(n153), .ZN(n2117) );
  NAND2 U4083 ( .A1(n27389), .A2(n156), .ZN(n2119) );
  NAND2 U4084 ( .A1(n27390), .A2(n159), .ZN(n2121) );
  NAND2 U4085 ( .A1(n27391), .A2(n162), .ZN(n2123) );
  NAND2 U4086 ( .A1(n27389), .A2(n165), .ZN(n2125) );
  NAND2 U4087 ( .A1(n27391), .A2(n10), .ZN(n2127) );
  NAND2 U4088 ( .A1(n27389), .A2(n11), .ZN(n2129) );
  NAND2 U4089 ( .A1(n27389), .A2(n12), .ZN(n2131) );
  NAND2 U4090 ( .A1(n27390), .A2(n24), .ZN(n2133) );
  NAND2 U4091 ( .A1(n27391), .A2(n27), .ZN(n2135) );
  NAND2 U4092 ( .A1(n27390), .A2(n30), .ZN(n2137) );
  NAND2 U4093 ( .A1(n27389), .A2(n33), .ZN(n2139) );
  NAND2 U4094 ( .A1(n27390), .A2(n36), .ZN(n2141) );
  NAND2 U4095 ( .A1(n27391), .A2(n39), .ZN(n2143) );
  NAND2 U4096 ( .A1(n27391), .A2(n168), .ZN(n2145) );
  NAND2 U4097 ( .A1(n27389), .A2(n171), .ZN(n2147) );
  NAND2 U4098 ( .A1(n27390), .A2(n174), .ZN(n2149) );
  NAND2 U4099 ( .A1(n27386), .A2(n23), .ZN(n2159) );
  NAND2 U4100 ( .A1(n27386), .A2(n5), .ZN(n2162) );
  NAND2 U4101 ( .A1(n27386), .A2(n6), .ZN(n2164) );
  NAND2 U4102 ( .A1(n27386), .A2(n7), .ZN(n2166) );
  NAND2 U4103 ( .A1(n27386), .A2(n8), .ZN(n2168) );
  NAND2 U4104 ( .A1(n27386), .A2(n9), .ZN(n2170) );
  NAND2 U4105 ( .A1(n27386), .A2(n42), .ZN(n2172) );
  NAND2 U4106 ( .A1(n27386), .A2(n45), .ZN(n2174) );
  NAND2 U4107 ( .A1(n27386), .A2(n48), .ZN(n2176) );
  NAND2 U4108 ( .A1(n27386), .A2(n51), .ZN(n2178) );
  NAND2 U4109 ( .A1(n27386), .A2(n54), .ZN(n2180) );
  NAND2 U4110 ( .A1(n27386), .A2(n57), .ZN(n2182) );
  NAND2 U4111 ( .A1(n27387), .A2(n60), .ZN(n2184) );
  NAND2 U4112 ( .A1(n27387), .A2(n63), .ZN(n2186) );
  NAND2 U4113 ( .A1(n27387), .A2(n66), .ZN(n2188) );
  NAND2 U4114 ( .A1(n27387), .A2(n69), .ZN(n2190) );
  NAND2 U4115 ( .A1(n27387), .A2(n72), .ZN(n2192) );
  NAND2 U4116 ( .A1(n27387), .A2(n75), .ZN(n2194) );
  NAND2 U4117 ( .A1(n27387), .A2(n78), .ZN(n2196) );
  NAND2 U4118 ( .A1(n27387), .A2(n81), .ZN(n2198) );
  NAND2 U4119 ( .A1(n27387), .A2(n84), .ZN(n2200) );
  NAND2 U4120 ( .A1(n27387), .A2(n87), .ZN(n2202) );
  NAND2 U4121 ( .A1(n27387), .A2(n90), .ZN(n2204) );
  NAND2 U4122 ( .A1(n27387), .A2(n93), .ZN(n2206) );
  NAND2 U4123 ( .A1(n27388), .A2(n96), .ZN(n2208) );
  NAND2 U4124 ( .A1(n27388), .A2(n99), .ZN(n2210) );
  NAND2 U4125 ( .A1(n27388), .A2(n102), .ZN(n2212) );
  NAND2 U4126 ( .A1(n27388), .A2(n105), .ZN(n2214) );
  NAND2 U4127 ( .A1(n27388), .A2(n108), .ZN(n2216) );
  NAND2 U4128 ( .A1(n27388), .A2(n111), .ZN(n2218) );
  NAND2 U4129 ( .A1(n27388), .A2(n114), .ZN(n2220) );
  NAND2 U4130 ( .A1(n27388), .A2(n117), .ZN(n2222) );
  NAND2 U4131 ( .A1(n27388), .A2(n120), .ZN(n2224) );
  NAND2 U4132 ( .A1(n27388), .A2(n123), .ZN(n2226) );
  NAND2 U4133 ( .A1(n27388), .A2(n126), .ZN(n2228) );
  NAND2 U4134 ( .A1(n27388), .A2(n129), .ZN(n2230) );
  NAND2 U4135 ( .A1(n27387), .A2(n132), .ZN(n2232) );
  NAND2 U4136 ( .A1(n27388), .A2(n135), .ZN(n2234) );
  NAND2 U4137 ( .A1(n27386), .A2(n138), .ZN(n2236) );
  NAND2 U4138 ( .A1(n27387), .A2(n141), .ZN(n2238) );
  NAND2 U4139 ( .A1(n27388), .A2(n144), .ZN(n2240) );
  NAND2 U4140 ( .A1(n27386), .A2(n147), .ZN(n2242) );
  NAND2 U4141 ( .A1(n27387), .A2(n150), .ZN(n2244) );
  NAND2 U4142 ( .A1(n27388), .A2(n153), .ZN(n2246) );
  NAND2 U4143 ( .A1(n27386), .A2(n156), .ZN(n2248) );
  NAND2 U4144 ( .A1(n27387), .A2(n159), .ZN(n2250) );
  NAND2 U4145 ( .A1(n27388), .A2(n162), .ZN(n2252) );
  NAND2 U4146 ( .A1(n27386), .A2(n165), .ZN(n2254) );
  NAND2 U4147 ( .A1(n27388), .A2(n10), .ZN(n2256) );
  NAND2 U4148 ( .A1(n27386), .A2(n11), .ZN(n2258) );
  NAND2 U4149 ( .A1(n27386), .A2(n12), .ZN(n2260) );
  NAND2 U4150 ( .A1(n27387), .A2(n24), .ZN(n2262) );
  NAND2 U4151 ( .A1(n27388), .A2(n27), .ZN(n2264) );
  NAND2 U4152 ( .A1(n27387), .A2(n30), .ZN(n2266) );
  NAND2 U4153 ( .A1(n27386), .A2(n33), .ZN(n2268) );
  NAND2 U4154 ( .A1(n27387), .A2(n36), .ZN(n2270) );
  NAND2 U4155 ( .A1(n27388), .A2(n39), .ZN(n2272) );
  NAND2 U4156 ( .A1(n27388), .A2(n168), .ZN(n2274) );
  NAND2 U4157 ( .A1(n27386), .A2(n171), .ZN(n2276) );
  NAND2 U4158 ( .A1(n27387), .A2(n174), .ZN(n2278) );
  NAND2 U4159 ( .A1(n27383), .A2(n23), .ZN(n2289) );
  NAND2 U4160 ( .A1(n27383), .A2(n5), .ZN(n2292) );
  NAND2 U4161 ( .A1(n27383), .A2(n6), .ZN(n2294) );
  NAND2 U4162 ( .A1(n27383), .A2(n7), .ZN(n2296) );
  NAND2 U4163 ( .A1(n27383), .A2(n8), .ZN(n2298) );
  NAND2 U4164 ( .A1(n27383), .A2(n9), .ZN(n2300) );
  NAND2 U4165 ( .A1(n27383), .A2(n42), .ZN(n2302) );
  NAND2 U4166 ( .A1(n27383), .A2(n45), .ZN(n2304) );
  NAND2 U4167 ( .A1(n27383), .A2(n48), .ZN(n2306) );
  NAND2 U4168 ( .A1(n27383), .A2(n51), .ZN(n2308) );
  NAND2 U4169 ( .A1(n27383), .A2(n54), .ZN(n2310) );
  NAND2 U4170 ( .A1(n27383), .A2(n57), .ZN(n2312) );
  NAND2 U4171 ( .A1(n27384), .A2(n60), .ZN(n2314) );
  NAND2 U4172 ( .A1(n27384), .A2(n63), .ZN(n2316) );
  NAND2 U4173 ( .A1(n27384), .A2(n66), .ZN(n2318) );
  NAND2 U4174 ( .A1(n27384), .A2(n69), .ZN(n2320) );
  NAND2 U4175 ( .A1(n27384), .A2(n72), .ZN(n2322) );
  NAND2 U4176 ( .A1(n27384), .A2(n75), .ZN(n2324) );
  NAND2 U4177 ( .A1(n27384), .A2(n78), .ZN(n2326) );
  NAND2 U4178 ( .A1(n27384), .A2(n81), .ZN(n2328) );
  NAND2 U4179 ( .A1(n27384), .A2(n84), .ZN(n2330) );
  NAND2 U4180 ( .A1(n27384), .A2(n87), .ZN(n2332) );
  NAND2 U4181 ( .A1(n27384), .A2(n90), .ZN(n2334) );
  NAND2 U4182 ( .A1(n27384), .A2(n93), .ZN(n2336) );
  NAND2 U4183 ( .A1(n27385), .A2(n96), .ZN(n2338) );
  NAND2 U4184 ( .A1(n27385), .A2(n99), .ZN(n2340) );
  NAND2 U4185 ( .A1(n27385), .A2(n102), .ZN(n2342) );
  NAND2 U4186 ( .A1(n27385), .A2(n105), .ZN(n2344) );
  NAND2 U4187 ( .A1(n27385), .A2(n108), .ZN(n2346) );
  NAND2 U4188 ( .A1(n27385), .A2(n111), .ZN(n2348) );
  NAND2 U4189 ( .A1(n27385), .A2(n114), .ZN(n2350) );
  NAND2 U4190 ( .A1(n27385), .A2(n117), .ZN(n2352) );
  NAND2 U4191 ( .A1(n27385), .A2(n120), .ZN(n2354) );
  NAND2 U4192 ( .A1(n27385), .A2(n123), .ZN(n2356) );
  NAND2 U4193 ( .A1(n27385), .A2(n126), .ZN(n2358) );
  NAND2 U4194 ( .A1(n27385), .A2(n129), .ZN(n2360) );
  NAND2 U4195 ( .A1(n27384), .A2(n132), .ZN(n2362) );
  NAND2 U4196 ( .A1(n27385), .A2(n135), .ZN(n2364) );
  NAND2 U4197 ( .A1(n27383), .A2(n138), .ZN(n2366) );
  NAND2 U4198 ( .A1(n27384), .A2(n141), .ZN(n2368) );
  NAND2 U4199 ( .A1(n27385), .A2(n144), .ZN(n2370) );
  NAND2 U4200 ( .A1(n27383), .A2(n147), .ZN(n2372) );
  NAND2 U4201 ( .A1(n27384), .A2(n150), .ZN(n2374) );
  NAND2 U4202 ( .A1(n27385), .A2(n153), .ZN(n2376) );
  NAND2 U4203 ( .A1(n27383), .A2(n156), .ZN(n2378) );
  NAND2 U4204 ( .A1(n27384), .A2(n159), .ZN(n2380) );
  NAND2 U4205 ( .A1(n27385), .A2(n162), .ZN(n2382) );
  NAND2 U4206 ( .A1(n27383), .A2(n165), .ZN(n2384) );
  NAND2 U4207 ( .A1(n27385), .A2(n10), .ZN(n2386) );
  NAND2 U4208 ( .A1(n27383), .A2(n11), .ZN(n2388) );
  NAND2 U4209 ( .A1(n27383), .A2(n12), .ZN(n2390) );
  NAND2 U4210 ( .A1(n27384), .A2(n24), .ZN(n2392) );
  NAND2 U4211 ( .A1(n27385), .A2(n27), .ZN(n2394) );
  NAND2 U4212 ( .A1(n27384), .A2(n30), .ZN(n2396) );
  NAND2 U4213 ( .A1(n27383), .A2(n33), .ZN(n2398) );
  NAND2 U4214 ( .A1(n27384), .A2(n36), .ZN(n2400) );
  NAND2 U4215 ( .A1(n27385), .A2(n39), .ZN(n2402) );
  NAND2 U4216 ( .A1(n27385), .A2(n168), .ZN(n2404) );
  NAND2 U4217 ( .A1(n27383), .A2(n171), .ZN(n2406) );
  NAND2 U4218 ( .A1(n27384), .A2(n174), .ZN(n2408) );
  NAND2 U4219 ( .A1(n27380), .A2(n23), .ZN(n2418) );
  NAND2 U4220 ( .A1(n27380), .A2(n5), .ZN(n2421) );
  NAND2 U4221 ( .A1(n27380), .A2(n6), .ZN(n2423) );
  NAND2 U4222 ( .A1(n27380), .A2(n7), .ZN(n2425) );
  NAND2 U4223 ( .A1(n27380), .A2(n8), .ZN(n2427) );
  NAND2 U4224 ( .A1(n27380), .A2(n9), .ZN(n2429) );
  NAND2 U4225 ( .A1(n27380), .A2(n42), .ZN(n2431) );
  NAND2 U4226 ( .A1(n27380), .A2(n45), .ZN(n2433) );
  NAND2 U4227 ( .A1(n27380), .A2(n48), .ZN(n2435) );
  NAND2 U4228 ( .A1(n27380), .A2(n51), .ZN(n2437) );
  NAND2 U4229 ( .A1(n27380), .A2(n54), .ZN(n2439) );
  NAND2 U4230 ( .A1(n27380), .A2(n57), .ZN(n2441) );
  NAND2 U4231 ( .A1(n27381), .A2(n60), .ZN(n2443) );
  NAND2 U4232 ( .A1(n27381), .A2(n63), .ZN(n2445) );
  NAND2 U4233 ( .A1(n27381), .A2(n66), .ZN(n2447) );
  NAND2 U4234 ( .A1(n27381), .A2(n69), .ZN(n2449) );
  NAND2 U4235 ( .A1(n27381), .A2(n72), .ZN(n2451) );
  NAND2 U4236 ( .A1(n27381), .A2(n75), .ZN(n2453) );
  NAND2 U4237 ( .A1(n27381), .A2(n78), .ZN(n2455) );
  NAND2 U4238 ( .A1(n27381), .A2(n81), .ZN(n2457) );
  NAND2 U4239 ( .A1(n27381), .A2(n84), .ZN(n2459) );
  NAND2 U4240 ( .A1(n27381), .A2(n87), .ZN(n2461) );
  NAND2 U4241 ( .A1(n27381), .A2(n90), .ZN(n2463) );
  NAND2 U4242 ( .A1(n27381), .A2(n93), .ZN(n2465) );
  NAND2 U4243 ( .A1(n27382), .A2(n96), .ZN(n2467) );
  NAND2 U4244 ( .A1(n27382), .A2(n99), .ZN(n2469) );
  NAND2 U4245 ( .A1(n27382), .A2(n102), .ZN(n2471) );
  NAND2 U4246 ( .A1(n27382), .A2(n105), .ZN(n2473) );
  NAND2 U4247 ( .A1(n27382), .A2(n108), .ZN(n2475) );
  NAND2 U4248 ( .A1(n27382), .A2(n111), .ZN(n2477) );
  NAND2 U4249 ( .A1(n27382), .A2(n114), .ZN(n2479) );
  NAND2 U4250 ( .A1(n27382), .A2(n117), .ZN(n2481) );
  NAND2 U4251 ( .A1(n27382), .A2(n120), .ZN(n2483) );
  NAND2 U4252 ( .A1(n27382), .A2(n123), .ZN(n2485) );
  NAND2 U4253 ( .A1(n27382), .A2(n126), .ZN(n2487) );
  NAND2 U4254 ( .A1(n27382), .A2(n129), .ZN(n2489) );
  NAND2 U4255 ( .A1(n27381), .A2(n132), .ZN(n2491) );
  NAND2 U4256 ( .A1(n27382), .A2(n135), .ZN(n2493) );
  NAND2 U4257 ( .A1(n27380), .A2(n138), .ZN(n2495) );
  NAND2 U4258 ( .A1(n27381), .A2(n141), .ZN(n2497) );
  NAND2 U4259 ( .A1(n27382), .A2(n144), .ZN(n2499) );
  NAND2 U4260 ( .A1(n27380), .A2(n147), .ZN(n2501) );
  NAND2 U4261 ( .A1(n27381), .A2(n150), .ZN(n2503) );
  NAND2 U4262 ( .A1(n27382), .A2(n153), .ZN(n2505) );
  NAND2 U4263 ( .A1(n27380), .A2(n156), .ZN(n2507) );
  NAND2 U4264 ( .A1(n27381), .A2(n159), .ZN(n2509) );
  NAND2 U4265 ( .A1(n27382), .A2(n162), .ZN(n2511) );
  NAND2 U4266 ( .A1(n27380), .A2(n165), .ZN(n2513) );
  NAND2 U4267 ( .A1(n27382), .A2(n10), .ZN(n2515) );
  NAND2 U4268 ( .A1(n27380), .A2(n11), .ZN(n2517) );
  NAND2 U4269 ( .A1(n27380), .A2(n12), .ZN(n2519) );
  NAND2 U4270 ( .A1(n27381), .A2(n24), .ZN(n2521) );
  NAND2 U4271 ( .A1(n27382), .A2(n27), .ZN(n2523) );
  NAND2 U4272 ( .A1(n27381), .A2(n30), .ZN(n2525) );
  NAND2 U4273 ( .A1(n27380), .A2(n33), .ZN(n2527) );
  NAND2 U4274 ( .A1(n27381), .A2(n36), .ZN(n2529) );
  NAND2 U4275 ( .A1(n27382), .A2(n39), .ZN(n2531) );
  NAND2 U4276 ( .A1(n27382), .A2(n168), .ZN(n2533) );
  NAND2 U4277 ( .A1(n27380), .A2(n171), .ZN(n2535) );
  NAND2 U4278 ( .A1(n27381), .A2(n174), .ZN(n2537) );
  NAND2 U4279 ( .A1(n27377), .A2(n23), .ZN(n2547) );
  NAND2 U4280 ( .A1(n27377), .A2(n5), .ZN(n2550) );
  NAND2 U4281 ( .A1(n27377), .A2(n6), .ZN(n2552) );
  NAND2 U4282 ( .A1(n27377), .A2(n7), .ZN(n2554) );
  NAND2 U4283 ( .A1(n27377), .A2(n8), .ZN(n2556) );
  NAND2 U4284 ( .A1(n27377), .A2(n9), .ZN(n2558) );
  NAND2 U4285 ( .A1(n27377), .A2(n42), .ZN(n2560) );
  NAND2 U4286 ( .A1(n27377), .A2(n45), .ZN(n2562) );
  NAND2 U4287 ( .A1(n27377), .A2(n48), .ZN(n2564) );
  NAND2 U4288 ( .A1(n27377), .A2(n51), .ZN(n2566) );
  NAND2 U4289 ( .A1(n27377), .A2(n54), .ZN(n2568) );
  NAND2 U4290 ( .A1(n27377), .A2(n57), .ZN(n2570) );
  NAND2 U4291 ( .A1(n27378), .A2(n60), .ZN(n2572) );
  NAND2 U4292 ( .A1(n27378), .A2(n63), .ZN(n2574) );
  NAND2 U4293 ( .A1(n27378), .A2(n66), .ZN(n2576) );
  NAND2 U4294 ( .A1(n27378), .A2(n69), .ZN(n2578) );
  NAND2 U4295 ( .A1(n27378), .A2(n72), .ZN(n2580) );
  NAND2 U4296 ( .A1(n27378), .A2(n75), .ZN(n2582) );
  NAND2 U4297 ( .A1(n27378), .A2(n78), .ZN(n2584) );
  NAND2 U4298 ( .A1(n27378), .A2(n81), .ZN(n2586) );
  NAND2 U4299 ( .A1(n27378), .A2(n84), .ZN(n2588) );
  NAND2 U4300 ( .A1(n27378), .A2(n87), .ZN(n2590) );
  NAND2 U4301 ( .A1(n27378), .A2(n90), .ZN(n2592) );
  NAND2 U4302 ( .A1(n27378), .A2(n93), .ZN(n2594) );
  NAND2 U4303 ( .A1(n27379), .A2(n96), .ZN(n2596) );
  NAND2 U4304 ( .A1(n27379), .A2(n99), .ZN(n2598) );
  NAND2 U4305 ( .A1(n27379), .A2(n102), .ZN(n2600) );
  NAND2 U4306 ( .A1(n27379), .A2(n105), .ZN(n2602) );
  NAND2 U4307 ( .A1(n27379), .A2(n108), .ZN(n2604) );
  NAND2 U4308 ( .A1(n27379), .A2(n111), .ZN(n2606) );
  NAND2 U4309 ( .A1(n27379), .A2(n114), .ZN(n2608) );
  NAND2 U4310 ( .A1(n27379), .A2(n117), .ZN(n2610) );
  NAND2 U4311 ( .A1(n27379), .A2(n120), .ZN(n2612) );
  NAND2 U4312 ( .A1(n27379), .A2(n123), .ZN(n2614) );
  NAND2 U4313 ( .A1(n27379), .A2(n126), .ZN(n2616) );
  NAND2 U4314 ( .A1(n27379), .A2(n129), .ZN(n2618) );
  NAND2 U4315 ( .A1(n27378), .A2(n132), .ZN(n2620) );
  NAND2 U4316 ( .A1(n27379), .A2(n135), .ZN(n2622) );
  NAND2 U4317 ( .A1(n27377), .A2(n138), .ZN(n2624) );
  NAND2 U4318 ( .A1(n27378), .A2(n141), .ZN(n2626) );
  NAND2 U4319 ( .A1(n27379), .A2(n144), .ZN(n2628) );
  NAND2 U4320 ( .A1(n27377), .A2(n147), .ZN(n2630) );
  NAND2 U4321 ( .A1(n27378), .A2(n150), .ZN(n2632) );
  NAND2 U4322 ( .A1(n27379), .A2(n153), .ZN(n2634) );
  NAND2 U4323 ( .A1(n27377), .A2(n156), .ZN(n2636) );
  NAND2 U4324 ( .A1(n27378), .A2(n159), .ZN(n2638) );
  NAND2 U4325 ( .A1(n27379), .A2(n162), .ZN(n2640) );
  NAND2 U4326 ( .A1(n27377), .A2(n165), .ZN(n2642) );
  NAND2 U4327 ( .A1(n27379), .A2(n10), .ZN(n2644) );
  NAND2 U4328 ( .A1(n27377), .A2(n11), .ZN(n2646) );
  NAND2 U4329 ( .A1(n27377), .A2(n12), .ZN(n2648) );
  NAND2 U4330 ( .A1(n27378), .A2(n24), .ZN(n2650) );
  NAND2 U4331 ( .A1(n27379), .A2(n27), .ZN(n2652) );
  NAND2 U4332 ( .A1(n27378), .A2(n30), .ZN(n2654) );
  NAND2 U4333 ( .A1(n27377), .A2(n33), .ZN(n2656) );
  NAND2 U4334 ( .A1(n27378), .A2(n36), .ZN(n2658) );
  NAND2 U4335 ( .A1(n27379), .A2(n39), .ZN(n2660) );
  NAND2 U4336 ( .A1(n27379), .A2(n168), .ZN(n2662) );
  NAND2 U4337 ( .A1(n27377), .A2(n171), .ZN(n2664) );
  NAND2 U4338 ( .A1(n27378), .A2(n174), .ZN(n2666) );
  NAND2 U4339 ( .A1(n27374), .A2(n23), .ZN(n2676) );
  NAND2 U4340 ( .A1(n27371), .A2(n23), .ZN(n2805) );
  NAND2 U4341 ( .A1(n27369), .A2(n23), .ZN(n2934) );
  NAND2 U4342 ( .A1(n27365), .A2(n23), .ZN(n3063) );
  NAND2 U4343 ( .A1(n27364), .A2(n23), .ZN(n3192) );
  NAND2 U4344 ( .A1(n27359), .A2(n23), .ZN(n3322) );
  NAND2 U4345 ( .A1(n27356), .A2(n23), .ZN(n3451) );
  NAND2 U4346 ( .A1(n27353), .A2(n23), .ZN(n3580) );
  NAND2 U4347 ( .A1(n27350), .A2(n23), .ZN(n3709) );
  NAND2 U4348 ( .A1(n27347), .A2(n23), .ZN(n3838) );
  NAND2 U4349 ( .A1(n27344), .A2(n23), .ZN(n3967) );
  NAND2 U4350 ( .A1(n27341), .A2(n23), .ZN(n4096) );
  NAND2 U4351 ( .A1(n5), .A2(n27434), .ZN(n25) );
  NAND2 U4352 ( .A1(n6), .A2(n27434), .ZN(n28) );
  NAND2 U4353 ( .A1(n7), .A2(n27434), .ZN(n31) );
  NAND2 U4354 ( .A1(n8), .A2(n27434), .ZN(n34) );
  NAND2 U4355 ( .A1(n9), .A2(n27434), .ZN(n37) );
  NAND2 U4356 ( .A1(n42), .A2(n27434), .ZN(n40) );
  NAND2 U4357 ( .A1(n45), .A2(n27434), .ZN(n43) );
  NAND2 U4358 ( .A1(n48), .A2(n27434), .ZN(n46) );
  NAND2 U4359 ( .A1(n51), .A2(n27434), .ZN(n49) );
  NAND2 U4360 ( .A1(n54), .A2(n27434), .ZN(n52) );
  NAND2 U4361 ( .A1(n57), .A2(n27434), .ZN(n55) );
  NAND2 U4362 ( .A1(n60), .A2(n27435), .ZN(n58) );
  NAND2 U4363 ( .A1(n63), .A2(n27435), .ZN(n61) );
  NAND2 U4364 ( .A1(n66), .A2(n27435), .ZN(n64) );
  NAND2 U4365 ( .A1(n69), .A2(n27435), .ZN(n67) );
  NAND2 U4366 ( .A1(n72), .A2(n27435), .ZN(n70) );
  NAND2 U4367 ( .A1(n75), .A2(n27435), .ZN(n73) );
  NAND2 U4368 ( .A1(n78), .A2(n27435), .ZN(n76) );
  NAND2 U4369 ( .A1(n81), .A2(n27435), .ZN(n79) );
  NAND2 U4370 ( .A1(n84), .A2(n27435), .ZN(n82) );
  NAND2 U4371 ( .A1(n87), .A2(n27435), .ZN(n85) );
  NAND2 U4372 ( .A1(n90), .A2(n27435), .ZN(n88) );
  NAND2 U4373 ( .A1(n93), .A2(n27435), .ZN(n91) );
  NAND2 U4374 ( .A1(n96), .A2(n27436), .ZN(n94) );
  NAND2 U4375 ( .A1(n99), .A2(n27436), .ZN(n97) );
  NAND2 U4376 ( .A1(n102), .A2(n27436), .ZN(n100) );
  NAND2 U4377 ( .A1(n105), .A2(n27436), .ZN(n103) );
  NAND2 U4378 ( .A1(n108), .A2(n27436), .ZN(n106) );
  NAND2 U4379 ( .A1(n111), .A2(n27436), .ZN(n109) );
  NAND2 U4380 ( .A1(n114), .A2(n27436), .ZN(n112) );
  NAND2 U4381 ( .A1(n117), .A2(n27436), .ZN(n115) );
  NAND2 U4382 ( .A1(n120), .A2(n27436), .ZN(n118) );
  NAND2 U4383 ( .A1(n123), .A2(n27436), .ZN(n121) );
  NAND2 U4384 ( .A1(n126), .A2(n27436), .ZN(n124) );
  NAND2 U4385 ( .A1(n129), .A2(n27436), .ZN(n127) );
  NAND2 U4386 ( .A1(n132), .A2(n27435), .ZN(n130) );
  NAND2 U4387 ( .A1(n135), .A2(n27435), .ZN(n133) );
  NAND2 U4388 ( .A1(n138), .A2(n27434), .ZN(n136) );
  NAND2 U4389 ( .A1(n141), .A2(n27436), .ZN(n139) );
  NAND2 U4390 ( .A1(n144), .A2(n27435), .ZN(n142) );
  NAND2 U4391 ( .A1(n147), .A2(n27434), .ZN(n145) );
  NAND2 U4392 ( .A1(n150), .A2(n27436), .ZN(n148) );
  NAND2 U4393 ( .A1(n153), .A2(n27435), .ZN(n151) );
  NAND2 U4394 ( .A1(n156), .A2(n27434), .ZN(n154) );
  NAND2 U4395 ( .A1(n159), .A2(n27434), .ZN(n157) );
  NAND2 U4396 ( .A1(n162), .A2(n27436), .ZN(n160) );
  NAND2 U4397 ( .A1(n165), .A2(n27435), .ZN(n163) );
  NAND2 U4398 ( .A1(n10), .A2(n27434), .ZN(n166) );
  NAND2 U4399 ( .A1(n11), .A2(n27436), .ZN(n169) );
  NAND2 U4400 ( .A1(n12), .A2(n27435), .ZN(n172) );
  NAND2 U4401 ( .A1(n24), .A2(n27434), .ZN(n175) );
  NAND2 U4402 ( .A1(n27), .A2(n27436), .ZN(n178) );
  NAND2 U4403 ( .A1(n30), .A2(n27435), .ZN(n181) );
  NAND2 U4404 ( .A1(n33), .A2(n27434), .ZN(n184) );
  NAND2 U4405 ( .A1(n36), .A2(n27436), .ZN(n187) );
  NAND2 U4406 ( .A1(n39), .A2(n27436), .ZN(n190) );
  NAND2 U4407 ( .A1(n168), .A2(n27434), .ZN(n193) );
  NAND2 U4408 ( .A1(n171), .A2(n27436), .ZN(n196) );
  NAND2 U4409 ( .A1(n174), .A2(n27435), .ZN(n199) );
  NAND2 U4410 ( .A1(n1), .A2(n27435), .ZN(n202) );
  NAND2 U4411 ( .A1(n2), .A2(n27434), .ZN(n205) );
  NAND2 U4412 ( .A1(n3), .A2(n27434), .ZN(n208) );
  NAND2 U4413 ( .A1(n4), .A2(n27436), .ZN(n211) );
  NAND2 U4414 ( .A1(n27432), .A2(n1), .ZN(n337) );
  NAND2 U4415 ( .A1(n27432), .A2(n2), .ZN(n339) );
  NAND2 U4416 ( .A1(n27433), .A2(n3), .ZN(n341) );
  NAND2 U4417 ( .A1(n27431), .A2(n4), .ZN(n343) );
  NAND2 U4418 ( .A1(n27429), .A2(n1), .ZN(n467) );
  NAND2 U4419 ( .A1(n27429), .A2(n2), .ZN(n469) );
  NAND2 U4420 ( .A1(n27430), .A2(n3), .ZN(n471) );
  NAND2 U4421 ( .A1(n27428), .A2(n4), .ZN(n473) );
  NAND2 U4422 ( .A1(n27426), .A2(n1), .ZN(n597) );
  NAND2 U4423 ( .A1(n27426), .A2(n2), .ZN(n599) );
  NAND2 U4424 ( .A1(n27427), .A2(n3), .ZN(n601) );
  NAND2 U4425 ( .A1(n27425), .A2(n4), .ZN(n603) );
  NAND2 U4426 ( .A1(n27423), .A2(n1), .ZN(n727) );
  NAND2 U4427 ( .A1(n27423), .A2(n2), .ZN(n729) );
  NAND2 U4428 ( .A1(n27424), .A2(n3), .ZN(n731) );
  NAND2 U4429 ( .A1(n27422), .A2(n4), .ZN(n733) );
  NAND2 U4430 ( .A1(n27420), .A2(n1), .ZN(n857) );
  NAND2 U4431 ( .A1(n27420), .A2(n2), .ZN(n859) );
  NAND2 U4432 ( .A1(n27421), .A2(n3), .ZN(n861) );
  NAND2 U4433 ( .A1(n27419), .A2(n4), .ZN(n863) );
  NAND2 U4434 ( .A1(n27417), .A2(n1), .ZN(n987) );
  NAND2 U4435 ( .A1(n27417), .A2(n2), .ZN(n989) );
  NAND2 U4436 ( .A1(n27418), .A2(n3), .ZN(n991) );
  NAND2 U4437 ( .A1(n27416), .A2(n4), .ZN(n993) );
  NAND2 U4438 ( .A1(n27414), .A2(n1), .ZN(n1117) );
  NAND2 U4439 ( .A1(n27414), .A2(n2), .ZN(n1119) );
  NAND2 U4440 ( .A1(n27415), .A2(n3), .ZN(n1121) );
  NAND2 U4441 ( .A1(n27412), .A2(n1), .ZN(n1247) );
  NAND2 U4442 ( .A1(n27412), .A2(n2), .ZN(n1249) );
  NAND2 U4443 ( .A1(n27410), .A2(n3), .ZN(n1251) );
  NAND2 U4444 ( .A1(n27411), .A2(n4), .ZN(n1253) );
  NAND2 U4445 ( .A1(n27409), .A2(n1), .ZN(n1377) );
  NAND2 U4446 ( .A1(n27409), .A2(n2), .ZN(n1379) );
  NAND2 U4447 ( .A1(n27407), .A2(n3), .ZN(n1381) );
  NAND2 U4448 ( .A1(n27408), .A2(n4), .ZN(n1383) );
  NAND2 U4449 ( .A1(n27406), .A2(n1), .ZN(n1506) );
  NAND2 U4450 ( .A1(n27406), .A2(n2), .ZN(n1508) );
  NAND2 U4451 ( .A1(n27404), .A2(n3), .ZN(n1510) );
  NAND2 U4452 ( .A1(n27405), .A2(n4), .ZN(n1512) );
  NAND2 U4453 ( .A1(n27403), .A2(n1), .ZN(n1635) );
  NAND2 U4454 ( .A1(n27403), .A2(n2), .ZN(n1637) );
  NAND2 U4455 ( .A1(n27401), .A2(n3), .ZN(n1639) );
  NAND2 U4456 ( .A1(n27402), .A2(n4), .ZN(n1641) );
  NAND2 U4457 ( .A1(n27400), .A2(n1), .ZN(n1764) );
  NAND2 U4458 ( .A1(n27400), .A2(n2), .ZN(n1766) );
  NAND2 U4459 ( .A1(n27398), .A2(n3), .ZN(n1768) );
  NAND2 U4460 ( .A1(n27399), .A2(n4), .ZN(n1770) );
  NAND2 U4461 ( .A1(n27397), .A2(n1), .ZN(n1893) );
  NAND2 U4462 ( .A1(n27397), .A2(n2), .ZN(n1895) );
  NAND2 U4463 ( .A1(n27395), .A2(n3), .ZN(n1897) );
  NAND2 U4464 ( .A1(n27396), .A2(n4), .ZN(n1899) );
  NAND2 U4465 ( .A1(n27394), .A2(n1), .ZN(n2022) );
  NAND2 U4466 ( .A1(n27394), .A2(n2), .ZN(n2024) );
  NAND2 U4467 ( .A1(n27392), .A2(n3), .ZN(n2026) );
  NAND2 U4468 ( .A1(n27393), .A2(n4), .ZN(n2028) );
  NAND2 U4469 ( .A1(n27391), .A2(n1), .ZN(n2151) );
  NAND2 U4470 ( .A1(n27391), .A2(n2), .ZN(n2153) );
  NAND2 U4471 ( .A1(n27389), .A2(n3), .ZN(n2155) );
  NAND2 U4472 ( .A1(n27388), .A2(n1), .ZN(n2280) );
  NAND2 U4473 ( .A1(n27388), .A2(n2), .ZN(n2282) );
  NAND2 U4474 ( .A1(n27386), .A2(n3), .ZN(n2284) );
  NAND2 U4475 ( .A1(n27387), .A2(n4), .ZN(n2286) );
  NAND2 U4476 ( .A1(n27385), .A2(n1), .ZN(n2410) );
  NAND2 U4477 ( .A1(n27385), .A2(n2), .ZN(n2412) );
  NAND2 U4478 ( .A1(n27383), .A2(n3), .ZN(n2414) );
  NAND2 U4479 ( .A1(n27384), .A2(n4), .ZN(n2416) );
  NAND2 U4480 ( .A1(n27382), .A2(n1), .ZN(n2539) );
  NAND2 U4481 ( .A1(n27382), .A2(n2), .ZN(n2541) );
  NAND2 U4482 ( .A1(n27380), .A2(n3), .ZN(n2543) );
  NAND2 U4483 ( .A1(n27381), .A2(n4), .ZN(n2545) );
  NAND2 U4484 ( .A1(n27379), .A2(n1), .ZN(n2668) );
  NAND2 U4485 ( .A1(n27379), .A2(n2), .ZN(n2670) );
  NAND2 U4486 ( .A1(n27377), .A2(n3), .ZN(n2672) );
  NAND2 U4487 ( .A1(n27378), .A2(n4), .ZN(n2674) );
  I_NAND2 U4488 ( .A1(n3190), .B1(n29481), .ZN(n3191) );
  I_NAND2 U4489 ( .A1(n4239), .B1(n29439), .ZN(n4240) );
  BUF U4490 ( .I(n29494), .Z(n29492) );
  NAND2 U4491 ( .A1(n27413), .A2(n4), .ZN(n1123) );
  NAND2 U4492 ( .A1(n27390), .A2(n4), .ZN(n2157) );
  BUF U4493 ( .I(n29494), .Z(n29493) );
  BUF U4494 ( .I(n29494), .Z(n29491) );
  BUF U4495 ( .I(n29578), .Z(n29552) );
  BUF U4496 ( .I(n29578), .Z(n29553) );
  BUF U4497 ( .I(n29576), .Z(n29557) );
  BUF U4498 ( .I(n29576), .Z(n29558) );
  BUF U4499 ( .I(n29576), .Z(n29559) );
  BUF U4500 ( .I(n29575), .Z(n29560) );
  BUF U4501 ( .I(n29577), .Z(n29554) );
  BUF U4502 ( .I(n29577), .Z(n29555) );
  BUF U4503 ( .I(n29577), .Z(n29556) );
  BUF U4504 ( .I(n29573), .Z(n29567) );
  BUF U4505 ( .I(n29573), .Z(n29568) );
  BUF U4506 ( .I(n29574), .Z(n29563) );
  BUF U4507 ( .I(n29575), .Z(n29561) );
  BUF U4508 ( .I(n29575), .Z(n29562) );
  BUF U4509 ( .I(n29573), .Z(n29566) );
  BUF U4510 ( .I(n29574), .Z(n29564) );
  BUF U4511 ( .I(n29574), .Z(n29565) );
  BUF U4512 ( .I(n29570), .Z(n29496) );
  BUF U4513 ( .I(n29570), .Z(n29495) );
  BUF U4514 ( .I(n29569), .Z(n29500) );
  BUF U4515 ( .I(n29569), .Z(n29499) );
  BUF U4516 ( .I(n29569), .Z(n29498) );
  BUF U4517 ( .I(n29570), .Z(n29497) );
  BUF U4518 ( .I(n27023), .Z(n27024) );
  BUF U4519 ( .I(n27023), .Z(n27025) );
  BUF U4520 ( .I(n26878), .Z(n26892) );
  BUF U4521 ( .I(n26403), .Z(n26417) );
  BUF U4522 ( .I(n26878), .Z(n26891) );
  BUF U4523 ( .I(n26403), .Z(n26416) );
  BUF U4524 ( .I(n26877), .Z(n26896) );
  BUF U4525 ( .I(n26402), .Z(n26421) );
  BUF U4526 ( .I(n26875), .Z(n26901) );
  BUF U4527 ( .I(n26400), .Z(n26426) );
  BUF U4528 ( .I(n26875), .Z(n26900) );
  BUF U4529 ( .I(n26400), .Z(n26425) );
  BUF U4530 ( .I(n26874), .Z(n26905) );
  BUF U4531 ( .I(n26399), .Z(n26430) );
  BUF U4532 ( .I(n26872), .Z(n26909) );
  BUF U4533 ( .I(n26397), .Z(n26434) );
  BUF U4534 ( .I(n26871), .Z(n26914) );
  BUF U4535 ( .I(n26396), .Z(n26439) );
  BUF U4536 ( .I(n26871), .Z(n26913) );
  BUF U4537 ( .I(n26396), .Z(n26438) );
  BUF U4538 ( .I(n26883), .Z(n27021) );
  BUF U4539 ( .I(n26883), .Z(n27022) );
  BUF U4540 ( .I(n26888), .Z(n27007) );
  BUF U4541 ( .I(n26887), .Z(n27008) );
  BUF U4542 ( .I(n26887), .Z(n27009) );
  BUF U4543 ( .I(n26887), .Z(n27010) );
  BUF U4544 ( .I(n26877), .Z(n26895) );
  BUF U4545 ( .I(n26402), .Z(n26420) );
  BUF U4546 ( .I(n26877), .Z(n26894) );
  BUF U4547 ( .I(n26878), .Z(n26893) );
  BUF U4548 ( .I(n26403), .Z(n26418) );
  BUF U4549 ( .I(n26876), .Z(n26897) );
  BUF U4550 ( .I(n26401), .Z(n26422) );
  BUF U4551 ( .I(n26876), .Z(n26899) );
  BUF U4552 ( .I(n26401), .Z(n26424) );
  BUF U4553 ( .I(n26876), .Z(n26898) );
  BUF U4554 ( .I(n26874), .Z(n26904) );
  BUF U4555 ( .I(n26399), .Z(n26429) );
  BUF U4556 ( .I(n26874), .Z(n26903) );
  BUF U4557 ( .I(n26399), .Z(n26428) );
  BUF U4558 ( .I(n26875), .Z(n26902) );
  BUF U4559 ( .I(n26400), .Z(n26427) );
  BUF U4560 ( .I(n26873), .Z(n26908) );
  BUF U4561 ( .I(n26398), .Z(n26433) );
  BUF U4562 ( .I(n26873), .Z(n26907) );
  BUF U4563 ( .I(n26873), .Z(n26906) );
  BUF U4564 ( .I(n26398), .Z(n26431) );
  BUF U4565 ( .I(n26872), .Z(n26910) );
  BUF U4566 ( .I(n26871), .Z(n26912) );
  BUF U4567 ( .I(n26396), .Z(n26437) );
  BUF U4568 ( .I(n26872), .Z(n26911) );
  BUF U4569 ( .I(n26397), .Z(n26436) );
  BUF U4570 ( .I(n26870), .Z(n26917) );
  BUF U4571 ( .I(n26395), .Z(n26442) );
  BUF U4572 ( .I(n26870), .Z(n26916) );
  BUF U4573 ( .I(n26870), .Z(n26915) );
  BUF U4574 ( .I(n26395), .Z(n26440) );
  BUF U4575 ( .I(n26886), .Z(n27011) );
  BUF U4576 ( .I(n26411), .Z(n26536) );
  BUF U4577 ( .I(n26886), .Z(n27012) );
  BUF U4578 ( .I(n26411), .Z(n26537) );
  BUF U4579 ( .I(n26884), .Z(n27018) );
  BUF U4580 ( .I(n26883), .Z(n27020) );
  BUF U4581 ( .I(n26884), .Z(n27019) );
  BUF U4582 ( .I(n26886), .Z(n27013) );
  BUF U4583 ( .I(n26885), .Z(n27014) );
  BUF U4584 ( .I(n26885), .Z(n27015) );
  BUF U4585 ( .I(n26884), .Z(n27017) );
  BUF U4586 ( .I(n26885), .Z(n27016) );
  BUF U4587 ( .I(n26890), .Z(n26999) );
  BUF U4588 ( .I(n26415), .Z(n26524) );
  BUF U4589 ( .I(n26889), .Z(n27004) );
  BUF U4590 ( .I(n26888), .Z(n27005) );
  BUF U4591 ( .I(n26888), .Z(n27006) );
  BUF U4592 ( .I(n26890), .Z(n27000) );
  BUF U4593 ( .I(n26890), .Z(n27001) );
  BUF U4594 ( .I(n26889), .Z(n27002) );
  BUF U4595 ( .I(n26889), .Z(n27003) );
  BUF U4596 ( .I(n26193), .Z(n26196) );
  BUF U4597 ( .I(n26193), .Z(n26195) );
  BUF U4598 ( .I(n26189), .Z(n26206) );
  BUF U4599 ( .I(n26190), .Z(n26205) );
  BUF U4600 ( .I(n26186), .Z(n26216) );
  BUF U4601 ( .I(n26186), .Z(n26215) );
  BUF U4602 ( .I(n26187), .Z(n26214) );
  BUF U4603 ( .I(n26183), .Z(n26225) );
  BUF U4604 ( .I(n26183), .Z(n26224) );
  BUF U4605 ( .I(n26180), .Z(n26235) );
  BUF U4606 ( .I(n26180), .Z(n26234) );
  BUF U4607 ( .I(n26176), .Z(n26245) );
  BUF U4608 ( .I(n26177), .Z(n26244) );
  BUF U4609 ( .I(n26173), .Z(n26255) );
  BUF U4610 ( .I(n26173), .Z(n26254) );
  BUF U4611 ( .I(n26170), .Z(n26265) );
  BUF U4612 ( .I(n26170), .Z(n26264) );
  BUF U4613 ( .I(n26190), .Z(n26204) );
  BUF U4614 ( .I(n26190), .Z(n26203) );
  BUF U4615 ( .I(n26191), .Z(n26202) );
  BUF U4616 ( .I(n26192), .Z(n26198) );
  BUF U4617 ( .I(n26192), .Z(n26197) );
  BUF U4618 ( .I(n26191), .Z(n26201) );
  BUF U4619 ( .I(n26191), .Z(n26200) );
  BUF U4620 ( .I(n26192), .Z(n26199) );
  BUF U4621 ( .I(n26187), .Z(n26213) );
  BUF U4622 ( .I(n26187), .Z(n26212) );
  BUF U4623 ( .I(n26189), .Z(n26208) );
  BUF U4624 ( .I(n26189), .Z(n26207) );
  BUF U4625 ( .I(n26188), .Z(n26211) );
  BUF U4626 ( .I(n26188), .Z(n26210) );
  BUF U4627 ( .I(n26188), .Z(n26209) );
  BUF U4628 ( .I(n26184), .Z(n26223) );
  BUF U4629 ( .I(n26184), .Z(n26222) );
  BUF U4630 ( .I(n26186), .Z(n26217) );
  BUF U4631 ( .I(n26184), .Z(n26221) );
  BUF U4632 ( .I(n26185), .Z(n26220) );
  BUF U4633 ( .I(n26185), .Z(n26218) );
  BUF U4634 ( .I(n26185), .Z(n26219) );
  BUF U4635 ( .I(n26180), .Z(n26233) );
  BUF U4636 ( .I(n26181), .Z(n26232) );
  BUF U4637 ( .I(n26183), .Z(n26226) );
  BUF U4638 ( .I(n26182), .Z(n26227) );
  BUF U4639 ( .I(n26181), .Z(n26231) );
  BUF U4640 ( .I(n26181), .Z(n26230) );
  BUF U4641 ( .I(n26182), .Z(n26228) );
  BUF U4642 ( .I(n26182), .Z(n26229) );
  BUF U4643 ( .I(n26177), .Z(n26243) );
  BUF U4644 ( .I(n26177), .Z(n26242) );
  BUF U4645 ( .I(n26178), .Z(n26241) );
  BUF U4646 ( .I(n26179), .Z(n26236) );
  BUF U4647 ( .I(n26179), .Z(n26237) );
  BUF U4648 ( .I(n26178), .Z(n26240) );
  BUF U4649 ( .I(n26178), .Z(n26239) );
  BUF U4650 ( .I(n26179), .Z(n26238) );
  BUF U4651 ( .I(n26174), .Z(n26253) );
  BUF U4652 ( .I(n26174), .Z(n26252) );
  BUF U4653 ( .I(n26174), .Z(n26251) );
  BUF U4654 ( .I(n26176), .Z(n26247) );
  BUF U4655 ( .I(n26176), .Z(n26246) );
  BUF U4656 ( .I(n26175), .Z(n26250) );
  BUF U4657 ( .I(n26175), .Z(n26249) );
  BUF U4658 ( .I(n26175), .Z(n26248) );
  BUF U4659 ( .I(n26170), .Z(n26263) );
  BUF U4660 ( .I(n26171), .Z(n26262) );
  BUF U4661 ( .I(n26171), .Z(n26261) );
  BUF U4662 ( .I(n26172), .Z(n26257) );
  BUF U4663 ( .I(n26173), .Z(n26256) );
  BUF U4664 ( .I(n26171), .Z(n26260) );
  BUF U4665 ( .I(n26172), .Z(n26259) );
  BUF U4666 ( .I(n26172), .Z(n26258) );
  BUF U4667 ( .I(n26168), .Z(n26271) );
  BUF U4668 ( .I(n26169), .Z(n26267) );
  BUF U4669 ( .I(n26169), .Z(n26266) );
  BUF U4670 ( .I(n26168), .Z(n26270) );
  BUF U4671 ( .I(n26168), .Z(n26269) );
  BUF U4672 ( .I(n26169), .Z(n26268) );
  BUF U4673 ( .I(n26193), .Z(n26194) );
  BUF U4674 ( .I(n26548), .Z(n26549) );
  BUF U4675 ( .I(n26548), .Z(n26550) );
  BUF U4676 ( .I(n26311), .Z(n26314) );
  BUF U4677 ( .I(n26311), .Z(n26313) );
  BUF U4678 ( .I(n26307), .Z(n26324) );
  BUF U4679 ( .I(n26308), .Z(n26323) );
  BUF U4680 ( .I(n26304), .Z(n26334) );
  BUF U4681 ( .I(n26304), .Z(n26333) );
  BUF U4682 ( .I(n26305), .Z(n26332) );
  BUF U4683 ( .I(n26301), .Z(n26343) );
  BUF U4684 ( .I(n26301), .Z(n26342) );
  BUF U4685 ( .I(n26298), .Z(n26353) );
  BUF U4686 ( .I(n26298), .Z(n26352) );
  BUF U4687 ( .I(n26294), .Z(n26363) );
  BUF U4688 ( .I(n26295), .Z(n26362) );
  BUF U4689 ( .I(n26291), .Z(n26373) );
  BUF U4690 ( .I(n26291), .Z(n26372) );
  BUF U4691 ( .I(n26288), .Z(n26383) );
  BUF U4692 ( .I(n26288), .Z(n26382) );
  BUF U4693 ( .I(n26308), .Z(n26322) );
  BUF U4694 ( .I(n26308), .Z(n26321) );
  BUF U4695 ( .I(n26309), .Z(n26320) );
  BUF U4696 ( .I(n26310), .Z(n26316) );
  BUF U4697 ( .I(n26310), .Z(n26315) );
  BUF U4698 ( .I(n26309), .Z(n26319) );
  BUF U4699 ( .I(n26309), .Z(n26318) );
  BUF U4700 ( .I(n26310), .Z(n26317) );
  BUF U4701 ( .I(n26305), .Z(n26331) );
  BUF U4702 ( .I(n26305), .Z(n26330) );
  BUF U4703 ( .I(n26307), .Z(n26326) );
  BUF U4704 ( .I(n26307), .Z(n26325) );
  BUF U4705 ( .I(n26306), .Z(n26329) );
  BUF U4706 ( .I(n26306), .Z(n26328) );
  BUF U4707 ( .I(n26306), .Z(n26327) );
  BUF U4708 ( .I(n26302), .Z(n26341) );
  BUF U4709 ( .I(n26302), .Z(n26340) );
  BUF U4710 ( .I(n26304), .Z(n26335) );
  BUF U4711 ( .I(n26302), .Z(n26339) );
  BUF U4712 ( .I(n26303), .Z(n26338) );
  BUF U4713 ( .I(n26303), .Z(n26336) );
  BUF U4714 ( .I(n26303), .Z(n26337) );
  BUF U4715 ( .I(n26298), .Z(n26351) );
  BUF U4716 ( .I(n26299), .Z(n26350) );
  BUF U4717 ( .I(n26301), .Z(n26344) );
  BUF U4718 ( .I(n26300), .Z(n26345) );
  BUF U4719 ( .I(n26299), .Z(n26349) );
  BUF U4720 ( .I(n26299), .Z(n26348) );
  BUF U4721 ( .I(n26300), .Z(n26346) );
  BUF U4722 ( .I(n26300), .Z(n26347) );
  BUF U4723 ( .I(n26295), .Z(n26361) );
  BUF U4724 ( .I(n26295), .Z(n26360) );
  BUF U4725 ( .I(n26296), .Z(n26359) );
  BUF U4726 ( .I(n26297), .Z(n26354) );
  BUF U4727 ( .I(n26297), .Z(n26355) );
  BUF U4728 ( .I(n26296), .Z(n26358) );
  BUF U4729 ( .I(n26296), .Z(n26357) );
  BUF U4730 ( .I(n26297), .Z(n26356) );
  BUF U4731 ( .I(n26292), .Z(n26371) );
  BUF U4732 ( .I(n26292), .Z(n26370) );
  BUF U4733 ( .I(n26292), .Z(n26369) );
  BUF U4734 ( .I(n26294), .Z(n26365) );
  BUF U4735 ( .I(n26294), .Z(n26364) );
  BUF U4736 ( .I(n26293), .Z(n26368) );
  BUF U4737 ( .I(n26293), .Z(n26367) );
  BUF U4738 ( .I(n26293), .Z(n26366) );
  BUF U4739 ( .I(n26288), .Z(n26381) );
  BUF U4740 ( .I(n26289), .Z(n26380) );
  BUF U4741 ( .I(n26289), .Z(n26379) );
  BUF U4742 ( .I(n26290), .Z(n26375) );
  BUF U4743 ( .I(n26291), .Z(n26374) );
  BUF U4744 ( .I(n26289), .Z(n26378) );
  BUF U4745 ( .I(n26290), .Z(n26377) );
  BUF U4746 ( .I(n26290), .Z(n26376) );
  BUF U4747 ( .I(n26286), .Z(n26389) );
  BUF U4748 ( .I(n26287), .Z(n26385) );
  BUF U4749 ( .I(n26287), .Z(n26384) );
  BUF U4750 ( .I(n26286), .Z(n26388) );
  BUF U4751 ( .I(n26286), .Z(n26387) );
  BUF U4752 ( .I(n26287), .Z(n26386) );
  BUF U4753 ( .I(n26311), .Z(n26312) );
  BUF U4754 ( .I(n26408), .Z(n26546) );
  BUF U4755 ( .I(n26408), .Z(n26547) );
  BUF U4756 ( .I(n26413), .Z(n26532) );
  BUF U4757 ( .I(n26412), .Z(n26533) );
  BUF U4758 ( .I(n26412), .Z(n26534) );
  BUF U4759 ( .I(n26412), .Z(n26535) );
  BUF U4760 ( .I(n26402), .Z(n26419) );
  BUF U4761 ( .I(n26401), .Z(n26423) );
  BUF U4762 ( .I(n26398), .Z(n26432) );
  BUF U4763 ( .I(n26397), .Z(n26435) );
  BUF U4764 ( .I(n26395), .Z(n26441) );
  BUF U4765 ( .I(n26409), .Z(n26543) );
  BUF U4766 ( .I(n26408), .Z(n26545) );
  BUF U4767 ( .I(n26409), .Z(n26544) );
  BUF U4768 ( .I(n26411), .Z(n26538) );
  BUF U4769 ( .I(n26410), .Z(n26539) );
  BUF U4770 ( .I(n26410), .Z(n26540) );
  BUF U4771 ( .I(n26409), .Z(n26542) );
  BUF U4772 ( .I(n26410), .Z(n26541) );
  BUF U4773 ( .I(n26414), .Z(n26529) );
  BUF U4774 ( .I(n26413), .Z(n26530) );
  BUF U4775 ( .I(n26413), .Z(n26531) );
  BUF U4776 ( .I(n26415), .Z(n26525) );
  BUF U4777 ( .I(n26415), .Z(n26526) );
  BUF U4778 ( .I(n26414), .Z(n26527) );
  BUF U4779 ( .I(n26414), .Z(n26528) );
  INV U4780 ( .I(n1128), .ZN(n27374) );
  INV U4781 ( .I(n1128), .ZN(n27375) );
  INV U4782 ( .I(n1128), .ZN(n27376) );
  INV U4783 ( .I(n1258), .ZN(n27371) );
  INV U4784 ( .I(n1258), .ZN(n27372) );
  INV U4785 ( .I(n1258), .ZN(n27373) );
  INV U4786 ( .I(n1387), .ZN(n27368) );
  INV U4787 ( .I(n1387), .ZN(n27369) );
  INV U4788 ( .I(n1387), .ZN(n27370) );
  INV U4789 ( .I(n1645), .ZN(n27362) );
  INV U4790 ( .I(n1645), .ZN(n27363) );
  INV U4791 ( .I(n1645), .ZN(n27364) );
  INV U4792 ( .I(n1774), .ZN(n27359) );
  INV U4793 ( .I(n1774), .ZN(n27360) );
  INV U4794 ( .I(n1774), .ZN(n27361) );
  INV U4795 ( .I(n1903), .ZN(n27356) );
  INV U4796 ( .I(n1903), .ZN(n27357) );
  INV U4797 ( .I(n1903), .ZN(n27358) );
  INV U4798 ( .I(n2032), .ZN(n27353) );
  INV U4799 ( .I(n2032), .ZN(n27354) );
  INV U4800 ( .I(n2032), .ZN(n27355) );
  INV U4801 ( .I(n2161), .ZN(n27350) );
  INV U4802 ( .I(n2161), .ZN(n27351) );
  INV U4803 ( .I(n2161), .ZN(n27352) );
  INV U4804 ( .I(n2291), .ZN(n27347) );
  INV U4805 ( .I(n2291), .ZN(n27348) );
  INV U4806 ( .I(n2291), .ZN(n27349) );
  INV U4807 ( .I(n2420), .ZN(n27344) );
  INV U4808 ( .I(n2420), .ZN(n27345) );
  INV U4809 ( .I(n2420), .ZN(n27346) );
  NAND2 U4810 ( .A1(n27374), .A2(n5), .ZN(n2679) );
  NAND2 U4811 ( .A1(n27374), .A2(n6), .ZN(n2681) );
  NAND2 U4812 ( .A1(n27374), .A2(n7), .ZN(n2683) );
  NAND2 U4813 ( .A1(n27374), .A2(n8), .ZN(n2685) );
  NAND2 U4814 ( .A1(n27374), .A2(n9), .ZN(n2687) );
  NAND2 U4815 ( .A1(n27374), .A2(n42), .ZN(n2689) );
  NAND2 U4816 ( .A1(n27374), .A2(n45), .ZN(n2691) );
  NAND2 U4817 ( .A1(n27374), .A2(n48), .ZN(n2693) );
  NAND2 U4818 ( .A1(n27374), .A2(n51), .ZN(n2695) );
  NAND2 U4819 ( .A1(n27374), .A2(n54), .ZN(n2697) );
  NAND2 U4820 ( .A1(n27374), .A2(n57), .ZN(n2699) );
  NAND2 U4821 ( .A1(n27375), .A2(n60), .ZN(n2701) );
  NAND2 U4822 ( .A1(n27375), .A2(n63), .ZN(n2703) );
  NAND2 U4823 ( .A1(n27376), .A2(n66), .ZN(n2705) );
  NAND2 U4824 ( .A1(n27374), .A2(n69), .ZN(n2707) );
  NAND2 U4825 ( .A1(n27376), .A2(n72), .ZN(n2709) );
  NAND2 U4826 ( .A1(n27375), .A2(n75), .ZN(n2711) );
  NAND2 U4827 ( .A1(n27376), .A2(n78), .ZN(n2713) );
  NAND2 U4828 ( .A1(n27374), .A2(n81), .ZN(n2715) );
  NAND2 U4829 ( .A1(n27374), .A2(n84), .ZN(n2717) );
  NAND2 U4830 ( .A1(n27375), .A2(n87), .ZN(n2719) );
  NAND2 U4831 ( .A1(n27376), .A2(n90), .ZN(n2721) );
  NAND2 U4832 ( .A1(n27374), .A2(n93), .ZN(n2723) );
  NAND2 U4833 ( .A1(n27375), .A2(n96), .ZN(n2725) );
  NAND2 U4834 ( .A1(n27375), .A2(n99), .ZN(n2727) );
  NAND2 U4835 ( .A1(n27375), .A2(n102), .ZN(n2729) );
  NAND2 U4836 ( .A1(n27375), .A2(n105), .ZN(n2731) );
  NAND2 U4837 ( .A1(n27375), .A2(n108), .ZN(n2733) );
  NAND2 U4838 ( .A1(n27375), .A2(n111), .ZN(n2735) );
  NAND2 U4839 ( .A1(n27375), .A2(n114), .ZN(n2737) );
  NAND2 U4840 ( .A1(n27375), .A2(n117), .ZN(n2739) );
  NAND2 U4841 ( .A1(n27375), .A2(n120), .ZN(n2741) );
  NAND2 U4842 ( .A1(n27375), .A2(n123), .ZN(n2743) );
  NAND2 U4843 ( .A1(n27375), .A2(n126), .ZN(n2745) );
  NAND2 U4844 ( .A1(n27375), .A2(n129), .ZN(n2747) );
  NAND2 U4845 ( .A1(n27376), .A2(n132), .ZN(n2749) );
  NAND2 U4846 ( .A1(n27376), .A2(n135), .ZN(n2751) );
  NAND2 U4847 ( .A1(n27376), .A2(n138), .ZN(n2753) );
  NAND2 U4848 ( .A1(n27376), .A2(n141), .ZN(n2755) );
  NAND2 U4849 ( .A1(n27376), .A2(n144), .ZN(n2757) );
  NAND2 U4850 ( .A1(n27376), .A2(n147), .ZN(n2759) );
  NAND2 U4851 ( .A1(n27376), .A2(n150), .ZN(n2761) );
  NAND2 U4852 ( .A1(n27376), .A2(n153), .ZN(n2763) );
  NAND2 U4853 ( .A1(n27376), .A2(n156), .ZN(n2765) );
  NAND2 U4854 ( .A1(n27376), .A2(n159), .ZN(n2767) );
  NAND2 U4855 ( .A1(n27376), .A2(n162), .ZN(n2769) );
  NAND2 U4856 ( .A1(n27376), .A2(n165), .ZN(n2771) );
  NAND2 U4857 ( .A1(n27376), .A2(n10), .ZN(n2773) );
  NAND2 U4858 ( .A1(n27374), .A2(n11), .ZN(n2775) );
  NAND2 U4859 ( .A1(n27375), .A2(n12), .ZN(n2777) );
  NAND2 U4860 ( .A1(n27376), .A2(n24), .ZN(n2779) );
  NAND2 U4861 ( .A1(n27374), .A2(n27), .ZN(n2781) );
  NAND2 U4862 ( .A1(n27375), .A2(n30), .ZN(n2783) );
  NAND2 U4863 ( .A1(n27376), .A2(n33), .ZN(n2785) );
  NAND2 U4864 ( .A1(n27374), .A2(n36), .ZN(n2787) );
  NAND2 U4865 ( .A1(n27375), .A2(n39), .ZN(n2789) );
  NAND2 U4866 ( .A1(n27376), .A2(n168), .ZN(n2791) );
  NAND2 U4867 ( .A1(n27374), .A2(n171), .ZN(n2793) );
  NAND2 U4868 ( .A1(n27375), .A2(n174), .ZN(n2795) );
  NAND2 U4869 ( .A1(n27371), .A2(n5), .ZN(n2808) );
  NAND2 U4870 ( .A1(n27371), .A2(n6), .ZN(n2810) );
  NAND2 U4871 ( .A1(n27371), .A2(n7), .ZN(n2812) );
  NAND2 U4872 ( .A1(n27371), .A2(n8), .ZN(n2814) );
  NAND2 U4873 ( .A1(n27371), .A2(n9), .ZN(n2816) );
  NAND2 U4874 ( .A1(n27371), .A2(n42), .ZN(n2818) );
  NAND2 U4875 ( .A1(n27371), .A2(n45), .ZN(n2820) );
  NAND2 U4876 ( .A1(n27371), .A2(n48), .ZN(n2822) );
  NAND2 U4877 ( .A1(n27371), .A2(n51), .ZN(n2824) );
  NAND2 U4878 ( .A1(n27371), .A2(n54), .ZN(n2826) );
  NAND2 U4879 ( .A1(n27371), .A2(n57), .ZN(n2828) );
  NAND2 U4880 ( .A1(n27372), .A2(n60), .ZN(n2830) );
  NAND2 U4881 ( .A1(n27373), .A2(n63), .ZN(n2832) );
  NAND2 U4882 ( .A1(n27371), .A2(n66), .ZN(n2834) );
  NAND2 U4883 ( .A1(n27371), .A2(n69), .ZN(n2836) );
  NAND2 U4884 ( .A1(n27372), .A2(n72), .ZN(n2838) );
  NAND2 U4885 ( .A1(n27373), .A2(n75), .ZN(n2840) );
  NAND2 U4886 ( .A1(n27371), .A2(n78), .ZN(n2842) );
  NAND2 U4887 ( .A1(n27372), .A2(n81), .ZN(n2844) );
  NAND2 U4888 ( .A1(n27372), .A2(n84), .ZN(n2846) );
  NAND2 U4889 ( .A1(n27373), .A2(n87), .ZN(n2848) );
  NAND2 U4890 ( .A1(n27371), .A2(n90), .ZN(n2850) );
  NAND2 U4891 ( .A1(n27373), .A2(n93), .ZN(n2852) );
  NAND2 U4892 ( .A1(n27372), .A2(n96), .ZN(n2854) );
  NAND2 U4893 ( .A1(n27372), .A2(n99), .ZN(n2856) );
  NAND2 U4894 ( .A1(n27372), .A2(n102), .ZN(n2858) );
  NAND2 U4895 ( .A1(n27372), .A2(n105), .ZN(n2860) );
  NAND2 U4896 ( .A1(n27372), .A2(n108), .ZN(n2862) );
  NAND2 U4897 ( .A1(n27372), .A2(n111), .ZN(n2864) );
  NAND2 U4898 ( .A1(n27372), .A2(n114), .ZN(n2866) );
  NAND2 U4899 ( .A1(n27372), .A2(n117), .ZN(n2868) );
  NAND2 U4900 ( .A1(n27372), .A2(n120), .ZN(n2870) );
  NAND2 U4901 ( .A1(n27372), .A2(n123), .ZN(n2872) );
  NAND2 U4902 ( .A1(n27372), .A2(n126), .ZN(n2874) );
  NAND2 U4903 ( .A1(n27372), .A2(n129), .ZN(n2876) );
  NAND2 U4904 ( .A1(n27373), .A2(n132), .ZN(n2878) );
  NAND2 U4905 ( .A1(n27373), .A2(n135), .ZN(n2880) );
  NAND2 U4906 ( .A1(n27373), .A2(n138), .ZN(n2882) );
  NAND2 U4907 ( .A1(n27373), .A2(n141), .ZN(n2884) );
  NAND2 U4908 ( .A1(n27373), .A2(n144), .ZN(n2886) );
  NAND2 U4909 ( .A1(n27373), .A2(n147), .ZN(n2888) );
  NAND2 U4910 ( .A1(n27373), .A2(n150), .ZN(n2890) );
  NAND2 U4911 ( .A1(n27373), .A2(n153), .ZN(n2892) );
  NAND2 U4912 ( .A1(n27373), .A2(n156), .ZN(n2894) );
  NAND2 U4913 ( .A1(n27373), .A2(n159), .ZN(n2896) );
  NAND2 U4914 ( .A1(n27373), .A2(n162), .ZN(n2898) );
  NAND2 U4915 ( .A1(n27373), .A2(n165), .ZN(n2900) );
  NAND2 U4916 ( .A1(n27373), .A2(n10), .ZN(n2902) );
  NAND2 U4917 ( .A1(n27371), .A2(n11), .ZN(n2904) );
  NAND2 U4918 ( .A1(n27372), .A2(n12), .ZN(n2906) );
  NAND2 U4919 ( .A1(n27373), .A2(n24), .ZN(n2908) );
  NAND2 U4920 ( .A1(n27371), .A2(n27), .ZN(n2910) );
  NAND2 U4921 ( .A1(n27372), .A2(n30), .ZN(n2912) );
  NAND2 U4922 ( .A1(n27373), .A2(n33), .ZN(n2914) );
  NAND2 U4923 ( .A1(n27371), .A2(n36), .ZN(n2916) );
  NAND2 U4924 ( .A1(n27371), .A2(n39), .ZN(n2918) );
  NAND2 U4925 ( .A1(n27372), .A2(n168), .ZN(n2920) );
  NAND2 U4926 ( .A1(n27372), .A2(n171), .ZN(n2922) );
  NAND2 U4927 ( .A1(n27373), .A2(n174), .ZN(n2924) );
  NAND2 U4928 ( .A1(n27369), .A2(n5), .ZN(n2937) );
  NAND2 U4929 ( .A1(n27369), .A2(n6), .ZN(n2939) );
  NAND2 U4930 ( .A1(n27369), .A2(n7), .ZN(n2941) );
  NAND2 U4931 ( .A1(n27370), .A2(n8), .ZN(n2943) );
  NAND2 U4932 ( .A1(n27368), .A2(n9), .ZN(n2945) );
  NAND2 U4933 ( .A1(n27370), .A2(n42), .ZN(n2947) );
  NAND2 U4934 ( .A1(n27368), .A2(n45), .ZN(n2949) );
  NAND2 U4935 ( .A1(n27370), .A2(n48), .ZN(n2951) );
  NAND2 U4936 ( .A1(n27369), .A2(n51), .ZN(n2953) );
  NAND2 U4937 ( .A1(n27370), .A2(n54), .ZN(n2955) );
  NAND2 U4938 ( .A1(n27368), .A2(n57), .ZN(n2957) );
  NAND2 U4939 ( .A1(n27368), .A2(n60), .ZN(n2959) );
  NAND2 U4940 ( .A1(n27368), .A2(n63), .ZN(n2961) );
  NAND2 U4941 ( .A1(n27368), .A2(n66), .ZN(n2963) );
  NAND2 U4942 ( .A1(n27368), .A2(n69), .ZN(n2965) );
  NAND2 U4943 ( .A1(n27368), .A2(n72), .ZN(n2967) );
  NAND2 U4944 ( .A1(n27368), .A2(n75), .ZN(n2969) );
  NAND2 U4945 ( .A1(n27368), .A2(n78), .ZN(n2971) );
  NAND2 U4946 ( .A1(n27368), .A2(n81), .ZN(n2973) );
  NAND2 U4947 ( .A1(n27368), .A2(n84), .ZN(n2975) );
  NAND2 U4948 ( .A1(n27368), .A2(n87), .ZN(n2977) );
  NAND2 U4949 ( .A1(n27368), .A2(n90), .ZN(n2979) );
  NAND2 U4950 ( .A1(n27368), .A2(n93), .ZN(n2981) );
  NAND2 U4951 ( .A1(n27369), .A2(n96), .ZN(n2983) );
  NAND2 U4952 ( .A1(n27369), .A2(n99), .ZN(n2985) );
  NAND2 U4953 ( .A1(n27369), .A2(n102), .ZN(n2987) );
  NAND2 U4954 ( .A1(n27369), .A2(n105), .ZN(n2989) );
  NAND2 U4955 ( .A1(n27369), .A2(n108), .ZN(n2991) );
  NAND2 U4956 ( .A1(n27369), .A2(n111), .ZN(n2993) );
  NAND2 U4957 ( .A1(n27369), .A2(n114), .ZN(n2995) );
  NAND2 U4958 ( .A1(n27369), .A2(n117), .ZN(n2997) );
  NAND2 U4959 ( .A1(n27369), .A2(n120), .ZN(n2999) );
  NAND2 U4960 ( .A1(n27369), .A2(n123), .ZN(n3001) );
  NAND2 U4961 ( .A1(n27369), .A2(n126), .ZN(n3003) );
  NAND2 U4962 ( .A1(n27369), .A2(n129), .ZN(n3005) );
  NAND2 U4963 ( .A1(n27370), .A2(n132), .ZN(n3007) );
  NAND2 U4964 ( .A1(n27370), .A2(n135), .ZN(n3009) );
  NAND2 U4965 ( .A1(n27370), .A2(n138), .ZN(n3011) );
  NAND2 U4966 ( .A1(n27370), .A2(n141), .ZN(n3013) );
  NAND2 U4967 ( .A1(n27370), .A2(n144), .ZN(n3015) );
  NAND2 U4968 ( .A1(n27370), .A2(n147), .ZN(n3017) );
  NAND2 U4969 ( .A1(n27370), .A2(n150), .ZN(n3019) );
  NAND2 U4970 ( .A1(n27370), .A2(n153), .ZN(n3021) );
  NAND2 U4971 ( .A1(n27370), .A2(n156), .ZN(n3023) );
  NAND2 U4972 ( .A1(n27370), .A2(n159), .ZN(n3025) );
  NAND2 U4973 ( .A1(n27370), .A2(n162), .ZN(n3027) );
  NAND2 U4974 ( .A1(n27370), .A2(n165), .ZN(n3029) );
  NAND2 U4975 ( .A1(n27370), .A2(n10), .ZN(n3031) );
  NAND2 U4976 ( .A1(n27368), .A2(n11), .ZN(n3033) );
  NAND2 U4977 ( .A1(n27369), .A2(n12), .ZN(n3035) );
  NAND2 U4978 ( .A1(n27370), .A2(n24), .ZN(n3037) );
  NAND2 U4979 ( .A1(n27368), .A2(n27), .ZN(n3039) );
  NAND2 U4980 ( .A1(n27369), .A2(n30), .ZN(n3041) );
  NAND2 U4981 ( .A1(n27370), .A2(n33), .ZN(n3043) );
  NAND2 U4982 ( .A1(n27368), .A2(n36), .ZN(n3045) );
  NAND2 U4983 ( .A1(n27368), .A2(n39), .ZN(n3047) );
  NAND2 U4984 ( .A1(n27370), .A2(n168), .ZN(n3049) );
  NAND2 U4985 ( .A1(n27368), .A2(n171), .ZN(n3051) );
  NAND2 U4986 ( .A1(n27369), .A2(n174), .ZN(n3053) );
  NAND2 U4987 ( .A1(n27365), .A2(n5), .ZN(n3066) );
  NAND2 U4988 ( .A1(n27365), .A2(n6), .ZN(n3068) );
  NAND2 U4989 ( .A1(n27365), .A2(n7), .ZN(n3070) );
  NAND2 U4990 ( .A1(n27365), .A2(n8), .ZN(n3072) );
  NAND2 U4991 ( .A1(n27365), .A2(n9), .ZN(n3074) );
  NAND2 U4992 ( .A1(n27365), .A2(n42), .ZN(n3076) );
  NAND2 U4993 ( .A1(n27365), .A2(n45), .ZN(n3078) );
  NAND2 U4994 ( .A1(n27365), .A2(n48), .ZN(n3080) );
  NAND2 U4995 ( .A1(n27365), .A2(n51), .ZN(n3082) );
  NAND2 U4996 ( .A1(n27365), .A2(n54), .ZN(n3084) );
  NAND2 U4997 ( .A1(n27365), .A2(n57), .ZN(n3086) );
  NAND2 U4998 ( .A1(n27366), .A2(n60), .ZN(n3088) );
  NAND2 U4999 ( .A1(n27366), .A2(n63), .ZN(n3090) );
  NAND2 U5000 ( .A1(n27367), .A2(n66), .ZN(n3092) );
  NAND2 U5001 ( .A1(n27365), .A2(n69), .ZN(n3094) );
  NAND2 U5002 ( .A1(n27367), .A2(n72), .ZN(n3096) );
  NAND2 U5003 ( .A1(n27366), .A2(n75), .ZN(n3098) );
  NAND2 U5004 ( .A1(n27367), .A2(n78), .ZN(n3100) );
  NAND2 U5005 ( .A1(n27365), .A2(n81), .ZN(n3102) );
  NAND2 U5006 ( .A1(n27365), .A2(n84), .ZN(n3104) );
  NAND2 U5007 ( .A1(n27366), .A2(n87), .ZN(n3106) );
  NAND2 U5008 ( .A1(n27367), .A2(n90), .ZN(n3108) );
  NAND2 U5009 ( .A1(n27365), .A2(n93), .ZN(n3110) );
  NAND2 U5010 ( .A1(n27366), .A2(n96), .ZN(n3112) );
  NAND2 U5011 ( .A1(n27366), .A2(n99), .ZN(n3114) );
  NAND2 U5012 ( .A1(n27366), .A2(n102), .ZN(n3116) );
  NAND2 U5013 ( .A1(n27366), .A2(n105), .ZN(n3118) );
  NAND2 U5014 ( .A1(n27366), .A2(n108), .ZN(n3120) );
  NAND2 U5015 ( .A1(n27366), .A2(n111), .ZN(n3122) );
  NAND2 U5016 ( .A1(n27366), .A2(n114), .ZN(n3124) );
  NAND2 U5017 ( .A1(n27366), .A2(n117), .ZN(n3126) );
  NAND2 U5018 ( .A1(n27366), .A2(n120), .ZN(n3128) );
  NAND2 U5019 ( .A1(n27366), .A2(n123), .ZN(n3130) );
  NAND2 U5020 ( .A1(n27366), .A2(n126), .ZN(n3132) );
  NAND2 U5021 ( .A1(n27366), .A2(n129), .ZN(n3134) );
  NAND2 U5022 ( .A1(n27367), .A2(n132), .ZN(n3136) );
  NAND2 U5023 ( .A1(n27367), .A2(n135), .ZN(n3138) );
  NAND2 U5024 ( .A1(n27367), .A2(n138), .ZN(n3140) );
  NAND2 U5025 ( .A1(n27367), .A2(n141), .ZN(n3142) );
  NAND2 U5026 ( .A1(n27367), .A2(n144), .ZN(n3144) );
  NAND2 U5027 ( .A1(n27367), .A2(n147), .ZN(n3146) );
  NAND2 U5028 ( .A1(n27367), .A2(n150), .ZN(n3148) );
  NAND2 U5029 ( .A1(n27367), .A2(n153), .ZN(n3150) );
  NAND2 U5030 ( .A1(n27367), .A2(n156), .ZN(n3152) );
  NAND2 U5031 ( .A1(n27367), .A2(n159), .ZN(n3154) );
  NAND2 U5032 ( .A1(n27367), .A2(n162), .ZN(n3156) );
  NAND2 U5033 ( .A1(n27367), .A2(n165), .ZN(n3158) );
  NAND2 U5034 ( .A1(n27367), .A2(n10), .ZN(n3160) );
  NAND2 U5035 ( .A1(n27365), .A2(n11), .ZN(n3162) );
  NAND2 U5036 ( .A1(n27366), .A2(n12), .ZN(n3164) );
  NAND2 U5037 ( .A1(n27367), .A2(n24), .ZN(n3166) );
  NAND2 U5038 ( .A1(n27365), .A2(n27), .ZN(n3168) );
  NAND2 U5039 ( .A1(n27366), .A2(n30), .ZN(n3170) );
  NAND2 U5040 ( .A1(n27367), .A2(n33), .ZN(n3172) );
  NAND2 U5041 ( .A1(n27365), .A2(n36), .ZN(n3174) );
  NAND2 U5042 ( .A1(n27366), .A2(n39), .ZN(n3176) );
  NAND2 U5043 ( .A1(n27367), .A2(n168), .ZN(n3178) );
  NAND2 U5044 ( .A1(n27365), .A2(n171), .ZN(n3180) );
  NAND2 U5045 ( .A1(n27366), .A2(n174), .ZN(n3182) );
  NAND2 U5046 ( .A1(n27362), .A2(n5), .ZN(n3195) );
  NAND2 U5047 ( .A1(n27362), .A2(n6), .ZN(n3197) );
  NAND2 U5048 ( .A1(n27363), .A2(n7), .ZN(n3199) );
  NAND2 U5049 ( .A1(n27364), .A2(n8), .ZN(n3201) );
  NAND2 U5050 ( .A1(n27362), .A2(n9), .ZN(n3203) );
  NAND2 U5051 ( .A1(n27363), .A2(n42), .ZN(n3205) );
  NAND2 U5052 ( .A1(n27363), .A2(n45), .ZN(n3207) );
  NAND2 U5053 ( .A1(n27364), .A2(n48), .ZN(n3209) );
  NAND2 U5054 ( .A1(n27362), .A2(n51), .ZN(n3211) );
  NAND2 U5055 ( .A1(n27364), .A2(n54), .ZN(n3213) );
  NAND2 U5056 ( .A1(n27363), .A2(n57), .ZN(n3215) );
  NAND2 U5057 ( .A1(n27362), .A2(n60), .ZN(n3217) );
  NAND2 U5058 ( .A1(n27362), .A2(n63), .ZN(n3219) );
  NAND2 U5059 ( .A1(n27362), .A2(n66), .ZN(n3221) );
  NAND2 U5060 ( .A1(n27362), .A2(n69), .ZN(n3223) );
  NAND2 U5061 ( .A1(n27362), .A2(n72), .ZN(n3225) );
  NAND2 U5062 ( .A1(n27362), .A2(n75), .ZN(n3227) );
  NAND2 U5063 ( .A1(n27362), .A2(n78), .ZN(n3229) );
  NAND2 U5064 ( .A1(n27362), .A2(n81), .ZN(n3231) );
  NAND2 U5065 ( .A1(n27362), .A2(n84), .ZN(n3233) );
  NAND2 U5066 ( .A1(n27362), .A2(n87), .ZN(n3235) );
  NAND2 U5067 ( .A1(n27362), .A2(n90), .ZN(n3237) );
  NAND2 U5068 ( .A1(n27362), .A2(n93), .ZN(n3239) );
  NAND2 U5069 ( .A1(n27363), .A2(n96), .ZN(n3241) );
  NAND2 U5070 ( .A1(n27363), .A2(n99), .ZN(n3243) );
  NAND2 U5071 ( .A1(n27363), .A2(n102), .ZN(n3245) );
  NAND2 U5072 ( .A1(n27363), .A2(n105), .ZN(n3247) );
  NAND2 U5073 ( .A1(n27363), .A2(n108), .ZN(n3249) );
  NAND2 U5074 ( .A1(n27363), .A2(n111), .ZN(n3251) );
  NAND2 U5075 ( .A1(n27363), .A2(n114), .ZN(n3253) );
  NAND2 U5076 ( .A1(n27363), .A2(n117), .ZN(n3255) );
  NAND2 U5077 ( .A1(n27363), .A2(n120), .ZN(n3257) );
  NAND2 U5078 ( .A1(n27363), .A2(n123), .ZN(n3259) );
  NAND2 U5079 ( .A1(n27363), .A2(n126), .ZN(n3261) );
  NAND2 U5080 ( .A1(n27363), .A2(n129), .ZN(n3263) );
  NAND2 U5081 ( .A1(n27364), .A2(n132), .ZN(n3265) );
  NAND2 U5082 ( .A1(n27364), .A2(n135), .ZN(n3267) );
  NAND2 U5083 ( .A1(n27364), .A2(n138), .ZN(n3269) );
  NAND2 U5084 ( .A1(n27364), .A2(n141), .ZN(n3271) );
  NAND2 U5085 ( .A1(n27364), .A2(n144), .ZN(n3273) );
  NAND2 U5086 ( .A1(n27364), .A2(n147), .ZN(n3275) );
  NAND2 U5087 ( .A1(n27364), .A2(n150), .ZN(n3277) );
  NAND2 U5088 ( .A1(n27364), .A2(n153), .ZN(n3279) );
  NAND2 U5089 ( .A1(n27364), .A2(n156), .ZN(n3281) );
  NAND2 U5090 ( .A1(n27364), .A2(n159), .ZN(n3283) );
  NAND2 U5091 ( .A1(n27364), .A2(n162), .ZN(n3285) );
  NAND2 U5092 ( .A1(n27364), .A2(n165), .ZN(n3287) );
  NAND2 U5093 ( .A1(n27363), .A2(n10), .ZN(n3289) );
  NAND2 U5094 ( .A1(n27364), .A2(n11), .ZN(n3291) );
  NAND2 U5095 ( .A1(n27362), .A2(n12), .ZN(n3293) );
  NAND2 U5096 ( .A1(n27363), .A2(n24), .ZN(n3295) );
  NAND2 U5097 ( .A1(n27364), .A2(n27), .ZN(n3297) );
  NAND2 U5098 ( .A1(n27362), .A2(n30), .ZN(n3299) );
  NAND2 U5099 ( .A1(n27363), .A2(n33), .ZN(n3301) );
  NAND2 U5100 ( .A1(n27364), .A2(n36), .ZN(n3303) );
  NAND2 U5101 ( .A1(n27362), .A2(n39), .ZN(n3305) );
  NAND2 U5102 ( .A1(n27363), .A2(n168), .ZN(n3307) );
  NAND2 U5103 ( .A1(n27364), .A2(n171), .ZN(n3309) );
  NAND2 U5104 ( .A1(n27362), .A2(n174), .ZN(n3311) );
  NAND2 U5105 ( .A1(n27359), .A2(n5), .ZN(n3325) );
  NAND2 U5106 ( .A1(n27359), .A2(n6), .ZN(n3327) );
  NAND2 U5107 ( .A1(n27359), .A2(n7), .ZN(n3329) );
  NAND2 U5108 ( .A1(n27359), .A2(n8), .ZN(n3331) );
  NAND2 U5109 ( .A1(n27359), .A2(n9), .ZN(n3333) );
  NAND2 U5110 ( .A1(n27359), .A2(n42), .ZN(n3335) );
  NAND2 U5111 ( .A1(n27359), .A2(n45), .ZN(n3337) );
  NAND2 U5112 ( .A1(n27359), .A2(n48), .ZN(n3339) );
  NAND2 U5113 ( .A1(n27359), .A2(n51), .ZN(n3341) );
  NAND2 U5114 ( .A1(n27359), .A2(n54), .ZN(n3343) );
  NAND2 U5115 ( .A1(n27359), .A2(n57), .ZN(n3345) );
  NAND2 U5116 ( .A1(n27360), .A2(n60), .ZN(n3347) );
  NAND2 U5117 ( .A1(n27360), .A2(n63), .ZN(n3349) );
  NAND2 U5118 ( .A1(n27361), .A2(n66), .ZN(n3351) );
  NAND2 U5119 ( .A1(n27359), .A2(n69), .ZN(n3353) );
  NAND2 U5120 ( .A1(n27361), .A2(n72), .ZN(n3355) );
  NAND2 U5121 ( .A1(n27360), .A2(n75), .ZN(n3357) );
  NAND2 U5122 ( .A1(n27361), .A2(n78), .ZN(n3359) );
  NAND2 U5123 ( .A1(n27359), .A2(n81), .ZN(n3361) );
  NAND2 U5124 ( .A1(n27359), .A2(n84), .ZN(n3363) );
  NAND2 U5125 ( .A1(n27360), .A2(n87), .ZN(n3365) );
  NAND2 U5126 ( .A1(n27361), .A2(n90), .ZN(n3367) );
  NAND2 U5127 ( .A1(n27359), .A2(n93), .ZN(n3369) );
  NAND2 U5128 ( .A1(n27360), .A2(n96), .ZN(n3371) );
  NAND2 U5129 ( .A1(n27360), .A2(n99), .ZN(n3373) );
  NAND2 U5130 ( .A1(n27360), .A2(n102), .ZN(n3375) );
  NAND2 U5131 ( .A1(n27360), .A2(n105), .ZN(n3377) );
  NAND2 U5132 ( .A1(n27360), .A2(n108), .ZN(n3379) );
  NAND2 U5133 ( .A1(n27360), .A2(n111), .ZN(n3381) );
  NAND2 U5134 ( .A1(n27360), .A2(n114), .ZN(n3383) );
  NAND2 U5135 ( .A1(n27360), .A2(n117), .ZN(n3385) );
  NAND2 U5136 ( .A1(n27360), .A2(n120), .ZN(n3387) );
  NAND2 U5137 ( .A1(n27360), .A2(n123), .ZN(n3389) );
  NAND2 U5138 ( .A1(n27360), .A2(n126), .ZN(n3391) );
  NAND2 U5139 ( .A1(n27360), .A2(n129), .ZN(n3393) );
  NAND2 U5140 ( .A1(n27361), .A2(n132), .ZN(n3395) );
  NAND2 U5141 ( .A1(n27361), .A2(n135), .ZN(n3397) );
  NAND2 U5142 ( .A1(n27361), .A2(n138), .ZN(n3399) );
  NAND2 U5143 ( .A1(n27361), .A2(n141), .ZN(n3401) );
  NAND2 U5144 ( .A1(n27361), .A2(n144), .ZN(n3403) );
  NAND2 U5145 ( .A1(n27361), .A2(n147), .ZN(n3405) );
  NAND2 U5146 ( .A1(n27361), .A2(n150), .ZN(n3407) );
  NAND2 U5147 ( .A1(n27361), .A2(n153), .ZN(n3409) );
  NAND2 U5148 ( .A1(n27361), .A2(n156), .ZN(n3411) );
  NAND2 U5149 ( .A1(n27361), .A2(n159), .ZN(n3413) );
  NAND2 U5150 ( .A1(n27361), .A2(n162), .ZN(n3415) );
  NAND2 U5151 ( .A1(n27361), .A2(n165), .ZN(n3417) );
  NAND2 U5152 ( .A1(n27361), .A2(n10), .ZN(n3419) );
  NAND2 U5153 ( .A1(n27359), .A2(n11), .ZN(n3421) );
  NAND2 U5154 ( .A1(n27360), .A2(n12), .ZN(n3423) );
  NAND2 U5155 ( .A1(n27361), .A2(n24), .ZN(n3425) );
  NAND2 U5156 ( .A1(n27359), .A2(n27), .ZN(n3427) );
  NAND2 U5157 ( .A1(n27360), .A2(n30), .ZN(n3429) );
  NAND2 U5158 ( .A1(n27361), .A2(n33), .ZN(n3431) );
  NAND2 U5159 ( .A1(n27359), .A2(n36), .ZN(n3433) );
  NAND2 U5160 ( .A1(n27360), .A2(n39), .ZN(n3435) );
  NAND2 U5161 ( .A1(n27361), .A2(n168), .ZN(n3437) );
  NAND2 U5162 ( .A1(n27359), .A2(n171), .ZN(n3439) );
  NAND2 U5163 ( .A1(n27360), .A2(n174), .ZN(n3441) );
  NAND2 U5164 ( .A1(n27356), .A2(n5), .ZN(n3454) );
  NAND2 U5165 ( .A1(n27356), .A2(n6), .ZN(n3456) );
  NAND2 U5166 ( .A1(n27356), .A2(n7), .ZN(n3458) );
  NAND2 U5167 ( .A1(n27356), .A2(n8), .ZN(n3460) );
  NAND2 U5168 ( .A1(n27356), .A2(n9), .ZN(n3462) );
  NAND2 U5169 ( .A1(n27356), .A2(n42), .ZN(n3464) );
  NAND2 U5170 ( .A1(n27356), .A2(n45), .ZN(n3466) );
  NAND2 U5171 ( .A1(n27356), .A2(n48), .ZN(n3468) );
  NAND2 U5172 ( .A1(n27356), .A2(n51), .ZN(n3470) );
  NAND2 U5173 ( .A1(n27356), .A2(n54), .ZN(n3472) );
  NAND2 U5174 ( .A1(n27356), .A2(n57), .ZN(n3474) );
  NAND2 U5175 ( .A1(n27357), .A2(n60), .ZN(n3476) );
  NAND2 U5176 ( .A1(n27357), .A2(n63), .ZN(n3478) );
  NAND2 U5177 ( .A1(n27358), .A2(n66), .ZN(n3480) );
  NAND2 U5178 ( .A1(n27356), .A2(n69), .ZN(n3482) );
  NAND2 U5179 ( .A1(n27358), .A2(n72), .ZN(n3484) );
  NAND2 U5180 ( .A1(n27357), .A2(n75), .ZN(n3486) );
  NAND2 U5181 ( .A1(n27358), .A2(n78), .ZN(n3488) );
  NAND2 U5182 ( .A1(n27356), .A2(n81), .ZN(n3490) );
  NAND2 U5183 ( .A1(n27356), .A2(n84), .ZN(n3492) );
  NAND2 U5184 ( .A1(n27357), .A2(n87), .ZN(n3494) );
  NAND2 U5185 ( .A1(n27358), .A2(n90), .ZN(n3496) );
  NAND2 U5186 ( .A1(n27356), .A2(n93), .ZN(n3498) );
  NAND2 U5187 ( .A1(n27357), .A2(n96), .ZN(n3500) );
  NAND2 U5188 ( .A1(n27357), .A2(n99), .ZN(n3502) );
  NAND2 U5189 ( .A1(n27357), .A2(n102), .ZN(n3504) );
  NAND2 U5190 ( .A1(n27357), .A2(n105), .ZN(n3506) );
  NAND2 U5191 ( .A1(n27357), .A2(n108), .ZN(n3508) );
  NAND2 U5192 ( .A1(n27357), .A2(n111), .ZN(n3510) );
  NAND2 U5193 ( .A1(n27357), .A2(n114), .ZN(n3512) );
  NAND2 U5194 ( .A1(n27357), .A2(n117), .ZN(n3514) );
  NAND2 U5195 ( .A1(n27357), .A2(n120), .ZN(n3516) );
  NAND2 U5196 ( .A1(n27357), .A2(n123), .ZN(n3518) );
  NAND2 U5197 ( .A1(n27357), .A2(n126), .ZN(n3520) );
  NAND2 U5198 ( .A1(n27357), .A2(n129), .ZN(n3522) );
  NAND2 U5199 ( .A1(n27358), .A2(n132), .ZN(n3524) );
  NAND2 U5200 ( .A1(n27358), .A2(n135), .ZN(n3526) );
  NAND2 U5201 ( .A1(n27358), .A2(n138), .ZN(n3528) );
  NAND2 U5202 ( .A1(n27358), .A2(n141), .ZN(n3530) );
  NAND2 U5203 ( .A1(n27358), .A2(n144), .ZN(n3532) );
  NAND2 U5204 ( .A1(n27358), .A2(n147), .ZN(n3534) );
  NAND2 U5205 ( .A1(n27358), .A2(n150), .ZN(n3536) );
  NAND2 U5206 ( .A1(n27358), .A2(n153), .ZN(n3538) );
  NAND2 U5207 ( .A1(n27358), .A2(n156), .ZN(n3540) );
  NAND2 U5208 ( .A1(n27358), .A2(n159), .ZN(n3542) );
  NAND2 U5209 ( .A1(n27358), .A2(n162), .ZN(n3544) );
  NAND2 U5210 ( .A1(n27358), .A2(n165), .ZN(n3546) );
  NAND2 U5211 ( .A1(n27358), .A2(n10), .ZN(n3548) );
  NAND2 U5212 ( .A1(n27356), .A2(n11), .ZN(n3550) );
  NAND2 U5213 ( .A1(n27357), .A2(n12), .ZN(n3552) );
  NAND2 U5214 ( .A1(n27358), .A2(n24), .ZN(n3554) );
  NAND2 U5215 ( .A1(n27356), .A2(n27), .ZN(n3556) );
  NAND2 U5216 ( .A1(n27357), .A2(n30), .ZN(n3558) );
  NAND2 U5217 ( .A1(n27358), .A2(n33), .ZN(n3560) );
  NAND2 U5218 ( .A1(n27356), .A2(n36), .ZN(n3562) );
  NAND2 U5219 ( .A1(n27357), .A2(n39), .ZN(n3564) );
  NAND2 U5220 ( .A1(n27358), .A2(n168), .ZN(n3566) );
  NAND2 U5221 ( .A1(n27356), .A2(n171), .ZN(n3568) );
  NAND2 U5222 ( .A1(n27357), .A2(n174), .ZN(n3570) );
  NAND2 U5223 ( .A1(n27353), .A2(n5), .ZN(n3583) );
  NAND2 U5224 ( .A1(n27353), .A2(n6), .ZN(n3585) );
  NAND2 U5225 ( .A1(n27353), .A2(n7), .ZN(n3587) );
  NAND2 U5226 ( .A1(n27353), .A2(n8), .ZN(n3589) );
  NAND2 U5227 ( .A1(n27353), .A2(n9), .ZN(n3591) );
  NAND2 U5228 ( .A1(n27353), .A2(n42), .ZN(n3593) );
  NAND2 U5229 ( .A1(n27353), .A2(n45), .ZN(n3595) );
  NAND2 U5230 ( .A1(n27353), .A2(n48), .ZN(n3597) );
  NAND2 U5231 ( .A1(n27353), .A2(n51), .ZN(n3599) );
  NAND2 U5232 ( .A1(n27353), .A2(n54), .ZN(n3601) );
  NAND2 U5233 ( .A1(n27353), .A2(n57), .ZN(n3603) );
  NAND2 U5234 ( .A1(n27354), .A2(n60), .ZN(n3605) );
  NAND2 U5235 ( .A1(n27354), .A2(n63), .ZN(n3607) );
  NAND2 U5236 ( .A1(n27355), .A2(n66), .ZN(n3609) );
  NAND2 U5237 ( .A1(n27353), .A2(n69), .ZN(n3611) );
  NAND2 U5238 ( .A1(n27355), .A2(n72), .ZN(n3613) );
  NAND2 U5239 ( .A1(n27354), .A2(n75), .ZN(n3615) );
  NAND2 U5240 ( .A1(n27355), .A2(n78), .ZN(n3617) );
  NAND2 U5241 ( .A1(n27353), .A2(n81), .ZN(n3619) );
  NAND2 U5242 ( .A1(n27353), .A2(n84), .ZN(n3621) );
  NAND2 U5243 ( .A1(n27354), .A2(n87), .ZN(n3623) );
  NAND2 U5244 ( .A1(n27355), .A2(n90), .ZN(n3625) );
  NAND2 U5245 ( .A1(n27353), .A2(n93), .ZN(n3627) );
  NAND2 U5246 ( .A1(n27354), .A2(n96), .ZN(n3629) );
  NAND2 U5247 ( .A1(n27354), .A2(n99), .ZN(n3631) );
  NAND2 U5248 ( .A1(n27354), .A2(n102), .ZN(n3633) );
  NAND2 U5249 ( .A1(n27354), .A2(n105), .ZN(n3635) );
  NAND2 U5250 ( .A1(n27354), .A2(n108), .ZN(n3637) );
  NAND2 U5251 ( .A1(n27354), .A2(n111), .ZN(n3639) );
  NAND2 U5252 ( .A1(n27354), .A2(n114), .ZN(n3641) );
  NAND2 U5253 ( .A1(n27354), .A2(n117), .ZN(n3643) );
  NAND2 U5254 ( .A1(n27354), .A2(n120), .ZN(n3645) );
  NAND2 U5255 ( .A1(n27354), .A2(n123), .ZN(n3647) );
  NAND2 U5256 ( .A1(n27354), .A2(n126), .ZN(n3649) );
  NAND2 U5257 ( .A1(n27354), .A2(n129), .ZN(n3651) );
  NAND2 U5258 ( .A1(n27355), .A2(n132), .ZN(n3653) );
  NAND2 U5259 ( .A1(n27355), .A2(n135), .ZN(n3655) );
  NAND2 U5260 ( .A1(n27355), .A2(n138), .ZN(n3657) );
  NAND2 U5261 ( .A1(n27355), .A2(n141), .ZN(n3659) );
  NAND2 U5262 ( .A1(n27355), .A2(n144), .ZN(n3661) );
  NAND2 U5263 ( .A1(n27355), .A2(n147), .ZN(n3663) );
  NAND2 U5264 ( .A1(n27355), .A2(n150), .ZN(n3665) );
  NAND2 U5265 ( .A1(n27355), .A2(n153), .ZN(n3667) );
  NAND2 U5266 ( .A1(n27355), .A2(n156), .ZN(n3669) );
  NAND2 U5267 ( .A1(n27355), .A2(n159), .ZN(n3671) );
  NAND2 U5268 ( .A1(n27355), .A2(n162), .ZN(n3673) );
  NAND2 U5269 ( .A1(n27355), .A2(n165), .ZN(n3675) );
  NAND2 U5270 ( .A1(n27355), .A2(n10), .ZN(n3677) );
  NAND2 U5271 ( .A1(n27353), .A2(n11), .ZN(n3679) );
  NAND2 U5272 ( .A1(n27354), .A2(n12), .ZN(n3681) );
  NAND2 U5273 ( .A1(n27355), .A2(n24), .ZN(n3683) );
  NAND2 U5274 ( .A1(n27353), .A2(n27), .ZN(n3685) );
  NAND2 U5275 ( .A1(n27354), .A2(n30), .ZN(n3687) );
  NAND2 U5276 ( .A1(n27355), .A2(n33), .ZN(n3689) );
  NAND2 U5277 ( .A1(n27353), .A2(n36), .ZN(n3691) );
  NAND2 U5278 ( .A1(n27354), .A2(n39), .ZN(n3693) );
  NAND2 U5279 ( .A1(n27355), .A2(n168), .ZN(n3695) );
  NAND2 U5280 ( .A1(n27353), .A2(n171), .ZN(n3697) );
  NAND2 U5281 ( .A1(n27354), .A2(n174), .ZN(n3699) );
  NAND2 U5282 ( .A1(n27350), .A2(n5), .ZN(n3712) );
  NAND2 U5283 ( .A1(n27350), .A2(n6), .ZN(n3714) );
  NAND2 U5284 ( .A1(n27350), .A2(n7), .ZN(n3716) );
  NAND2 U5285 ( .A1(n27350), .A2(n8), .ZN(n3718) );
  NAND2 U5286 ( .A1(n27350), .A2(n9), .ZN(n3720) );
  NAND2 U5287 ( .A1(n27350), .A2(n42), .ZN(n3722) );
  NAND2 U5288 ( .A1(n27350), .A2(n45), .ZN(n3724) );
  NAND2 U5289 ( .A1(n27350), .A2(n48), .ZN(n3726) );
  NAND2 U5290 ( .A1(n27350), .A2(n51), .ZN(n3728) );
  NAND2 U5291 ( .A1(n27350), .A2(n54), .ZN(n3730) );
  NAND2 U5292 ( .A1(n27350), .A2(n57), .ZN(n3732) );
  NAND2 U5293 ( .A1(n27351), .A2(n60), .ZN(n3734) );
  NAND2 U5294 ( .A1(n27351), .A2(n63), .ZN(n3736) );
  NAND2 U5295 ( .A1(n27352), .A2(n66), .ZN(n3738) );
  NAND2 U5296 ( .A1(n27350), .A2(n69), .ZN(n3740) );
  NAND2 U5297 ( .A1(n27352), .A2(n72), .ZN(n3742) );
  NAND2 U5298 ( .A1(n27351), .A2(n75), .ZN(n3744) );
  NAND2 U5299 ( .A1(n27352), .A2(n78), .ZN(n3746) );
  NAND2 U5300 ( .A1(n27350), .A2(n81), .ZN(n3748) );
  NAND2 U5301 ( .A1(n27350), .A2(n84), .ZN(n3750) );
  NAND2 U5302 ( .A1(n27351), .A2(n87), .ZN(n3752) );
  NAND2 U5303 ( .A1(n27352), .A2(n90), .ZN(n3754) );
  NAND2 U5304 ( .A1(n27350), .A2(n93), .ZN(n3756) );
  NAND2 U5305 ( .A1(n27351), .A2(n96), .ZN(n3758) );
  NAND2 U5306 ( .A1(n27351), .A2(n99), .ZN(n3760) );
  NAND2 U5307 ( .A1(n27351), .A2(n102), .ZN(n3762) );
  NAND2 U5308 ( .A1(n27351), .A2(n105), .ZN(n3764) );
  NAND2 U5309 ( .A1(n27351), .A2(n108), .ZN(n3766) );
  NAND2 U5310 ( .A1(n27351), .A2(n111), .ZN(n3768) );
  NAND2 U5311 ( .A1(n27351), .A2(n114), .ZN(n3770) );
  NAND2 U5312 ( .A1(n27351), .A2(n117), .ZN(n3772) );
  NAND2 U5313 ( .A1(n27351), .A2(n120), .ZN(n3774) );
  NAND2 U5314 ( .A1(n27351), .A2(n123), .ZN(n3776) );
  NAND2 U5315 ( .A1(n27351), .A2(n126), .ZN(n3778) );
  NAND2 U5316 ( .A1(n27351), .A2(n129), .ZN(n3780) );
  NAND2 U5317 ( .A1(n27352), .A2(n132), .ZN(n3782) );
  NAND2 U5318 ( .A1(n27352), .A2(n135), .ZN(n3784) );
  NAND2 U5319 ( .A1(n27352), .A2(n138), .ZN(n3786) );
  NAND2 U5320 ( .A1(n27352), .A2(n141), .ZN(n3788) );
  NAND2 U5321 ( .A1(n27352), .A2(n144), .ZN(n3790) );
  NAND2 U5322 ( .A1(n27352), .A2(n147), .ZN(n3792) );
  NAND2 U5323 ( .A1(n27352), .A2(n150), .ZN(n3794) );
  NAND2 U5324 ( .A1(n27352), .A2(n153), .ZN(n3796) );
  NAND2 U5325 ( .A1(n27352), .A2(n156), .ZN(n3798) );
  NAND2 U5326 ( .A1(n27352), .A2(n159), .ZN(n3800) );
  NAND2 U5327 ( .A1(n27352), .A2(n162), .ZN(n3802) );
  NAND2 U5328 ( .A1(n27352), .A2(n165), .ZN(n3804) );
  NAND2 U5329 ( .A1(n27352), .A2(n10), .ZN(n3806) );
  NAND2 U5330 ( .A1(n27350), .A2(n11), .ZN(n3808) );
  NAND2 U5331 ( .A1(n27351), .A2(n12), .ZN(n3810) );
  NAND2 U5332 ( .A1(n27352), .A2(n24), .ZN(n3812) );
  NAND2 U5333 ( .A1(n27350), .A2(n27), .ZN(n3814) );
  NAND2 U5334 ( .A1(n27351), .A2(n30), .ZN(n3816) );
  NAND2 U5335 ( .A1(n27352), .A2(n33), .ZN(n3818) );
  NAND2 U5336 ( .A1(n27350), .A2(n36), .ZN(n3820) );
  NAND2 U5337 ( .A1(n27351), .A2(n39), .ZN(n3822) );
  NAND2 U5338 ( .A1(n27352), .A2(n168), .ZN(n3824) );
  NAND2 U5339 ( .A1(n27350), .A2(n171), .ZN(n3826) );
  NAND2 U5340 ( .A1(n27351), .A2(n174), .ZN(n3828) );
  NAND2 U5341 ( .A1(n27347), .A2(n5), .ZN(n3841) );
  NAND2 U5342 ( .A1(n27347), .A2(n6), .ZN(n3843) );
  NAND2 U5343 ( .A1(n27347), .A2(n7), .ZN(n3845) );
  NAND2 U5344 ( .A1(n27347), .A2(n8), .ZN(n3847) );
  NAND2 U5345 ( .A1(n27347), .A2(n9), .ZN(n3849) );
  NAND2 U5346 ( .A1(n27347), .A2(n42), .ZN(n3851) );
  NAND2 U5347 ( .A1(n27347), .A2(n45), .ZN(n3853) );
  NAND2 U5348 ( .A1(n27347), .A2(n48), .ZN(n3855) );
  NAND2 U5349 ( .A1(n27347), .A2(n51), .ZN(n3857) );
  NAND2 U5350 ( .A1(n27347), .A2(n54), .ZN(n3859) );
  NAND2 U5351 ( .A1(n27347), .A2(n57), .ZN(n3861) );
  NAND2 U5352 ( .A1(n27348), .A2(n60), .ZN(n3863) );
  NAND2 U5353 ( .A1(n27348), .A2(n63), .ZN(n3865) );
  NAND2 U5354 ( .A1(n27349), .A2(n66), .ZN(n3867) );
  NAND2 U5355 ( .A1(n27347), .A2(n69), .ZN(n3869) );
  NAND2 U5356 ( .A1(n27349), .A2(n72), .ZN(n3871) );
  NAND2 U5357 ( .A1(n27348), .A2(n75), .ZN(n3873) );
  NAND2 U5358 ( .A1(n27349), .A2(n78), .ZN(n3875) );
  NAND2 U5359 ( .A1(n27347), .A2(n81), .ZN(n3877) );
  NAND2 U5360 ( .A1(n27347), .A2(n84), .ZN(n3879) );
  NAND2 U5361 ( .A1(n27348), .A2(n87), .ZN(n3881) );
  NAND2 U5362 ( .A1(n27349), .A2(n90), .ZN(n3883) );
  NAND2 U5363 ( .A1(n27347), .A2(n93), .ZN(n3885) );
  NAND2 U5364 ( .A1(n27348), .A2(n96), .ZN(n3887) );
  NAND2 U5365 ( .A1(n27348), .A2(n99), .ZN(n3889) );
  NAND2 U5366 ( .A1(n27348), .A2(n102), .ZN(n3891) );
  NAND2 U5367 ( .A1(n27348), .A2(n105), .ZN(n3893) );
  NAND2 U5368 ( .A1(n27348), .A2(n108), .ZN(n3895) );
  NAND2 U5369 ( .A1(n27348), .A2(n111), .ZN(n3897) );
  NAND2 U5370 ( .A1(n27348), .A2(n114), .ZN(n3899) );
  NAND2 U5371 ( .A1(n27348), .A2(n117), .ZN(n3901) );
  NAND2 U5372 ( .A1(n27348), .A2(n120), .ZN(n3903) );
  NAND2 U5373 ( .A1(n27348), .A2(n123), .ZN(n3905) );
  NAND2 U5374 ( .A1(n27348), .A2(n126), .ZN(n3907) );
  NAND2 U5375 ( .A1(n27348), .A2(n129), .ZN(n3909) );
  NAND2 U5376 ( .A1(n27349), .A2(n132), .ZN(n3911) );
  NAND2 U5377 ( .A1(n27349), .A2(n135), .ZN(n3913) );
  NAND2 U5378 ( .A1(n27349), .A2(n138), .ZN(n3915) );
  NAND2 U5379 ( .A1(n27349), .A2(n141), .ZN(n3917) );
  NAND2 U5380 ( .A1(n27349), .A2(n144), .ZN(n3919) );
  NAND2 U5381 ( .A1(n27349), .A2(n147), .ZN(n3921) );
  NAND2 U5382 ( .A1(n27349), .A2(n150), .ZN(n3923) );
  NAND2 U5383 ( .A1(n27349), .A2(n153), .ZN(n3925) );
  NAND2 U5384 ( .A1(n27349), .A2(n156), .ZN(n3927) );
  NAND2 U5385 ( .A1(n27349), .A2(n159), .ZN(n3929) );
  NAND2 U5386 ( .A1(n27349), .A2(n162), .ZN(n3931) );
  NAND2 U5387 ( .A1(n27349), .A2(n165), .ZN(n3933) );
  NAND2 U5388 ( .A1(n27349), .A2(n10), .ZN(n3935) );
  NAND2 U5389 ( .A1(n27347), .A2(n11), .ZN(n3937) );
  NAND2 U5390 ( .A1(n27348), .A2(n12), .ZN(n3939) );
  NAND2 U5391 ( .A1(n27349), .A2(n24), .ZN(n3941) );
  NAND2 U5392 ( .A1(n27347), .A2(n27), .ZN(n3943) );
  NAND2 U5393 ( .A1(n27348), .A2(n30), .ZN(n3945) );
  NAND2 U5394 ( .A1(n27349), .A2(n33), .ZN(n3947) );
  NAND2 U5395 ( .A1(n27347), .A2(n36), .ZN(n3949) );
  NAND2 U5396 ( .A1(n27348), .A2(n39), .ZN(n3951) );
  NAND2 U5397 ( .A1(n27349), .A2(n168), .ZN(n3953) );
  NAND2 U5398 ( .A1(n27347), .A2(n171), .ZN(n3955) );
  NAND2 U5399 ( .A1(n27348), .A2(n174), .ZN(n3957) );
  NAND2 U5400 ( .A1(n27344), .A2(n5), .ZN(n3970) );
  NAND2 U5401 ( .A1(n27344), .A2(n6), .ZN(n3972) );
  NAND2 U5402 ( .A1(n27344), .A2(n7), .ZN(n3974) );
  NAND2 U5403 ( .A1(n27344), .A2(n8), .ZN(n3976) );
  NAND2 U5404 ( .A1(n27344), .A2(n9), .ZN(n3978) );
  NAND2 U5405 ( .A1(n27344), .A2(n42), .ZN(n3980) );
  NAND2 U5406 ( .A1(n27344), .A2(n45), .ZN(n3982) );
  NAND2 U5407 ( .A1(n27344), .A2(n48), .ZN(n3984) );
  NAND2 U5408 ( .A1(n27344), .A2(n51), .ZN(n3986) );
  NAND2 U5409 ( .A1(n27344), .A2(n54), .ZN(n3988) );
  NAND2 U5410 ( .A1(n27344), .A2(n57), .ZN(n3990) );
  NAND2 U5411 ( .A1(n27345), .A2(n60), .ZN(n3992) );
  NAND2 U5412 ( .A1(n27345), .A2(n63), .ZN(n3994) );
  NAND2 U5413 ( .A1(n27346), .A2(n66), .ZN(n3996) );
  NAND2 U5414 ( .A1(n27344), .A2(n69), .ZN(n3998) );
  NAND2 U5415 ( .A1(n27346), .A2(n72), .ZN(n4000) );
  NAND2 U5416 ( .A1(n27345), .A2(n75), .ZN(n4002) );
  NAND2 U5417 ( .A1(n27346), .A2(n78), .ZN(n4004) );
  NAND2 U5418 ( .A1(n27344), .A2(n81), .ZN(n4006) );
  NAND2 U5419 ( .A1(n27344), .A2(n84), .ZN(n4008) );
  NAND2 U5420 ( .A1(n27345), .A2(n87), .ZN(n4010) );
  NAND2 U5421 ( .A1(n27346), .A2(n90), .ZN(n4012) );
  NAND2 U5422 ( .A1(n27344), .A2(n93), .ZN(n4014) );
  NAND2 U5423 ( .A1(n27345), .A2(n96), .ZN(n4016) );
  NAND2 U5424 ( .A1(n27345), .A2(n99), .ZN(n4018) );
  NAND2 U5425 ( .A1(n27345), .A2(n102), .ZN(n4020) );
  NAND2 U5426 ( .A1(n27345), .A2(n105), .ZN(n4022) );
  NAND2 U5427 ( .A1(n27345), .A2(n108), .ZN(n4024) );
  NAND2 U5428 ( .A1(n27345), .A2(n111), .ZN(n4026) );
  NAND2 U5429 ( .A1(n27345), .A2(n114), .ZN(n4028) );
  NAND2 U5430 ( .A1(n27345), .A2(n117), .ZN(n4030) );
  NAND2 U5431 ( .A1(n27345), .A2(n120), .ZN(n4032) );
  NAND2 U5432 ( .A1(n27345), .A2(n123), .ZN(n4034) );
  NAND2 U5433 ( .A1(n27345), .A2(n126), .ZN(n4036) );
  NAND2 U5434 ( .A1(n27345), .A2(n129), .ZN(n4038) );
  NAND2 U5435 ( .A1(n27346), .A2(n132), .ZN(n4040) );
  NAND2 U5436 ( .A1(n27346), .A2(n135), .ZN(n4042) );
  NAND2 U5437 ( .A1(n27346), .A2(n138), .ZN(n4044) );
  NAND2 U5438 ( .A1(n27346), .A2(n141), .ZN(n4046) );
  NAND2 U5439 ( .A1(n27346), .A2(n144), .ZN(n4048) );
  NAND2 U5440 ( .A1(n27346), .A2(n147), .ZN(n4050) );
  NAND2 U5441 ( .A1(n27346), .A2(n150), .ZN(n4052) );
  NAND2 U5442 ( .A1(n27346), .A2(n153), .ZN(n4054) );
  NAND2 U5443 ( .A1(n27346), .A2(n156), .ZN(n4056) );
  NAND2 U5444 ( .A1(n27346), .A2(n159), .ZN(n4058) );
  NAND2 U5445 ( .A1(n27346), .A2(n162), .ZN(n4060) );
  NAND2 U5446 ( .A1(n27346), .A2(n165), .ZN(n4062) );
  NAND2 U5447 ( .A1(n27346), .A2(n10), .ZN(n4064) );
  NAND2 U5448 ( .A1(n27344), .A2(n11), .ZN(n4066) );
  NAND2 U5449 ( .A1(n27345), .A2(n12), .ZN(n4068) );
  NAND2 U5450 ( .A1(n27346), .A2(n24), .ZN(n4070) );
  NAND2 U5451 ( .A1(n27344), .A2(n27), .ZN(n4072) );
  NAND2 U5452 ( .A1(n27345), .A2(n30), .ZN(n4074) );
  NAND2 U5453 ( .A1(n27346), .A2(n33), .ZN(n4076) );
  NAND2 U5454 ( .A1(n27344), .A2(n36), .ZN(n4078) );
  NAND2 U5455 ( .A1(n27345), .A2(n39), .ZN(n4080) );
  NAND2 U5456 ( .A1(n27346), .A2(n168), .ZN(n4082) );
  NAND2 U5457 ( .A1(n27344), .A2(n171), .ZN(n4084) );
  NAND2 U5458 ( .A1(n27345), .A2(n174), .ZN(n4086) );
  NAND2 U5459 ( .A1(n27341), .A2(n5), .ZN(n4101) );
  NAND2 U5460 ( .A1(n27341), .A2(n6), .ZN(n4104) );
  NAND2 U5461 ( .A1(n27341), .A2(n7), .ZN(n4107) );
  NAND2 U5462 ( .A1(n27341), .A2(n8), .ZN(n4110) );
  NAND2 U5463 ( .A1(n27341), .A2(n9), .ZN(n4113) );
  NAND2 U5464 ( .A1(n27341), .A2(n42), .ZN(n4116) );
  NAND2 U5465 ( .A1(n27341), .A2(n45), .ZN(n4119) );
  NAND2 U5466 ( .A1(n27341), .A2(n48), .ZN(n4122) );
  NAND2 U5467 ( .A1(n27341), .A2(n51), .ZN(n4125) );
  NAND2 U5468 ( .A1(n27341), .A2(n54), .ZN(n4127) );
  NAND2 U5469 ( .A1(n27341), .A2(n57), .ZN(n4129) );
  NAND2 U5470 ( .A1(n27342), .A2(n60), .ZN(n4131) );
  NAND2 U5471 ( .A1(n27342), .A2(n63), .ZN(n4133) );
  NAND2 U5472 ( .A1(n27343), .A2(n66), .ZN(n4135) );
  NAND2 U5473 ( .A1(n27341), .A2(n69), .ZN(n4137) );
  NAND2 U5474 ( .A1(n27343), .A2(n72), .ZN(n4139) );
  NAND2 U5475 ( .A1(n27342), .A2(n75), .ZN(n4142) );
  NAND2 U5476 ( .A1(n27343), .A2(n78), .ZN(n4144) );
  NAND2 U5477 ( .A1(n27341), .A2(n81), .ZN(n4146) );
  NAND2 U5478 ( .A1(n27341), .A2(n84), .ZN(n4148) );
  NAND2 U5479 ( .A1(n27342), .A2(n87), .ZN(n4150) );
  NAND2 U5480 ( .A1(n27343), .A2(n90), .ZN(n4152) );
  NAND2 U5481 ( .A1(n27341), .A2(n93), .ZN(n4154) );
  NAND2 U5482 ( .A1(n27342), .A2(n96), .ZN(n4156) );
  NAND2 U5483 ( .A1(n27342), .A2(n99), .ZN(n4159) );
  NAND2 U5484 ( .A1(n27342), .A2(n102), .ZN(n4161) );
  NAND2 U5485 ( .A1(n27342), .A2(n105), .ZN(n4163) );
  NAND2 U5486 ( .A1(n27342), .A2(n108), .ZN(n4165) );
  NAND2 U5487 ( .A1(n27342), .A2(n111), .ZN(n4167) );
  NAND2 U5488 ( .A1(n27342), .A2(n114), .ZN(n4169) );
  NAND2 U5489 ( .A1(n27342), .A2(n117), .ZN(n4171) );
  NAND2 U5490 ( .A1(n27342), .A2(n120), .ZN(n4173) );
  NAND2 U5491 ( .A1(n27342), .A2(n123), .ZN(n4176) );
  NAND2 U5492 ( .A1(n27342), .A2(n126), .ZN(n4178) );
  NAND2 U5493 ( .A1(n27342), .A2(n129), .ZN(n4180) );
  NAND2 U5494 ( .A1(n27343), .A2(n132), .ZN(n4182) );
  NAND2 U5495 ( .A1(n27343), .A2(n135), .ZN(n4184) );
  NAND2 U5496 ( .A1(n27343), .A2(n138), .ZN(n4186) );
  NAND2 U5497 ( .A1(n27343), .A2(n141), .ZN(n4188) );
  NAND2 U5498 ( .A1(n27343), .A2(n144), .ZN(n4190) );
  NAND2 U5499 ( .A1(n27343), .A2(n147), .ZN(n4193) );
  NAND2 U5500 ( .A1(n27343), .A2(n150), .ZN(n4195) );
  NAND2 U5501 ( .A1(n27343), .A2(n153), .ZN(n4197) );
  NAND2 U5502 ( .A1(n27343), .A2(n156), .ZN(n4199) );
  NAND2 U5503 ( .A1(n27343), .A2(n159), .ZN(n4201) );
  NAND2 U5504 ( .A1(n27343), .A2(n162), .ZN(n4203) );
  NAND2 U5505 ( .A1(n27343), .A2(n165), .ZN(n4205) );
  NAND2 U5506 ( .A1(n27343), .A2(n10), .ZN(n4207) );
  NAND2 U5507 ( .A1(n27341), .A2(n11), .ZN(n4210) );
  NAND2 U5508 ( .A1(n27342), .A2(n12), .ZN(n4212) );
  NAND2 U5509 ( .A1(n27343), .A2(n24), .ZN(n4214) );
  NAND2 U5510 ( .A1(n27341), .A2(n27), .ZN(n4216) );
  NAND2 U5511 ( .A1(n27342), .A2(n30), .ZN(n4218) );
  NAND2 U5512 ( .A1(n27343), .A2(n33), .ZN(n4220) );
  NAND2 U5513 ( .A1(n27341), .A2(n36), .ZN(n4222) );
  NAND2 U5514 ( .A1(n27342), .A2(n39), .ZN(n4224) );
  NAND2 U5515 ( .A1(n27343), .A2(n168), .ZN(n4227) );
  NAND2 U5516 ( .A1(n27341), .A2(n171), .ZN(n4229) );
  NAND2 U5517 ( .A1(n27342), .A2(n174), .ZN(n4231) );
  NAND2 U5518 ( .A1(n27375), .A2(n1), .ZN(n2797) );
  NAND2 U5519 ( .A1(n27375), .A2(n2), .ZN(n2799) );
  NAND2 U5520 ( .A1(n27376), .A2(n3), .ZN(n2801) );
  NAND2 U5521 ( .A1(n27374), .A2(n4), .ZN(n2803) );
  NAND2 U5522 ( .A1(n27371), .A2(n1), .ZN(n2926) );
  NAND2 U5523 ( .A1(n27372), .A2(n2), .ZN(n2928) );
  NAND2 U5524 ( .A1(n27373), .A2(n3), .ZN(n2930) );
  NAND2 U5525 ( .A1(n27371), .A2(n4), .ZN(n2932) );
  NAND2 U5526 ( .A1(n27370), .A2(n1), .ZN(n3055) );
  NAND2 U5527 ( .A1(n27369), .A2(n2), .ZN(n3057) );
  NAND2 U5528 ( .A1(n27370), .A2(n3), .ZN(n3059) );
  NAND2 U5529 ( .A1(n27368), .A2(n4), .ZN(n3061) );
  NAND2 U5530 ( .A1(n27366), .A2(n1), .ZN(n3184) );
  NAND2 U5531 ( .A1(n27366), .A2(n2), .ZN(n3186) );
  NAND2 U5532 ( .A1(n27367), .A2(n3), .ZN(n3188) );
  NAND2 U5533 ( .A1(n27363), .A2(n1), .ZN(n3313) );
  NAND2 U5534 ( .A1(n27363), .A2(n2), .ZN(n3315) );
  NAND2 U5535 ( .A1(n27364), .A2(n3), .ZN(n3317) );
  NAND2 U5536 ( .A1(n27362), .A2(n4), .ZN(n3319) );
  NAND2 U5537 ( .A1(n27360), .A2(n1), .ZN(n3443) );
  NAND2 U5538 ( .A1(n27360), .A2(n2), .ZN(n3445) );
  NAND2 U5539 ( .A1(n27361), .A2(n3), .ZN(n3447) );
  NAND2 U5540 ( .A1(n27359), .A2(n4), .ZN(n3449) );
  NAND2 U5541 ( .A1(n27357), .A2(n1), .ZN(n3572) );
  NAND2 U5542 ( .A1(n27357), .A2(n2), .ZN(n3574) );
  NAND2 U5543 ( .A1(n27358), .A2(n3), .ZN(n3576) );
  NAND2 U5544 ( .A1(n27356), .A2(n4), .ZN(n3578) );
  NAND2 U5545 ( .A1(n27354), .A2(n1), .ZN(n3701) );
  NAND2 U5546 ( .A1(n27354), .A2(n2), .ZN(n3703) );
  NAND2 U5547 ( .A1(n27355), .A2(n3), .ZN(n3705) );
  NAND2 U5548 ( .A1(n27353), .A2(n4), .ZN(n3707) );
  NAND2 U5549 ( .A1(n27351), .A2(n1), .ZN(n3830) );
  NAND2 U5550 ( .A1(n27351), .A2(n2), .ZN(n3832) );
  NAND2 U5551 ( .A1(n27352), .A2(n3), .ZN(n3834) );
  NAND2 U5552 ( .A1(n27350), .A2(n4), .ZN(n3836) );
  NAND2 U5553 ( .A1(n27348), .A2(n1), .ZN(n3959) );
  NAND2 U5554 ( .A1(n27348), .A2(n2), .ZN(n3961) );
  NAND2 U5555 ( .A1(n27349), .A2(n3), .ZN(n3963) );
  NAND2 U5556 ( .A1(n27347), .A2(n4), .ZN(n3965) );
  NAND2 U5557 ( .A1(n27345), .A2(n1), .ZN(n4088) );
  NAND2 U5558 ( .A1(n27345), .A2(n2), .ZN(n4090) );
  NAND2 U5559 ( .A1(n27346), .A2(n3), .ZN(n4092) );
  NAND2 U5560 ( .A1(n27344), .A2(n4), .ZN(n4094) );
  NAND2 U5561 ( .A1(n27342), .A2(n1), .ZN(n4233) );
  NAND2 U5562 ( .A1(n27342), .A2(n2), .ZN(n4235) );
  NAND2 U5563 ( .A1(n27343), .A2(n3), .ZN(n4237) );
  NAND2 U5564 ( .A1(n27365), .A2(n4), .ZN(n3190) );
  NAND2 U5565 ( .A1(n27341), .A2(n4), .ZN(n4239) );
  BUF U5566 ( .I(n29571), .Z(n29494) );
  BUF U5567 ( .I(n29572), .Z(n29571) );
  BUF U5568 ( .I(n29298), .Z(n29088) );
  BUF U5569 ( .I(n29063), .Z(n28853) );
  BUF U5570 ( .I(n28828), .Z(n28618) );
  BUF U5571 ( .I(n28593), .Z(n28383) );
  BUF U5572 ( .I(n28358), .Z(n28148) );
  BUF U5573 ( .I(n28123), .Z(n27913) );
  BUF U5574 ( .I(n27888), .Z(n27678) );
  BUF U5575 ( .I(n27653), .Z(n27443) );
  BUF U5576 ( .I(n29298), .Z(n29089) );
  BUF U5577 ( .I(n29063), .Z(n28854) );
  BUF U5578 ( .I(n28828), .Z(n28619) );
  BUF U5579 ( .I(n28593), .Z(n28384) );
  BUF U5580 ( .I(n28358), .Z(n28149) );
  BUF U5581 ( .I(n28123), .Z(n27914) );
  BUF U5582 ( .I(n27888), .Z(n27679) );
  BUF U5583 ( .I(n27653), .Z(n27444) );
  BUF U5584 ( .I(n29297), .Z(n29090) );
  BUF U5585 ( .I(n29062), .Z(n28855) );
  BUF U5586 ( .I(n28827), .Z(n28620) );
  BUF U5587 ( .I(n28592), .Z(n28385) );
  BUF U5588 ( .I(n28357), .Z(n28150) );
  BUF U5589 ( .I(n28122), .Z(n27915) );
  BUF U5590 ( .I(n27887), .Z(n27680) );
  BUF U5591 ( .I(n27652), .Z(n27445) );
  BUF U5592 ( .I(n29297), .Z(n29091) );
  BUF U5593 ( .I(n29062), .Z(n28856) );
  BUF U5594 ( .I(n28827), .Z(n28621) );
  BUF U5595 ( .I(n28592), .Z(n28386) );
  BUF U5596 ( .I(n28357), .Z(n28151) );
  BUF U5597 ( .I(n28122), .Z(n27916) );
  BUF U5598 ( .I(n27887), .Z(n27681) );
  BUF U5599 ( .I(n27652), .Z(n27446) );
  BUF U5600 ( .I(n29297), .Z(n29092) );
  BUF U5601 ( .I(n29062), .Z(n28857) );
  BUF U5602 ( .I(n28827), .Z(n28622) );
  BUF U5603 ( .I(n28592), .Z(n28387) );
  BUF U5604 ( .I(n28357), .Z(n28152) );
  BUF U5605 ( .I(n28122), .Z(n27917) );
  BUF U5606 ( .I(n27887), .Z(n27682) );
  BUF U5607 ( .I(n27652), .Z(n27447) );
  BUF U5608 ( .I(n29296), .Z(n29093) );
  BUF U5609 ( .I(n29061), .Z(n28858) );
  BUF U5610 ( .I(n28826), .Z(n28623) );
  BUF U5611 ( .I(n28591), .Z(n28388) );
  BUF U5612 ( .I(n28356), .Z(n28153) );
  BUF U5613 ( .I(n28121), .Z(n27918) );
  BUF U5614 ( .I(n27886), .Z(n27683) );
  BUF U5615 ( .I(n27651), .Z(n27448) );
  BUF U5616 ( .I(n29296), .Z(n29094) );
  BUF U5617 ( .I(n29061), .Z(n28859) );
  BUF U5618 ( .I(n28826), .Z(n28624) );
  BUF U5619 ( .I(n28591), .Z(n28389) );
  BUF U5620 ( .I(n28356), .Z(n28154) );
  BUF U5621 ( .I(n28121), .Z(n27919) );
  BUF U5622 ( .I(n27886), .Z(n27684) );
  BUF U5623 ( .I(n27651), .Z(n27449) );
  BUF U5624 ( .I(n29296), .Z(n29095) );
  BUF U5625 ( .I(n29061), .Z(n28860) );
  BUF U5626 ( .I(n28826), .Z(n28625) );
  BUF U5627 ( .I(n28591), .Z(n28390) );
  BUF U5628 ( .I(n28356), .Z(n28155) );
  BUF U5629 ( .I(n28121), .Z(n27920) );
  BUF U5630 ( .I(n27886), .Z(n27685) );
  BUF U5631 ( .I(n27651), .Z(n27450) );
  BUF U5632 ( .I(n29295), .Z(n29096) );
  BUF U5633 ( .I(n29060), .Z(n28861) );
  BUF U5634 ( .I(n28825), .Z(n28626) );
  BUF U5635 ( .I(n28590), .Z(n28391) );
  BUF U5636 ( .I(n28355), .Z(n28156) );
  BUF U5637 ( .I(n28120), .Z(n27921) );
  BUF U5638 ( .I(n27885), .Z(n27686) );
  BUF U5639 ( .I(n27650), .Z(n27451) );
  BUF U5640 ( .I(n29295), .Z(n29097) );
  BUF U5641 ( .I(n29060), .Z(n28862) );
  BUF U5642 ( .I(n28825), .Z(n28627) );
  BUF U5643 ( .I(n28590), .Z(n28392) );
  BUF U5644 ( .I(n28355), .Z(n28157) );
  BUF U5645 ( .I(n28120), .Z(n27922) );
  BUF U5646 ( .I(n27885), .Z(n27687) );
  BUF U5647 ( .I(n27650), .Z(n27452) );
  BUF U5648 ( .I(n29295), .Z(n29098) );
  BUF U5649 ( .I(n29060), .Z(n28863) );
  BUF U5650 ( .I(n28825), .Z(n28628) );
  BUF U5651 ( .I(n28590), .Z(n28393) );
  BUF U5652 ( .I(n28355), .Z(n28158) );
  BUF U5653 ( .I(n28120), .Z(n27923) );
  BUF U5654 ( .I(n27885), .Z(n27688) );
  BUF U5655 ( .I(n27650), .Z(n27453) );
  BUF U5656 ( .I(n29294), .Z(n29099) );
  BUF U5657 ( .I(n29059), .Z(n28864) );
  BUF U5658 ( .I(n28824), .Z(n28629) );
  BUF U5659 ( .I(n28589), .Z(n28394) );
  BUF U5660 ( .I(n28354), .Z(n28159) );
  BUF U5661 ( .I(n28119), .Z(n27924) );
  BUF U5662 ( .I(n27884), .Z(n27689) );
  BUF U5663 ( .I(n27649), .Z(n27454) );
  BUF U5664 ( .I(n29294), .Z(n29100) );
  BUF U5665 ( .I(n29059), .Z(n28865) );
  BUF U5666 ( .I(n28824), .Z(n28630) );
  BUF U5667 ( .I(n28589), .Z(n28395) );
  BUF U5668 ( .I(n28354), .Z(n28160) );
  BUF U5669 ( .I(n28119), .Z(n27925) );
  BUF U5670 ( .I(n27884), .Z(n27690) );
  BUF U5671 ( .I(n27649), .Z(n27455) );
  BUF U5672 ( .I(n29294), .Z(n29101) );
  BUF U5673 ( .I(n29059), .Z(n28866) );
  BUF U5674 ( .I(n28824), .Z(n28631) );
  BUF U5675 ( .I(n28589), .Z(n28396) );
  BUF U5676 ( .I(n28354), .Z(n28161) );
  BUF U5677 ( .I(n28119), .Z(n27926) );
  BUF U5678 ( .I(n27884), .Z(n27691) );
  BUF U5679 ( .I(n27649), .Z(n27456) );
  BUF U5680 ( .I(n29293), .Z(n29102) );
  BUF U5681 ( .I(n29058), .Z(n28867) );
  BUF U5682 ( .I(n28823), .Z(n28632) );
  BUF U5683 ( .I(n28588), .Z(n28397) );
  BUF U5684 ( .I(n28353), .Z(n28162) );
  BUF U5685 ( .I(n28118), .Z(n27927) );
  BUF U5686 ( .I(n27883), .Z(n27692) );
  BUF U5687 ( .I(n27648), .Z(n27457) );
  BUF U5688 ( .I(n29293), .Z(n29103) );
  BUF U5689 ( .I(n29058), .Z(n28868) );
  BUF U5690 ( .I(n28823), .Z(n28633) );
  BUF U5691 ( .I(n28588), .Z(n28398) );
  BUF U5692 ( .I(n28353), .Z(n28163) );
  BUF U5693 ( .I(n28118), .Z(n27928) );
  BUF U5694 ( .I(n27883), .Z(n27693) );
  BUF U5695 ( .I(n27648), .Z(n27458) );
  BUF U5696 ( .I(n29293), .Z(n29104) );
  BUF U5697 ( .I(n29058), .Z(n28869) );
  BUF U5698 ( .I(n28823), .Z(n28634) );
  BUF U5699 ( .I(n28588), .Z(n28399) );
  BUF U5700 ( .I(n28353), .Z(n28164) );
  BUF U5701 ( .I(n28118), .Z(n27929) );
  BUF U5702 ( .I(n27883), .Z(n27694) );
  BUF U5703 ( .I(n27648), .Z(n27459) );
  BUF U5704 ( .I(n29292), .Z(n29105) );
  BUF U5705 ( .I(n29057), .Z(n28870) );
  BUF U5706 ( .I(n28822), .Z(n28635) );
  BUF U5707 ( .I(n28587), .Z(n28400) );
  BUF U5708 ( .I(n28352), .Z(n28165) );
  BUF U5709 ( .I(n28117), .Z(n27930) );
  BUF U5710 ( .I(n27882), .Z(n27695) );
  BUF U5711 ( .I(n27647), .Z(n27460) );
  BUF U5712 ( .I(n29292), .Z(n29106) );
  BUF U5713 ( .I(n29057), .Z(n28871) );
  BUF U5714 ( .I(n28822), .Z(n28636) );
  BUF U5715 ( .I(n28587), .Z(n28401) );
  BUF U5716 ( .I(n28352), .Z(n28166) );
  BUF U5717 ( .I(n28117), .Z(n27931) );
  BUF U5718 ( .I(n27882), .Z(n27696) );
  BUF U5719 ( .I(n27647), .Z(n27461) );
  BUF U5720 ( .I(n29292), .Z(n29107) );
  BUF U5721 ( .I(n29057), .Z(n28872) );
  BUF U5722 ( .I(n28822), .Z(n28637) );
  BUF U5723 ( .I(n28587), .Z(n28402) );
  BUF U5724 ( .I(n28352), .Z(n28167) );
  BUF U5725 ( .I(n28117), .Z(n27932) );
  BUF U5726 ( .I(n27882), .Z(n27697) );
  BUF U5727 ( .I(n27647), .Z(n27462) );
  BUF U5728 ( .I(n29291), .Z(n29108) );
  BUF U5729 ( .I(n29056), .Z(n28873) );
  BUF U5730 ( .I(n28821), .Z(n28638) );
  BUF U5731 ( .I(n28586), .Z(n28403) );
  BUF U5732 ( .I(n28351), .Z(n28168) );
  BUF U5733 ( .I(n28116), .Z(n27933) );
  BUF U5734 ( .I(n27881), .Z(n27698) );
  BUF U5735 ( .I(n27646), .Z(n27463) );
  BUF U5736 ( .I(n29291), .Z(n29109) );
  BUF U5737 ( .I(n29056), .Z(n28874) );
  BUF U5738 ( .I(n28821), .Z(n28639) );
  BUF U5739 ( .I(n28586), .Z(n28404) );
  BUF U5740 ( .I(n28351), .Z(n28169) );
  BUF U5741 ( .I(n28116), .Z(n27934) );
  BUF U5742 ( .I(n27881), .Z(n27699) );
  BUF U5743 ( .I(n27646), .Z(n27464) );
  BUF U5744 ( .I(n29291), .Z(n29110) );
  BUF U5745 ( .I(n29056), .Z(n28875) );
  BUF U5746 ( .I(n28821), .Z(n28640) );
  BUF U5747 ( .I(n28586), .Z(n28405) );
  BUF U5748 ( .I(n28351), .Z(n28170) );
  BUF U5749 ( .I(n28116), .Z(n27935) );
  BUF U5750 ( .I(n27881), .Z(n27700) );
  BUF U5751 ( .I(n27646), .Z(n27465) );
  BUF U5752 ( .I(n29290), .Z(n29111) );
  BUF U5753 ( .I(n29055), .Z(n28876) );
  BUF U5754 ( .I(n28820), .Z(n28641) );
  BUF U5755 ( .I(n28585), .Z(n28406) );
  BUF U5756 ( .I(n28350), .Z(n28171) );
  BUF U5757 ( .I(n28115), .Z(n27936) );
  BUF U5758 ( .I(n27880), .Z(n27701) );
  BUF U5759 ( .I(n27645), .Z(n27466) );
  BUF U5760 ( .I(n29290), .Z(n29112) );
  BUF U5761 ( .I(n29055), .Z(n28877) );
  BUF U5762 ( .I(n28820), .Z(n28642) );
  BUF U5763 ( .I(n28585), .Z(n28407) );
  BUF U5764 ( .I(n28350), .Z(n28172) );
  BUF U5765 ( .I(n28115), .Z(n27937) );
  BUF U5766 ( .I(n27880), .Z(n27702) );
  BUF U5767 ( .I(n27645), .Z(n27467) );
  BUF U5768 ( .I(n29290), .Z(n29113) );
  BUF U5769 ( .I(n29055), .Z(n28878) );
  BUF U5770 ( .I(n28820), .Z(n28643) );
  BUF U5771 ( .I(n28585), .Z(n28408) );
  BUF U5772 ( .I(n28350), .Z(n28173) );
  BUF U5773 ( .I(n28115), .Z(n27938) );
  BUF U5774 ( .I(n27880), .Z(n27703) );
  BUF U5775 ( .I(n27645), .Z(n27468) );
  BUF U5776 ( .I(n29289), .Z(n29114) );
  BUF U5777 ( .I(n29054), .Z(n28879) );
  BUF U5778 ( .I(n28819), .Z(n28644) );
  BUF U5779 ( .I(n28584), .Z(n28409) );
  BUF U5780 ( .I(n28349), .Z(n28174) );
  BUF U5781 ( .I(n28114), .Z(n27939) );
  BUF U5782 ( .I(n27879), .Z(n27704) );
  BUF U5783 ( .I(n27644), .Z(n27469) );
  BUF U5784 ( .I(n29289), .Z(n29115) );
  BUF U5785 ( .I(n29054), .Z(n28880) );
  BUF U5786 ( .I(n28819), .Z(n28645) );
  BUF U5787 ( .I(n28584), .Z(n28410) );
  BUF U5788 ( .I(n28349), .Z(n28175) );
  BUF U5789 ( .I(n28114), .Z(n27940) );
  BUF U5790 ( .I(n27879), .Z(n27705) );
  BUF U5791 ( .I(n27644), .Z(n27470) );
  BUF U5792 ( .I(n29289), .Z(n29116) );
  BUF U5793 ( .I(n29054), .Z(n28881) );
  BUF U5794 ( .I(n28819), .Z(n28646) );
  BUF U5795 ( .I(n28584), .Z(n28411) );
  BUF U5796 ( .I(n28349), .Z(n28176) );
  BUF U5797 ( .I(n28114), .Z(n27941) );
  BUF U5798 ( .I(n27879), .Z(n27706) );
  BUF U5799 ( .I(n27644), .Z(n27471) );
  BUF U5800 ( .I(n29288), .Z(n29117) );
  BUF U5801 ( .I(n29053), .Z(n28882) );
  BUF U5802 ( .I(n28818), .Z(n28647) );
  BUF U5803 ( .I(n28583), .Z(n28412) );
  BUF U5804 ( .I(n28348), .Z(n28177) );
  BUF U5805 ( .I(n28113), .Z(n27942) );
  BUF U5806 ( .I(n27878), .Z(n27707) );
  BUF U5807 ( .I(n27643), .Z(n27472) );
  BUF U5808 ( .I(n29288), .Z(n29118) );
  BUF U5809 ( .I(n29053), .Z(n28883) );
  BUF U5810 ( .I(n28818), .Z(n28648) );
  BUF U5811 ( .I(n28583), .Z(n28413) );
  BUF U5812 ( .I(n28348), .Z(n28178) );
  BUF U5813 ( .I(n28113), .Z(n27943) );
  BUF U5814 ( .I(n27878), .Z(n27708) );
  BUF U5815 ( .I(n27643), .Z(n27473) );
  BUF U5816 ( .I(n29288), .Z(n29119) );
  BUF U5817 ( .I(n29053), .Z(n28884) );
  BUF U5818 ( .I(n28818), .Z(n28649) );
  BUF U5819 ( .I(n28583), .Z(n28414) );
  BUF U5820 ( .I(n28348), .Z(n28179) );
  BUF U5821 ( .I(n28113), .Z(n27944) );
  BUF U5822 ( .I(n27878), .Z(n27709) );
  BUF U5823 ( .I(n27643), .Z(n27474) );
  BUF U5824 ( .I(n29287), .Z(n29120) );
  BUF U5825 ( .I(n29052), .Z(n28885) );
  BUF U5826 ( .I(n28817), .Z(n28650) );
  BUF U5827 ( .I(n28582), .Z(n28415) );
  BUF U5828 ( .I(n28347), .Z(n28180) );
  BUF U5829 ( .I(n28112), .Z(n27945) );
  BUF U5830 ( .I(n27877), .Z(n27710) );
  BUF U5831 ( .I(n27642), .Z(n27475) );
  BUF U5832 ( .I(n29287), .Z(n29121) );
  BUF U5833 ( .I(n29052), .Z(n28886) );
  BUF U5834 ( .I(n28817), .Z(n28651) );
  BUF U5835 ( .I(n28582), .Z(n28416) );
  BUF U5836 ( .I(n28347), .Z(n28181) );
  BUF U5837 ( .I(n28112), .Z(n27946) );
  BUF U5838 ( .I(n27877), .Z(n27711) );
  BUF U5839 ( .I(n27642), .Z(n27476) );
  BUF U5840 ( .I(n29287), .Z(n29122) );
  BUF U5841 ( .I(n29052), .Z(n28887) );
  BUF U5842 ( .I(n28817), .Z(n28652) );
  BUF U5843 ( .I(n28582), .Z(n28417) );
  BUF U5844 ( .I(n28347), .Z(n28182) );
  BUF U5845 ( .I(n28112), .Z(n27947) );
  BUF U5846 ( .I(n27877), .Z(n27712) );
  BUF U5847 ( .I(n27642), .Z(n27477) );
  BUF U5848 ( .I(n29286), .Z(n29123) );
  BUF U5849 ( .I(n29051), .Z(n28888) );
  BUF U5850 ( .I(n28816), .Z(n28653) );
  BUF U5851 ( .I(n28581), .Z(n28418) );
  BUF U5852 ( .I(n28346), .Z(n28183) );
  BUF U5853 ( .I(n28111), .Z(n27948) );
  BUF U5854 ( .I(n27876), .Z(n27713) );
  BUF U5855 ( .I(n27641), .Z(n27478) );
  BUF U5856 ( .I(n29286), .Z(n29124) );
  BUF U5857 ( .I(n29051), .Z(n28889) );
  BUF U5858 ( .I(n28816), .Z(n28654) );
  BUF U5859 ( .I(n28581), .Z(n28419) );
  BUF U5860 ( .I(n28346), .Z(n28184) );
  BUF U5861 ( .I(n28111), .Z(n27949) );
  BUF U5862 ( .I(n27876), .Z(n27714) );
  BUF U5863 ( .I(n27641), .Z(n27479) );
  BUF U5864 ( .I(n29286), .Z(n29125) );
  BUF U5865 ( .I(n29051), .Z(n28890) );
  BUF U5866 ( .I(n28816), .Z(n28655) );
  BUF U5867 ( .I(n28581), .Z(n28420) );
  BUF U5868 ( .I(n28346), .Z(n28185) );
  BUF U5869 ( .I(n28111), .Z(n27950) );
  BUF U5870 ( .I(n27876), .Z(n27715) );
  BUF U5871 ( .I(n27641), .Z(n27480) );
  BUF U5872 ( .I(n29285), .Z(n29126) );
  BUF U5873 ( .I(n29050), .Z(n28891) );
  BUF U5874 ( .I(n28815), .Z(n28656) );
  BUF U5875 ( .I(n28580), .Z(n28421) );
  BUF U5876 ( .I(n28345), .Z(n28186) );
  BUF U5877 ( .I(n28110), .Z(n27951) );
  BUF U5878 ( .I(n27875), .Z(n27716) );
  BUF U5879 ( .I(n27640), .Z(n27481) );
  BUF U5880 ( .I(n29285), .Z(n29127) );
  BUF U5881 ( .I(n29050), .Z(n28892) );
  BUF U5882 ( .I(n28815), .Z(n28657) );
  BUF U5883 ( .I(n28580), .Z(n28422) );
  BUF U5884 ( .I(n28345), .Z(n28187) );
  BUF U5885 ( .I(n28110), .Z(n27952) );
  BUF U5886 ( .I(n27875), .Z(n27717) );
  BUF U5887 ( .I(n27640), .Z(n27482) );
  BUF U5888 ( .I(n29285), .Z(n29128) );
  BUF U5889 ( .I(n29050), .Z(n28893) );
  BUF U5890 ( .I(n28815), .Z(n28658) );
  BUF U5891 ( .I(n28580), .Z(n28423) );
  BUF U5892 ( .I(n28345), .Z(n28188) );
  BUF U5893 ( .I(n28110), .Z(n27953) );
  BUF U5894 ( .I(n27875), .Z(n27718) );
  BUF U5895 ( .I(n27640), .Z(n27483) );
  BUF U5896 ( .I(n29284), .Z(n29129) );
  BUF U5897 ( .I(n29049), .Z(n28894) );
  BUF U5898 ( .I(n28814), .Z(n28659) );
  BUF U5899 ( .I(n28579), .Z(n28424) );
  BUF U5900 ( .I(n28344), .Z(n28189) );
  BUF U5901 ( .I(n28109), .Z(n27954) );
  BUF U5902 ( .I(n27874), .Z(n27719) );
  BUF U5903 ( .I(n27639), .Z(n27484) );
  BUF U5904 ( .I(n29284), .Z(n29130) );
  BUF U5905 ( .I(n29049), .Z(n28895) );
  BUF U5906 ( .I(n28814), .Z(n28660) );
  BUF U5907 ( .I(n28579), .Z(n28425) );
  BUF U5908 ( .I(n28344), .Z(n28190) );
  BUF U5909 ( .I(n28109), .Z(n27955) );
  BUF U5910 ( .I(n27874), .Z(n27720) );
  BUF U5911 ( .I(n27639), .Z(n27485) );
  BUF U5912 ( .I(n29284), .Z(n29131) );
  BUF U5913 ( .I(n29049), .Z(n28896) );
  BUF U5914 ( .I(n28814), .Z(n28661) );
  BUF U5915 ( .I(n28579), .Z(n28426) );
  BUF U5916 ( .I(n28344), .Z(n28191) );
  BUF U5917 ( .I(n28109), .Z(n27956) );
  BUF U5918 ( .I(n27874), .Z(n27721) );
  BUF U5919 ( .I(n27639), .Z(n27486) );
  BUF U5920 ( .I(n29283), .Z(n29132) );
  BUF U5921 ( .I(n29048), .Z(n28897) );
  BUF U5922 ( .I(n28813), .Z(n28662) );
  BUF U5923 ( .I(n28578), .Z(n28427) );
  BUF U5924 ( .I(n28343), .Z(n28192) );
  BUF U5925 ( .I(n28108), .Z(n27957) );
  BUF U5926 ( .I(n27873), .Z(n27722) );
  BUF U5927 ( .I(n27638), .Z(n27487) );
  BUF U5928 ( .I(n29283), .Z(n29133) );
  BUF U5929 ( .I(n29048), .Z(n28898) );
  BUF U5930 ( .I(n28813), .Z(n28663) );
  BUF U5931 ( .I(n28578), .Z(n28428) );
  BUF U5932 ( .I(n28343), .Z(n28193) );
  BUF U5933 ( .I(n28108), .Z(n27958) );
  BUF U5934 ( .I(n27873), .Z(n27723) );
  BUF U5935 ( .I(n27638), .Z(n27488) );
  BUF U5936 ( .I(n29283), .Z(n29134) );
  BUF U5937 ( .I(n29048), .Z(n28899) );
  BUF U5938 ( .I(n28813), .Z(n28664) );
  BUF U5939 ( .I(n28578), .Z(n28429) );
  BUF U5940 ( .I(n28343), .Z(n28194) );
  BUF U5941 ( .I(n28108), .Z(n27959) );
  BUF U5942 ( .I(n27873), .Z(n27724) );
  BUF U5943 ( .I(n27638), .Z(n27489) );
  BUF U5944 ( .I(n29282), .Z(n29135) );
  BUF U5945 ( .I(n29047), .Z(n28900) );
  BUF U5946 ( .I(n28812), .Z(n28665) );
  BUF U5947 ( .I(n28577), .Z(n28430) );
  BUF U5948 ( .I(n28342), .Z(n28195) );
  BUF U5949 ( .I(n28107), .Z(n27960) );
  BUF U5950 ( .I(n27872), .Z(n27725) );
  BUF U5951 ( .I(n27637), .Z(n27490) );
  BUF U5952 ( .I(n29282), .Z(n29136) );
  BUF U5953 ( .I(n29047), .Z(n28901) );
  BUF U5954 ( .I(n28812), .Z(n28666) );
  BUF U5955 ( .I(n28577), .Z(n28431) );
  BUF U5956 ( .I(n28342), .Z(n28196) );
  BUF U5957 ( .I(n28107), .Z(n27961) );
  BUF U5958 ( .I(n27872), .Z(n27726) );
  BUF U5959 ( .I(n27637), .Z(n27491) );
  BUF U5960 ( .I(n29282), .Z(n29137) );
  BUF U5961 ( .I(n29047), .Z(n28902) );
  BUF U5962 ( .I(n28812), .Z(n28667) );
  BUF U5963 ( .I(n28577), .Z(n28432) );
  BUF U5964 ( .I(n28342), .Z(n28197) );
  BUF U5965 ( .I(n28107), .Z(n27962) );
  BUF U5966 ( .I(n27872), .Z(n27727) );
  BUF U5967 ( .I(n27637), .Z(n27492) );
  BUF U5968 ( .I(n29281), .Z(n29138) );
  BUF U5969 ( .I(n29046), .Z(n28903) );
  BUF U5970 ( .I(n28811), .Z(n28668) );
  BUF U5971 ( .I(n28576), .Z(n28433) );
  BUF U5972 ( .I(n28341), .Z(n28198) );
  BUF U5973 ( .I(n28106), .Z(n27963) );
  BUF U5974 ( .I(n27871), .Z(n27728) );
  BUF U5975 ( .I(n27636), .Z(n27493) );
  BUF U5976 ( .I(n29281), .Z(n29139) );
  BUF U5977 ( .I(n29046), .Z(n28904) );
  BUF U5978 ( .I(n28811), .Z(n28669) );
  BUF U5979 ( .I(n28576), .Z(n28434) );
  BUF U5980 ( .I(n28341), .Z(n28199) );
  BUF U5981 ( .I(n28106), .Z(n27964) );
  BUF U5982 ( .I(n27871), .Z(n27729) );
  BUF U5983 ( .I(n27636), .Z(n27494) );
  BUF U5984 ( .I(n29281), .Z(n29140) );
  BUF U5985 ( .I(n29046), .Z(n28905) );
  BUF U5986 ( .I(n28811), .Z(n28670) );
  BUF U5987 ( .I(n28576), .Z(n28435) );
  BUF U5988 ( .I(n28341), .Z(n28200) );
  BUF U5989 ( .I(n28106), .Z(n27965) );
  BUF U5990 ( .I(n27871), .Z(n27730) );
  BUF U5991 ( .I(n27636), .Z(n27495) );
  BUF U5992 ( .I(n29280), .Z(n29141) );
  BUF U5993 ( .I(n29045), .Z(n28906) );
  BUF U5994 ( .I(n28810), .Z(n28671) );
  BUF U5995 ( .I(n28575), .Z(n28436) );
  BUF U5996 ( .I(n28340), .Z(n28201) );
  BUF U5997 ( .I(n28105), .Z(n27966) );
  BUF U5998 ( .I(n27870), .Z(n27731) );
  BUF U5999 ( .I(n27635), .Z(n27496) );
  BUF U6000 ( .I(n29280), .Z(n29142) );
  BUF U6001 ( .I(n29045), .Z(n28907) );
  BUF U6002 ( .I(n28810), .Z(n28672) );
  BUF U6003 ( .I(n28575), .Z(n28437) );
  BUF U6004 ( .I(n28340), .Z(n28202) );
  BUF U6005 ( .I(n28105), .Z(n27967) );
  BUF U6006 ( .I(n27870), .Z(n27732) );
  BUF U6007 ( .I(n27635), .Z(n27497) );
  BUF U6008 ( .I(n29280), .Z(n29143) );
  BUF U6009 ( .I(n29045), .Z(n28908) );
  BUF U6010 ( .I(n28810), .Z(n28673) );
  BUF U6011 ( .I(n28575), .Z(n28438) );
  BUF U6012 ( .I(n28340), .Z(n28203) );
  BUF U6013 ( .I(n28105), .Z(n27968) );
  BUF U6014 ( .I(n27870), .Z(n27733) );
  BUF U6015 ( .I(n27635), .Z(n27498) );
  BUF U6016 ( .I(n29279), .Z(n29144) );
  BUF U6017 ( .I(n29044), .Z(n28909) );
  BUF U6018 ( .I(n28809), .Z(n28674) );
  BUF U6019 ( .I(n28574), .Z(n28439) );
  BUF U6020 ( .I(n28339), .Z(n28204) );
  BUF U6021 ( .I(n28104), .Z(n27969) );
  BUF U6022 ( .I(n27869), .Z(n27734) );
  BUF U6023 ( .I(n27634), .Z(n27499) );
  BUF U6024 ( .I(n29279), .Z(n29145) );
  BUF U6025 ( .I(n29044), .Z(n28910) );
  BUF U6026 ( .I(n28809), .Z(n28675) );
  BUF U6027 ( .I(n28574), .Z(n28440) );
  BUF U6028 ( .I(n28339), .Z(n28205) );
  BUF U6029 ( .I(n28104), .Z(n27970) );
  BUF U6030 ( .I(n27869), .Z(n27735) );
  BUF U6031 ( .I(n27634), .Z(n27500) );
  BUF U6032 ( .I(n29279), .Z(n29146) );
  BUF U6033 ( .I(n29044), .Z(n28911) );
  BUF U6034 ( .I(n28809), .Z(n28676) );
  BUF U6035 ( .I(n28574), .Z(n28441) );
  BUF U6036 ( .I(n28339), .Z(n28206) );
  BUF U6037 ( .I(n28104), .Z(n27971) );
  BUF U6038 ( .I(n27869), .Z(n27736) );
  BUF U6039 ( .I(n27634), .Z(n27501) );
  BUF U6040 ( .I(n29278), .Z(n29147) );
  BUF U6041 ( .I(n29043), .Z(n28912) );
  BUF U6042 ( .I(n28808), .Z(n28677) );
  BUF U6043 ( .I(n28573), .Z(n28442) );
  BUF U6044 ( .I(n28338), .Z(n28207) );
  BUF U6045 ( .I(n28103), .Z(n27972) );
  BUF U6046 ( .I(n27868), .Z(n27737) );
  BUF U6047 ( .I(n27633), .Z(n27502) );
  BUF U6048 ( .I(n29278), .Z(n29148) );
  BUF U6049 ( .I(n29043), .Z(n28913) );
  BUF U6050 ( .I(n28808), .Z(n28678) );
  BUF U6051 ( .I(n28573), .Z(n28443) );
  BUF U6052 ( .I(n28338), .Z(n28208) );
  BUF U6053 ( .I(n28103), .Z(n27973) );
  BUF U6054 ( .I(n27868), .Z(n27738) );
  BUF U6055 ( .I(n27633), .Z(n27503) );
  BUF U6056 ( .I(n29278), .Z(n29149) );
  BUF U6057 ( .I(n29043), .Z(n28914) );
  BUF U6058 ( .I(n28808), .Z(n28679) );
  BUF U6059 ( .I(n28573), .Z(n28444) );
  BUF U6060 ( .I(n28338), .Z(n28209) );
  BUF U6061 ( .I(n28103), .Z(n27974) );
  BUF U6062 ( .I(n27868), .Z(n27739) );
  BUF U6063 ( .I(n27633), .Z(n27504) );
  BUF U6064 ( .I(n29277), .Z(n29150) );
  BUF U6065 ( .I(n29042), .Z(n28915) );
  BUF U6066 ( .I(n28807), .Z(n28680) );
  BUF U6067 ( .I(n28572), .Z(n28445) );
  BUF U6068 ( .I(n28337), .Z(n28210) );
  BUF U6069 ( .I(n28102), .Z(n27975) );
  BUF U6070 ( .I(n27867), .Z(n27740) );
  BUF U6071 ( .I(n27632), .Z(n27505) );
  BUF U6072 ( .I(n29277), .Z(n29151) );
  BUF U6073 ( .I(n29042), .Z(n28916) );
  BUF U6074 ( .I(n28807), .Z(n28681) );
  BUF U6075 ( .I(n28572), .Z(n28446) );
  BUF U6076 ( .I(n28337), .Z(n28211) );
  BUF U6077 ( .I(n28102), .Z(n27976) );
  BUF U6078 ( .I(n27867), .Z(n27741) );
  BUF U6079 ( .I(n27632), .Z(n27506) );
  BUF U6080 ( .I(n29277), .Z(n29152) );
  BUF U6081 ( .I(n29042), .Z(n28917) );
  BUF U6082 ( .I(n28807), .Z(n28682) );
  BUF U6083 ( .I(n28572), .Z(n28447) );
  BUF U6084 ( .I(n28337), .Z(n28212) );
  BUF U6085 ( .I(n28102), .Z(n27977) );
  BUF U6086 ( .I(n27867), .Z(n27742) );
  BUF U6087 ( .I(n27632), .Z(n27507) );
  BUF U6088 ( .I(n29276), .Z(n29153) );
  BUF U6089 ( .I(n29041), .Z(n28918) );
  BUF U6090 ( .I(n28806), .Z(n28683) );
  BUF U6091 ( .I(n28571), .Z(n28448) );
  BUF U6092 ( .I(n28336), .Z(n28213) );
  BUF U6093 ( .I(n28101), .Z(n27978) );
  BUF U6094 ( .I(n27866), .Z(n27743) );
  BUF U6095 ( .I(n27631), .Z(n27508) );
  BUF U6096 ( .I(n29276), .Z(n29154) );
  BUF U6097 ( .I(n29041), .Z(n28919) );
  BUF U6098 ( .I(n28806), .Z(n28684) );
  BUF U6099 ( .I(n28571), .Z(n28449) );
  BUF U6100 ( .I(n28336), .Z(n28214) );
  BUF U6101 ( .I(n28101), .Z(n27979) );
  BUF U6102 ( .I(n27866), .Z(n27744) );
  BUF U6103 ( .I(n27631), .Z(n27509) );
  BUF U6104 ( .I(n29276), .Z(n29155) );
  BUF U6105 ( .I(n29041), .Z(n28920) );
  BUF U6106 ( .I(n28806), .Z(n28685) );
  BUF U6107 ( .I(n28571), .Z(n28450) );
  BUF U6108 ( .I(n28336), .Z(n28215) );
  BUF U6109 ( .I(n28101), .Z(n27980) );
  BUF U6110 ( .I(n27866), .Z(n27745) );
  BUF U6111 ( .I(n27631), .Z(n27510) );
  BUF U6112 ( .I(n29275), .Z(n29156) );
  BUF U6113 ( .I(n29040), .Z(n28921) );
  BUF U6114 ( .I(n28805), .Z(n28686) );
  BUF U6115 ( .I(n28570), .Z(n28451) );
  BUF U6116 ( .I(n28335), .Z(n28216) );
  BUF U6117 ( .I(n28100), .Z(n27981) );
  BUF U6118 ( .I(n27865), .Z(n27746) );
  BUF U6119 ( .I(n27630), .Z(n27511) );
  BUF U6120 ( .I(n29275), .Z(n29157) );
  BUF U6121 ( .I(n29040), .Z(n28922) );
  BUF U6122 ( .I(n28805), .Z(n28687) );
  BUF U6123 ( .I(n28570), .Z(n28452) );
  BUF U6124 ( .I(n28335), .Z(n28217) );
  BUF U6125 ( .I(n28100), .Z(n27982) );
  BUF U6126 ( .I(n27865), .Z(n27747) );
  BUF U6127 ( .I(n27630), .Z(n27512) );
  BUF U6128 ( .I(n29275), .Z(n29158) );
  BUF U6129 ( .I(n29040), .Z(n28923) );
  BUF U6130 ( .I(n28805), .Z(n28688) );
  BUF U6131 ( .I(n28570), .Z(n28453) );
  BUF U6132 ( .I(n28335), .Z(n28218) );
  BUF U6133 ( .I(n28100), .Z(n27983) );
  BUF U6134 ( .I(n27865), .Z(n27748) );
  BUF U6135 ( .I(n27630), .Z(n27513) );
  BUF U6136 ( .I(n29274), .Z(n29159) );
  BUF U6137 ( .I(n29039), .Z(n28924) );
  BUF U6138 ( .I(n28804), .Z(n28689) );
  BUF U6139 ( .I(n28569), .Z(n28454) );
  BUF U6140 ( .I(n28334), .Z(n28219) );
  BUF U6141 ( .I(n28099), .Z(n27984) );
  BUF U6142 ( .I(n27864), .Z(n27749) );
  BUF U6143 ( .I(n27629), .Z(n27514) );
  BUF U6144 ( .I(n29274), .Z(n29160) );
  BUF U6145 ( .I(n29039), .Z(n28925) );
  BUF U6146 ( .I(n28804), .Z(n28690) );
  BUF U6147 ( .I(n28569), .Z(n28455) );
  BUF U6148 ( .I(n28334), .Z(n28220) );
  BUF U6149 ( .I(n28099), .Z(n27985) );
  BUF U6150 ( .I(n27864), .Z(n27750) );
  BUF U6151 ( .I(n27629), .Z(n27515) );
  BUF U6152 ( .I(n29274), .Z(n29161) );
  BUF U6153 ( .I(n29039), .Z(n28926) );
  BUF U6154 ( .I(n28804), .Z(n28691) );
  BUF U6155 ( .I(n28569), .Z(n28456) );
  BUF U6156 ( .I(n28334), .Z(n28221) );
  BUF U6157 ( .I(n28099), .Z(n27986) );
  BUF U6158 ( .I(n27864), .Z(n27751) );
  BUF U6159 ( .I(n27629), .Z(n27516) );
  BUF U6160 ( .I(n29273), .Z(n29162) );
  BUF U6161 ( .I(n29038), .Z(n28927) );
  BUF U6162 ( .I(n28803), .Z(n28692) );
  BUF U6163 ( .I(n28568), .Z(n28457) );
  BUF U6164 ( .I(n28333), .Z(n28222) );
  BUF U6165 ( .I(n28098), .Z(n27987) );
  BUF U6166 ( .I(n27863), .Z(n27752) );
  BUF U6167 ( .I(n27628), .Z(n27517) );
  BUF U6168 ( .I(n29273), .Z(n29163) );
  BUF U6169 ( .I(n29038), .Z(n28928) );
  BUF U6170 ( .I(n28803), .Z(n28693) );
  BUF U6171 ( .I(n28568), .Z(n28458) );
  BUF U6172 ( .I(n28333), .Z(n28223) );
  BUF U6173 ( .I(n28098), .Z(n27988) );
  BUF U6174 ( .I(n27863), .Z(n27753) );
  BUF U6175 ( .I(n27628), .Z(n27518) );
  BUF U6176 ( .I(n29273), .Z(n29164) );
  BUF U6177 ( .I(n29038), .Z(n28929) );
  BUF U6178 ( .I(n28803), .Z(n28694) );
  BUF U6179 ( .I(n28568), .Z(n28459) );
  BUF U6180 ( .I(n28333), .Z(n28224) );
  BUF U6181 ( .I(n28098), .Z(n27989) );
  BUF U6182 ( .I(n27863), .Z(n27754) );
  BUF U6183 ( .I(n27628), .Z(n27519) );
  BUF U6184 ( .I(n29272), .Z(n29165) );
  BUF U6185 ( .I(n29037), .Z(n28930) );
  BUF U6186 ( .I(n28802), .Z(n28695) );
  BUF U6187 ( .I(n28567), .Z(n28460) );
  BUF U6188 ( .I(n28332), .Z(n28225) );
  BUF U6189 ( .I(n28097), .Z(n27990) );
  BUF U6190 ( .I(n27862), .Z(n27755) );
  BUF U6191 ( .I(n27627), .Z(n27520) );
  BUF U6192 ( .I(n29272), .Z(n29166) );
  BUF U6193 ( .I(n29037), .Z(n28931) );
  BUF U6194 ( .I(n28802), .Z(n28696) );
  BUF U6195 ( .I(n28567), .Z(n28461) );
  BUF U6196 ( .I(n28332), .Z(n28226) );
  BUF U6197 ( .I(n28097), .Z(n27991) );
  BUF U6198 ( .I(n27862), .Z(n27756) );
  BUF U6199 ( .I(n27627), .Z(n27521) );
  BUF U6200 ( .I(n29272), .Z(n29167) );
  BUF U6201 ( .I(n29037), .Z(n28932) );
  BUF U6202 ( .I(n28802), .Z(n28697) );
  BUF U6203 ( .I(n28567), .Z(n28462) );
  BUF U6204 ( .I(n28332), .Z(n28227) );
  BUF U6205 ( .I(n28097), .Z(n27992) );
  BUF U6206 ( .I(n27862), .Z(n27757) );
  BUF U6207 ( .I(n27627), .Z(n27522) );
  BUF U6208 ( .I(n29271), .Z(n29168) );
  BUF U6209 ( .I(n29036), .Z(n28933) );
  BUF U6210 ( .I(n28801), .Z(n28698) );
  BUF U6211 ( .I(n28566), .Z(n28463) );
  BUF U6212 ( .I(n28331), .Z(n28228) );
  BUF U6213 ( .I(n28096), .Z(n27993) );
  BUF U6214 ( .I(n27861), .Z(n27758) );
  BUF U6215 ( .I(n27626), .Z(n27523) );
  BUF U6216 ( .I(n29271), .Z(n29169) );
  BUF U6217 ( .I(n29036), .Z(n28934) );
  BUF U6218 ( .I(n28801), .Z(n28699) );
  BUF U6219 ( .I(n28566), .Z(n28464) );
  BUF U6220 ( .I(n28331), .Z(n28229) );
  BUF U6221 ( .I(n28096), .Z(n27994) );
  BUF U6222 ( .I(n27861), .Z(n27759) );
  BUF U6223 ( .I(n27626), .Z(n27524) );
  BUF U6224 ( .I(n29271), .Z(n29170) );
  BUF U6225 ( .I(n29036), .Z(n28935) );
  BUF U6226 ( .I(n28801), .Z(n28700) );
  BUF U6227 ( .I(n28566), .Z(n28465) );
  BUF U6228 ( .I(n28331), .Z(n28230) );
  BUF U6229 ( .I(n28096), .Z(n27995) );
  BUF U6230 ( .I(n27861), .Z(n27760) );
  BUF U6231 ( .I(n27626), .Z(n27525) );
  BUF U6232 ( .I(n29270), .Z(n29171) );
  BUF U6233 ( .I(n29035), .Z(n28936) );
  BUF U6234 ( .I(n28800), .Z(n28701) );
  BUF U6235 ( .I(n28565), .Z(n28466) );
  BUF U6236 ( .I(n28330), .Z(n28231) );
  BUF U6237 ( .I(n28095), .Z(n27996) );
  BUF U6238 ( .I(n27860), .Z(n27761) );
  BUF U6239 ( .I(n27625), .Z(n27526) );
  BUF U6240 ( .I(n29270), .Z(n29172) );
  BUF U6241 ( .I(n29035), .Z(n28937) );
  BUF U6242 ( .I(n28800), .Z(n28702) );
  BUF U6243 ( .I(n28565), .Z(n28467) );
  BUF U6244 ( .I(n28330), .Z(n28232) );
  BUF U6245 ( .I(n28095), .Z(n27997) );
  BUF U6246 ( .I(n27860), .Z(n27762) );
  BUF U6247 ( .I(n27625), .Z(n27527) );
  BUF U6248 ( .I(n29270), .Z(n29173) );
  BUF U6249 ( .I(n29035), .Z(n28938) );
  BUF U6250 ( .I(n28800), .Z(n28703) );
  BUF U6251 ( .I(n28565), .Z(n28468) );
  BUF U6252 ( .I(n28330), .Z(n28233) );
  BUF U6253 ( .I(n28095), .Z(n27998) );
  BUF U6254 ( .I(n27860), .Z(n27763) );
  BUF U6255 ( .I(n27625), .Z(n27528) );
  BUF U6256 ( .I(n29269), .Z(n29174) );
  BUF U6257 ( .I(n29034), .Z(n28939) );
  BUF U6258 ( .I(n28799), .Z(n28704) );
  BUF U6259 ( .I(n28564), .Z(n28469) );
  BUF U6260 ( .I(n28329), .Z(n28234) );
  BUF U6261 ( .I(n28094), .Z(n27999) );
  BUF U6262 ( .I(n27859), .Z(n27764) );
  BUF U6263 ( .I(n27624), .Z(n27529) );
  BUF U6264 ( .I(n29269), .Z(n29175) );
  BUF U6265 ( .I(n29034), .Z(n28940) );
  BUF U6266 ( .I(n28799), .Z(n28705) );
  BUF U6267 ( .I(n28564), .Z(n28470) );
  BUF U6268 ( .I(n28329), .Z(n28235) );
  BUF U6269 ( .I(n28094), .Z(n28000) );
  BUF U6270 ( .I(n27859), .Z(n27765) );
  BUF U6271 ( .I(n27624), .Z(n27530) );
  BUF U6272 ( .I(n29269), .Z(n29176) );
  BUF U6273 ( .I(n29034), .Z(n28941) );
  BUF U6274 ( .I(n28799), .Z(n28706) );
  BUF U6275 ( .I(n28564), .Z(n28471) );
  BUF U6276 ( .I(n28329), .Z(n28236) );
  BUF U6277 ( .I(n28094), .Z(n28001) );
  BUF U6278 ( .I(n27859), .Z(n27766) );
  BUF U6279 ( .I(n27624), .Z(n27531) );
  BUF U6280 ( .I(n29268), .Z(n29177) );
  BUF U6281 ( .I(n29033), .Z(n28942) );
  BUF U6282 ( .I(n28798), .Z(n28707) );
  BUF U6283 ( .I(n28563), .Z(n28472) );
  BUF U6284 ( .I(n28328), .Z(n28237) );
  BUF U6285 ( .I(n28093), .Z(n28002) );
  BUF U6286 ( .I(n27858), .Z(n27767) );
  BUF U6287 ( .I(n27623), .Z(n27532) );
  BUF U6288 ( .I(n29268), .Z(n29178) );
  BUF U6289 ( .I(n29033), .Z(n28943) );
  BUF U6290 ( .I(n28798), .Z(n28708) );
  BUF U6291 ( .I(n28563), .Z(n28473) );
  BUF U6292 ( .I(n28328), .Z(n28238) );
  BUF U6293 ( .I(n28093), .Z(n28003) );
  BUF U6294 ( .I(n27858), .Z(n27768) );
  BUF U6295 ( .I(n27623), .Z(n27533) );
  BUF U6296 ( .I(n29268), .Z(n29179) );
  BUF U6297 ( .I(n29033), .Z(n28944) );
  BUF U6298 ( .I(n28798), .Z(n28709) );
  BUF U6299 ( .I(n28563), .Z(n28474) );
  BUF U6300 ( .I(n28328), .Z(n28239) );
  BUF U6301 ( .I(n28093), .Z(n28004) );
  BUF U6302 ( .I(n27858), .Z(n27769) );
  BUF U6303 ( .I(n27623), .Z(n27534) );
  BUF U6304 ( .I(n29267), .Z(n29180) );
  BUF U6305 ( .I(n29032), .Z(n28945) );
  BUF U6306 ( .I(n28797), .Z(n28710) );
  BUF U6307 ( .I(n28562), .Z(n28475) );
  BUF U6308 ( .I(n28327), .Z(n28240) );
  BUF U6309 ( .I(n28092), .Z(n28005) );
  BUF U6310 ( .I(n27857), .Z(n27770) );
  BUF U6311 ( .I(n27622), .Z(n27535) );
  BUF U6312 ( .I(n29267), .Z(n29181) );
  BUF U6313 ( .I(n29032), .Z(n28946) );
  BUF U6314 ( .I(n28797), .Z(n28711) );
  BUF U6315 ( .I(n28562), .Z(n28476) );
  BUF U6316 ( .I(n28327), .Z(n28241) );
  BUF U6317 ( .I(n28092), .Z(n28006) );
  BUF U6318 ( .I(n27857), .Z(n27771) );
  BUF U6319 ( .I(n27622), .Z(n27536) );
  BUF U6320 ( .I(n29267), .Z(n29182) );
  BUF U6321 ( .I(n29032), .Z(n28947) );
  BUF U6322 ( .I(n28797), .Z(n28712) );
  BUF U6323 ( .I(n28562), .Z(n28477) );
  BUF U6324 ( .I(n28327), .Z(n28242) );
  BUF U6325 ( .I(n28092), .Z(n28007) );
  BUF U6326 ( .I(n27857), .Z(n27772) );
  BUF U6327 ( .I(n27622), .Z(n27537) );
  BUF U6328 ( .I(n29266), .Z(n29183) );
  BUF U6329 ( .I(n29031), .Z(n28948) );
  BUF U6330 ( .I(n28796), .Z(n28713) );
  BUF U6331 ( .I(n28561), .Z(n28478) );
  BUF U6332 ( .I(n28326), .Z(n28243) );
  BUF U6333 ( .I(n28091), .Z(n28008) );
  BUF U6334 ( .I(n27856), .Z(n27773) );
  BUF U6335 ( .I(n27621), .Z(n27538) );
  BUF U6336 ( .I(n29266), .Z(n29184) );
  BUF U6337 ( .I(n29031), .Z(n28949) );
  BUF U6338 ( .I(n28796), .Z(n28714) );
  BUF U6339 ( .I(n28561), .Z(n28479) );
  BUF U6340 ( .I(n28326), .Z(n28244) );
  BUF U6341 ( .I(n28091), .Z(n28009) );
  BUF U6342 ( .I(n27856), .Z(n27774) );
  BUF U6343 ( .I(n27621), .Z(n27539) );
  BUF U6344 ( .I(n29266), .Z(n29185) );
  BUF U6345 ( .I(n29031), .Z(n28950) );
  BUF U6346 ( .I(n28796), .Z(n28715) );
  BUF U6347 ( .I(n28561), .Z(n28480) );
  BUF U6348 ( .I(n28326), .Z(n28245) );
  BUF U6349 ( .I(n28091), .Z(n28010) );
  BUF U6350 ( .I(n27856), .Z(n27775) );
  BUF U6351 ( .I(n27621), .Z(n27540) );
  BUF U6352 ( .I(n29265), .Z(n29186) );
  BUF U6353 ( .I(n29030), .Z(n28951) );
  BUF U6354 ( .I(n28795), .Z(n28716) );
  BUF U6355 ( .I(n28560), .Z(n28481) );
  BUF U6356 ( .I(n28325), .Z(n28246) );
  BUF U6357 ( .I(n28090), .Z(n28011) );
  BUF U6358 ( .I(n27855), .Z(n27776) );
  BUF U6359 ( .I(n27620), .Z(n27541) );
  BUF U6360 ( .I(n29265), .Z(n29187) );
  BUF U6361 ( .I(n29030), .Z(n28952) );
  BUF U6362 ( .I(n28795), .Z(n28717) );
  BUF U6363 ( .I(n28560), .Z(n28482) );
  BUF U6364 ( .I(n28325), .Z(n28247) );
  BUF U6365 ( .I(n28090), .Z(n28012) );
  BUF U6366 ( .I(n27855), .Z(n27777) );
  BUF U6367 ( .I(n27620), .Z(n27542) );
  BUF U6368 ( .I(n29265), .Z(n29188) );
  BUF U6369 ( .I(n29030), .Z(n28953) );
  BUF U6370 ( .I(n28795), .Z(n28718) );
  BUF U6371 ( .I(n28560), .Z(n28483) );
  BUF U6372 ( .I(n28325), .Z(n28248) );
  BUF U6373 ( .I(n28090), .Z(n28013) );
  BUF U6374 ( .I(n27855), .Z(n27778) );
  BUF U6375 ( .I(n27620), .Z(n27543) );
  BUF U6376 ( .I(n29264), .Z(n29189) );
  BUF U6377 ( .I(n29029), .Z(n28954) );
  BUF U6378 ( .I(n28794), .Z(n28719) );
  BUF U6379 ( .I(n28559), .Z(n28484) );
  BUF U6380 ( .I(n28324), .Z(n28249) );
  BUF U6381 ( .I(n28089), .Z(n28014) );
  BUF U6382 ( .I(n27854), .Z(n27779) );
  BUF U6383 ( .I(n27619), .Z(n27544) );
  BUF U6384 ( .I(n29264), .Z(n29190) );
  BUF U6385 ( .I(n29029), .Z(n28955) );
  BUF U6386 ( .I(n28794), .Z(n28720) );
  BUF U6387 ( .I(n28559), .Z(n28485) );
  BUF U6388 ( .I(n28324), .Z(n28250) );
  BUF U6389 ( .I(n28089), .Z(n28015) );
  BUF U6390 ( .I(n27854), .Z(n27780) );
  BUF U6391 ( .I(n27619), .Z(n27545) );
  BUF U6392 ( .I(n29264), .Z(n29191) );
  BUF U6393 ( .I(n29029), .Z(n28956) );
  BUF U6394 ( .I(n28794), .Z(n28721) );
  BUF U6395 ( .I(n28559), .Z(n28486) );
  BUF U6396 ( .I(n28324), .Z(n28251) );
  BUF U6397 ( .I(n28089), .Z(n28016) );
  BUF U6398 ( .I(n27854), .Z(n27781) );
  BUF U6399 ( .I(n27619), .Z(n27546) );
  BUF U6400 ( .I(n29263), .Z(n29192) );
  BUF U6401 ( .I(n29028), .Z(n28957) );
  BUF U6402 ( .I(n28793), .Z(n28722) );
  BUF U6403 ( .I(n28558), .Z(n28487) );
  BUF U6404 ( .I(n28323), .Z(n28252) );
  BUF U6405 ( .I(n28088), .Z(n28017) );
  BUF U6406 ( .I(n27853), .Z(n27782) );
  BUF U6407 ( .I(n27618), .Z(n27547) );
  BUF U6408 ( .I(n29263), .Z(n29193) );
  BUF U6409 ( .I(n29028), .Z(n28958) );
  BUF U6410 ( .I(n28793), .Z(n28723) );
  BUF U6411 ( .I(n28558), .Z(n28488) );
  BUF U6412 ( .I(n28323), .Z(n28253) );
  BUF U6413 ( .I(n28088), .Z(n28018) );
  BUF U6414 ( .I(n27853), .Z(n27783) );
  BUF U6415 ( .I(n27618), .Z(n27548) );
  BUF U6416 ( .I(n29263), .Z(n29194) );
  BUF U6417 ( .I(n29028), .Z(n28959) );
  BUF U6418 ( .I(n28793), .Z(n28724) );
  BUF U6419 ( .I(n28558), .Z(n28489) );
  BUF U6420 ( .I(n28323), .Z(n28254) );
  BUF U6421 ( .I(n28088), .Z(n28019) );
  BUF U6422 ( .I(n27853), .Z(n27784) );
  BUF U6423 ( .I(n27618), .Z(n27549) );
  BUF U6424 ( .I(n29262), .Z(n29195) );
  BUF U6425 ( .I(n29027), .Z(n28960) );
  BUF U6426 ( .I(n28792), .Z(n28725) );
  BUF U6427 ( .I(n28557), .Z(n28490) );
  BUF U6428 ( .I(n28322), .Z(n28255) );
  BUF U6429 ( .I(n28087), .Z(n28020) );
  BUF U6430 ( .I(n27852), .Z(n27785) );
  BUF U6431 ( .I(n27617), .Z(n27550) );
  BUF U6432 ( .I(n29262), .Z(n29196) );
  BUF U6433 ( .I(n29027), .Z(n28961) );
  BUF U6434 ( .I(n28792), .Z(n28726) );
  BUF U6435 ( .I(n28557), .Z(n28491) );
  BUF U6436 ( .I(n28322), .Z(n28256) );
  BUF U6437 ( .I(n28087), .Z(n28021) );
  BUF U6438 ( .I(n27852), .Z(n27786) );
  BUF U6439 ( .I(n27617), .Z(n27551) );
  BUF U6440 ( .I(n29262), .Z(n29197) );
  BUF U6441 ( .I(n29027), .Z(n28962) );
  BUF U6442 ( .I(n28792), .Z(n28727) );
  BUF U6443 ( .I(n28557), .Z(n28492) );
  BUF U6444 ( .I(n28322), .Z(n28257) );
  BUF U6445 ( .I(n28087), .Z(n28022) );
  BUF U6446 ( .I(n27852), .Z(n27787) );
  BUF U6447 ( .I(n27617), .Z(n27552) );
  BUF U6448 ( .I(n29261), .Z(n29198) );
  BUF U6449 ( .I(n29026), .Z(n28963) );
  BUF U6450 ( .I(n28791), .Z(n28728) );
  BUF U6451 ( .I(n28556), .Z(n28493) );
  BUF U6452 ( .I(n28321), .Z(n28258) );
  BUF U6453 ( .I(n28086), .Z(n28023) );
  BUF U6454 ( .I(n27851), .Z(n27788) );
  BUF U6455 ( .I(n27616), .Z(n27553) );
  BUF U6456 ( .I(n29261), .Z(n29199) );
  BUF U6457 ( .I(n29026), .Z(n28964) );
  BUF U6458 ( .I(n28791), .Z(n28729) );
  BUF U6459 ( .I(n28556), .Z(n28494) );
  BUF U6460 ( .I(n28321), .Z(n28259) );
  BUF U6461 ( .I(n28086), .Z(n28024) );
  BUF U6462 ( .I(n27851), .Z(n27789) );
  BUF U6463 ( .I(n27616), .Z(n27554) );
  BUF U6464 ( .I(n29261), .Z(n29200) );
  BUF U6465 ( .I(n29026), .Z(n28965) );
  BUF U6466 ( .I(n28791), .Z(n28730) );
  BUF U6467 ( .I(n28556), .Z(n28495) );
  BUF U6468 ( .I(n28321), .Z(n28260) );
  BUF U6469 ( .I(n28086), .Z(n28025) );
  BUF U6470 ( .I(n27851), .Z(n27790) );
  BUF U6471 ( .I(n27616), .Z(n27555) );
  BUF U6472 ( .I(n29260), .Z(n29201) );
  BUF U6473 ( .I(n29025), .Z(n28966) );
  BUF U6474 ( .I(n28790), .Z(n28731) );
  BUF U6475 ( .I(n28555), .Z(n28496) );
  BUF U6476 ( .I(n28320), .Z(n28261) );
  BUF U6477 ( .I(n28085), .Z(n28026) );
  BUF U6478 ( .I(n27850), .Z(n27791) );
  BUF U6479 ( .I(n27615), .Z(n27556) );
  BUF U6480 ( .I(n29260), .Z(n29202) );
  BUF U6481 ( .I(n29025), .Z(n28967) );
  BUF U6482 ( .I(n28790), .Z(n28732) );
  BUF U6483 ( .I(n28555), .Z(n28497) );
  BUF U6484 ( .I(n28320), .Z(n28262) );
  BUF U6485 ( .I(n28085), .Z(n28027) );
  BUF U6486 ( .I(n27850), .Z(n27792) );
  BUF U6487 ( .I(n27615), .Z(n27557) );
  BUF U6488 ( .I(n29260), .Z(n29203) );
  BUF U6489 ( .I(n29025), .Z(n28968) );
  BUF U6490 ( .I(n28790), .Z(n28733) );
  BUF U6491 ( .I(n28555), .Z(n28498) );
  BUF U6492 ( .I(n28320), .Z(n28263) );
  BUF U6493 ( .I(n28085), .Z(n28028) );
  BUF U6494 ( .I(n27850), .Z(n27793) );
  BUF U6495 ( .I(n27615), .Z(n27558) );
  BUF U6496 ( .I(n29259), .Z(n29204) );
  BUF U6497 ( .I(n29024), .Z(n28969) );
  BUF U6498 ( .I(n28789), .Z(n28734) );
  BUF U6499 ( .I(n28554), .Z(n28499) );
  BUF U6500 ( .I(n28319), .Z(n28264) );
  BUF U6501 ( .I(n28084), .Z(n28029) );
  BUF U6502 ( .I(n27849), .Z(n27794) );
  BUF U6503 ( .I(n27614), .Z(n27559) );
  BUF U6504 ( .I(n29259), .Z(n29205) );
  BUF U6505 ( .I(n29024), .Z(n28970) );
  BUF U6506 ( .I(n28789), .Z(n28735) );
  BUF U6507 ( .I(n28554), .Z(n28500) );
  BUF U6508 ( .I(n28319), .Z(n28265) );
  BUF U6509 ( .I(n28084), .Z(n28030) );
  BUF U6510 ( .I(n27849), .Z(n27795) );
  BUF U6511 ( .I(n27614), .Z(n27560) );
  BUF U6512 ( .I(n29259), .Z(n29206) );
  BUF U6513 ( .I(n29024), .Z(n28971) );
  BUF U6514 ( .I(n28789), .Z(n28736) );
  BUF U6515 ( .I(n28554), .Z(n28501) );
  BUF U6516 ( .I(n28319), .Z(n28266) );
  BUF U6517 ( .I(n28084), .Z(n28031) );
  BUF U6518 ( .I(n27849), .Z(n27796) );
  BUF U6519 ( .I(n27614), .Z(n27561) );
  BUF U6520 ( .I(n29258), .Z(n29207) );
  BUF U6521 ( .I(n29023), .Z(n28972) );
  BUF U6522 ( .I(n28788), .Z(n28737) );
  BUF U6523 ( .I(n28553), .Z(n28502) );
  BUF U6524 ( .I(n28318), .Z(n28267) );
  BUF U6525 ( .I(n28083), .Z(n28032) );
  BUF U6526 ( .I(n27848), .Z(n27797) );
  BUF U6527 ( .I(n27613), .Z(n27562) );
  BUF U6528 ( .I(n29258), .Z(n29208) );
  BUF U6529 ( .I(n29023), .Z(n28973) );
  BUF U6530 ( .I(n28788), .Z(n28738) );
  BUF U6531 ( .I(n28553), .Z(n28503) );
  BUF U6532 ( .I(n28318), .Z(n28268) );
  BUF U6533 ( .I(n28083), .Z(n28033) );
  BUF U6534 ( .I(n27848), .Z(n27798) );
  BUF U6535 ( .I(n27613), .Z(n27563) );
  BUF U6536 ( .I(n29258), .Z(n29209) );
  BUF U6537 ( .I(n29023), .Z(n28974) );
  BUF U6538 ( .I(n28788), .Z(n28739) );
  BUF U6539 ( .I(n28553), .Z(n28504) );
  BUF U6540 ( .I(n28318), .Z(n28269) );
  BUF U6541 ( .I(n28083), .Z(n28034) );
  BUF U6542 ( .I(n27848), .Z(n27799) );
  BUF U6543 ( .I(n27613), .Z(n27564) );
  BUF U6544 ( .I(n29257), .Z(n29210) );
  BUF U6545 ( .I(n29022), .Z(n28975) );
  BUF U6546 ( .I(n28787), .Z(n28740) );
  BUF U6547 ( .I(n28552), .Z(n28505) );
  BUF U6548 ( .I(n28317), .Z(n28270) );
  BUF U6549 ( .I(n28082), .Z(n28035) );
  BUF U6550 ( .I(n27847), .Z(n27800) );
  BUF U6551 ( .I(n27612), .Z(n27565) );
  BUF U6552 ( .I(n29257), .Z(n29211) );
  BUF U6553 ( .I(n29022), .Z(n28976) );
  BUF U6554 ( .I(n28787), .Z(n28741) );
  BUF U6555 ( .I(n28552), .Z(n28506) );
  BUF U6556 ( .I(n28317), .Z(n28271) );
  BUF U6557 ( .I(n28082), .Z(n28036) );
  BUF U6558 ( .I(n27847), .Z(n27801) );
  BUF U6559 ( .I(n27612), .Z(n27566) );
  BUF U6560 ( .I(n29257), .Z(n29212) );
  BUF U6561 ( .I(n29022), .Z(n28977) );
  BUF U6562 ( .I(n28787), .Z(n28742) );
  BUF U6563 ( .I(n28552), .Z(n28507) );
  BUF U6564 ( .I(n28317), .Z(n28272) );
  BUF U6565 ( .I(n28082), .Z(n28037) );
  BUF U6566 ( .I(n27847), .Z(n27802) );
  BUF U6567 ( .I(n27612), .Z(n27567) );
  BUF U6568 ( .I(n29256), .Z(n29213) );
  BUF U6569 ( .I(n29021), .Z(n28978) );
  BUF U6570 ( .I(n28786), .Z(n28743) );
  BUF U6571 ( .I(n28551), .Z(n28508) );
  BUF U6572 ( .I(n28316), .Z(n28273) );
  BUF U6573 ( .I(n28081), .Z(n28038) );
  BUF U6574 ( .I(n27846), .Z(n27803) );
  BUF U6575 ( .I(n27611), .Z(n27568) );
  BUF U6576 ( .I(n29256), .Z(n29214) );
  BUF U6577 ( .I(n29021), .Z(n28979) );
  BUF U6578 ( .I(n28786), .Z(n28744) );
  BUF U6579 ( .I(n28551), .Z(n28509) );
  BUF U6580 ( .I(n28316), .Z(n28274) );
  BUF U6581 ( .I(n28081), .Z(n28039) );
  BUF U6582 ( .I(n27846), .Z(n27804) );
  BUF U6583 ( .I(n27611), .Z(n27569) );
  BUF U6584 ( .I(n29256), .Z(n29215) );
  BUF U6585 ( .I(n29021), .Z(n28980) );
  BUF U6586 ( .I(n28786), .Z(n28745) );
  BUF U6587 ( .I(n28551), .Z(n28510) );
  BUF U6588 ( .I(n28316), .Z(n28275) );
  BUF U6589 ( .I(n28081), .Z(n28040) );
  BUF U6590 ( .I(n27846), .Z(n27805) );
  BUF U6591 ( .I(n27611), .Z(n27570) );
  BUF U6592 ( .I(n29255), .Z(n29216) );
  BUF U6593 ( .I(n29020), .Z(n28981) );
  BUF U6594 ( .I(n28785), .Z(n28746) );
  BUF U6595 ( .I(n28550), .Z(n28511) );
  BUF U6596 ( .I(n28315), .Z(n28276) );
  BUF U6597 ( .I(n28080), .Z(n28041) );
  BUF U6598 ( .I(n27845), .Z(n27806) );
  BUF U6599 ( .I(n27610), .Z(n27571) );
  BUF U6600 ( .I(n29255), .Z(n29217) );
  BUF U6601 ( .I(n29020), .Z(n28982) );
  BUF U6602 ( .I(n28785), .Z(n28747) );
  BUF U6603 ( .I(n28550), .Z(n28512) );
  BUF U6604 ( .I(n28315), .Z(n28277) );
  BUF U6605 ( .I(n28080), .Z(n28042) );
  BUF U6606 ( .I(n27845), .Z(n27807) );
  BUF U6607 ( .I(n27610), .Z(n27572) );
  BUF U6608 ( .I(n29255), .Z(n29218) );
  BUF U6609 ( .I(n29020), .Z(n28983) );
  BUF U6610 ( .I(n28785), .Z(n28748) );
  BUF U6611 ( .I(n28550), .Z(n28513) );
  BUF U6612 ( .I(n28315), .Z(n28278) );
  BUF U6613 ( .I(n28080), .Z(n28043) );
  BUF U6614 ( .I(n27845), .Z(n27808) );
  BUF U6615 ( .I(n27610), .Z(n27573) );
  BUF U6616 ( .I(n29254), .Z(n29219) );
  BUF U6617 ( .I(n29019), .Z(n28984) );
  BUF U6618 ( .I(n28784), .Z(n28749) );
  BUF U6619 ( .I(n28549), .Z(n28514) );
  BUF U6620 ( .I(n28314), .Z(n28279) );
  BUF U6621 ( .I(n28079), .Z(n28044) );
  BUF U6622 ( .I(n27844), .Z(n27809) );
  BUF U6623 ( .I(n27609), .Z(n27574) );
  BUF U6624 ( .I(n29254), .Z(n29220) );
  BUF U6625 ( .I(n29019), .Z(n28985) );
  BUF U6626 ( .I(n28784), .Z(n28750) );
  BUF U6627 ( .I(n28549), .Z(n28515) );
  BUF U6628 ( .I(n28314), .Z(n28280) );
  BUF U6629 ( .I(n28079), .Z(n28045) );
  BUF U6630 ( .I(n27844), .Z(n27810) );
  BUF U6631 ( .I(n27609), .Z(n27575) );
  BUF U6632 ( .I(n29254), .Z(n29221) );
  BUF U6633 ( .I(n29019), .Z(n28986) );
  BUF U6634 ( .I(n28784), .Z(n28751) );
  BUF U6635 ( .I(n28549), .Z(n28516) );
  BUF U6636 ( .I(n28314), .Z(n28281) );
  BUF U6637 ( .I(n28079), .Z(n28046) );
  BUF U6638 ( .I(n27844), .Z(n27811) );
  BUF U6639 ( .I(n27609), .Z(n27576) );
  BUF U6640 ( .I(n29253), .Z(n29222) );
  BUF U6641 ( .I(n29018), .Z(n28987) );
  BUF U6642 ( .I(n28783), .Z(n28752) );
  BUF U6643 ( .I(n28548), .Z(n28517) );
  BUF U6644 ( .I(n28313), .Z(n28282) );
  BUF U6645 ( .I(n28078), .Z(n28047) );
  BUF U6646 ( .I(n27843), .Z(n27812) );
  BUF U6647 ( .I(n27608), .Z(n27577) );
  BUF U6648 ( .I(n29253), .Z(n29223) );
  BUF U6649 ( .I(n29018), .Z(n28988) );
  BUF U6650 ( .I(n28783), .Z(n28753) );
  BUF U6651 ( .I(n28548), .Z(n28518) );
  BUF U6652 ( .I(n28313), .Z(n28283) );
  BUF U6653 ( .I(n28078), .Z(n28048) );
  BUF U6654 ( .I(n27843), .Z(n27813) );
  BUF U6655 ( .I(n27608), .Z(n27578) );
  BUF U6656 ( .I(n29253), .Z(n29224) );
  BUF U6657 ( .I(n29018), .Z(n28989) );
  BUF U6658 ( .I(n28783), .Z(n28754) );
  BUF U6659 ( .I(n28548), .Z(n28519) );
  BUF U6660 ( .I(n28313), .Z(n28284) );
  BUF U6661 ( .I(n28078), .Z(n28049) );
  BUF U6662 ( .I(n27843), .Z(n27814) );
  BUF U6663 ( .I(n27608), .Z(n27579) );
  BUF U6664 ( .I(n29252), .Z(n29225) );
  BUF U6665 ( .I(n29017), .Z(n28990) );
  BUF U6666 ( .I(n28782), .Z(n28755) );
  BUF U6667 ( .I(n28547), .Z(n28520) );
  BUF U6668 ( .I(n28312), .Z(n28285) );
  BUF U6669 ( .I(n28077), .Z(n28050) );
  BUF U6670 ( .I(n27842), .Z(n27815) );
  BUF U6671 ( .I(n27607), .Z(n27580) );
  BUF U6672 ( .I(n29252), .Z(n29226) );
  BUF U6673 ( .I(n29017), .Z(n28991) );
  BUF U6674 ( .I(n28782), .Z(n28756) );
  BUF U6675 ( .I(n28547), .Z(n28521) );
  BUF U6676 ( .I(n28312), .Z(n28286) );
  BUF U6677 ( .I(n28077), .Z(n28051) );
  BUF U6678 ( .I(n27842), .Z(n27816) );
  BUF U6679 ( .I(n27607), .Z(n27581) );
  BUF U6680 ( .I(n29252), .Z(n29227) );
  BUF U6681 ( .I(n29017), .Z(n28992) );
  BUF U6682 ( .I(n28782), .Z(n28757) );
  BUF U6683 ( .I(n28547), .Z(n28522) );
  BUF U6684 ( .I(n28312), .Z(n28287) );
  BUF U6685 ( .I(n28077), .Z(n28052) );
  BUF U6686 ( .I(n27842), .Z(n27817) );
  BUF U6687 ( .I(n27607), .Z(n27582) );
  BUF U6688 ( .I(n29251), .Z(n29228) );
  BUF U6689 ( .I(n29016), .Z(n28993) );
  BUF U6690 ( .I(n28781), .Z(n28758) );
  BUF U6691 ( .I(n28546), .Z(n28523) );
  BUF U6692 ( .I(n28311), .Z(n28288) );
  BUF U6693 ( .I(n28076), .Z(n28053) );
  BUF U6694 ( .I(n27841), .Z(n27818) );
  BUF U6695 ( .I(n27606), .Z(n27583) );
  BUF U6696 ( .I(n29251), .Z(n29229) );
  BUF U6697 ( .I(n29016), .Z(n28994) );
  BUF U6698 ( .I(n28781), .Z(n28759) );
  BUF U6699 ( .I(n28546), .Z(n28524) );
  BUF U6700 ( .I(n28311), .Z(n28289) );
  BUF U6701 ( .I(n28076), .Z(n28054) );
  BUF U6702 ( .I(n27841), .Z(n27819) );
  BUF U6703 ( .I(n27606), .Z(n27584) );
  BUF U6704 ( .I(n29251), .Z(n29230) );
  BUF U6705 ( .I(n29016), .Z(n28995) );
  BUF U6706 ( .I(n28781), .Z(n28760) );
  BUF U6707 ( .I(n28546), .Z(n28525) );
  BUF U6708 ( .I(n28311), .Z(n28290) );
  BUF U6709 ( .I(n28076), .Z(n28055) );
  BUF U6710 ( .I(n27841), .Z(n27820) );
  BUF U6711 ( .I(n27606), .Z(n27585) );
  BUF U6712 ( .I(n29250), .Z(n29231) );
  BUF U6713 ( .I(n29015), .Z(n28996) );
  BUF U6714 ( .I(n28780), .Z(n28761) );
  BUF U6715 ( .I(n28545), .Z(n28526) );
  BUF U6716 ( .I(n28310), .Z(n28291) );
  BUF U6717 ( .I(n28075), .Z(n28056) );
  BUF U6718 ( .I(n27840), .Z(n27821) );
  BUF U6719 ( .I(n27605), .Z(n27586) );
  BUF U6720 ( .I(n29250), .Z(n29232) );
  BUF U6721 ( .I(n29015), .Z(n28997) );
  BUF U6722 ( .I(n28780), .Z(n28762) );
  BUF U6723 ( .I(n28545), .Z(n28527) );
  BUF U6724 ( .I(n28310), .Z(n28292) );
  BUF U6725 ( .I(n28075), .Z(n28057) );
  BUF U6726 ( .I(n27840), .Z(n27822) );
  BUF U6727 ( .I(n27605), .Z(n27587) );
  BUF U6728 ( .I(n29250), .Z(n29233) );
  BUF U6729 ( .I(n29015), .Z(n28998) );
  BUF U6730 ( .I(n28780), .Z(n28763) );
  BUF U6731 ( .I(n28545), .Z(n28528) );
  BUF U6732 ( .I(n28310), .Z(n28293) );
  BUF U6733 ( .I(n28075), .Z(n28058) );
  BUF U6734 ( .I(n27840), .Z(n27823) );
  BUF U6735 ( .I(n27605), .Z(n27588) );
  BUF U6736 ( .I(n29249), .Z(n29234) );
  BUF U6737 ( .I(n29014), .Z(n28999) );
  BUF U6738 ( .I(n28779), .Z(n28764) );
  BUF U6739 ( .I(n28544), .Z(n28529) );
  BUF U6740 ( .I(n28309), .Z(n28294) );
  BUF U6741 ( .I(n28074), .Z(n28059) );
  BUF U6742 ( .I(n27839), .Z(n27824) );
  BUF U6743 ( .I(n27604), .Z(n27589) );
  BUF U6744 ( .I(n29249), .Z(n29235) );
  BUF U6745 ( .I(n29014), .Z(n29000) );
  BUF U6746 ( .I(n28779), .Z(n28765) );
  BUF U6747 ( .I(n28544), .Z(n28530) );
  BUF U6748 ( .I(n28309), .Z(n28295) );
  BUF U6749 ( .I(n28074), .Z(n28060) );
  BUF U6750 ( .I(n27839), .Z(n27825) );
  BUF U6751 ( .I(n27604), .Z(n27590) );
  BUF U6752 ( .I(n29249), .Z(n29236) );
  BUF U6753 ( .I(n29014), .Z(n29001) );
  BUF U6754 ( .I(n28779), .Z(n28766) );
  BUF U6755 ( .I(n28544), .Z(n28531) );
  BUF U6756 ( .I(n28309), .Z(n28296) );
  BUF U6757 ( .I(n28074), .Z(n28061) );
  BUF U6758 ( .I(n27839), .Z(n27826) );
  BUF U6759 ( .I(n27604), .Z(n27591) );
  BUF U6760 ( .I(n29248), .Z(n29237) );
  BUF U6761 ( .I(n29013), .Z(n29002) );
  BUF U6762 ( .I(n28778), .Z(n28767) );
  BUF U6763 ( .I(n28543), .Z(n28532) );
  BUF U6764 ( .I(n28308), .Z(n28297) );
  BUF U6765 ( .I(n28073), .Z(n28062) );
  BUF U6766 ( .I(n27838), .Z(n27827) );
  BUF U6767 ( .I(n27603), .Z(n27592) );
  BUF U6768 ( .I(n29248), .Z(n29238) );
  BUF U6769 ( .I(n29013), .Z(n29003) );
  BUF U6770 ( .I(n28778), .Z(n28768) );
  BUF U6771 ( .I(n28543), .Z(n28533) );
  BUF U6772 ( .I(n28308), .Z(n28298) );
  BUF U6773 ( .I(n28073), .Z(n28063) );
  BUF U6774 ( .I(n27838), .Z(n27828) );
  BUF U6775 ( .I(n27603), .Z(n27593) );
  BUF U6776 ( .I(n29248), .Z(n29239) );
  BUF U6777 ( .I(n29013), .Z(n29004) );
  BUF U6778 ( .I(n28778), .Z(n28769) );
  BUF U6779 ( .I(n28543), .Z(n28534) );
  BUF U6780 ( .I(n28308), .Z(n28299) );
  BUF U6781 ( .I(n28073), .Z(n28064) );
  BUF U6782 ( .I(n27838), .Z(n27829) );
  BUF U6783 ( .I(n27603), .Z(n27594) );
  BUF U6784 ( .I(n29247), .Z(n29240) );
  BUF U6785 ( .I(n29012), .Z(n29005) );
  BUF U6786 ( .I(n28777), .Z(n28770) );
  BUF U6787 ( .I(n28542), .Z(n28535) );
  BUF U6788 ( .I(n28307), .Z(n28300) );
  BUF U6789 ( .I(n28072), .Z(n28065) );
  BUF U6790 ( .I(n27837), .Z(n27830) );
  BUF U6791 ( .I(n27602), .Z(n27595) );
  BUF U6792 ( .I(n29247), .Z(n29241) );
  BUF U6793 ( .I(n29012), .Z(n29006) );
  BUF U6794 ( .I(n28777), .Z(n28771) );
  BUF U6795 ( .I(n28542), .Z(n28536) );
  BUF U6796 ( .I(n28307), .Z(n28301) );
  BUF U6797 ( .I(n28072), .Z(n28066) );
  BUF U6798 ( .I(n27837), .Z(n27831) );
  BUF U6799 ( .I(n27602), .Z(n27596) );
  BUF U6800 ( .I(n29247), .Z(n29242) );
  BUF U6801 ( .I(n29012), .Z(n29007) );
  BUF U6802 ( .I(n28777), .Z(n28772) );
  BUF U6803 ( .I(n28542), .Z(n28537) );
  BUF U6804 ( .I(n28307), .Z(n28302) );
  BUF U6805 ( .I(n28072), .Z(n28067) );
  BUF U6806 ( .I(n27837), .Z(n27832) );
  BUF U6807 ( .I(n27602), .Z(n27597) );
  BUF U6808 ( .I(n29246), .Z(n29243) );
  BUF U6809 ( .I(n29011), .Z(n29008) );
  BUF U6810 ( .I(n28776), .Z(n28773) );
  BUF U6811 ( .I(n28541), .Z(n28538) );
  BUF U6812 ( .I(n28306), .Z(n28303) );
  BUF U6813 ( .I(n28071), .Z(n28068) );
  BUF U6814 ( .I(n27836), .Z(n27833) );
  BUF U6815 ( .I(n27601), .Z(n27598) );
  BUF U6816 ( .I(n29246), .Z(n29244) );
  BUF U6817 ( .I(n29011), .Z(n29009) );
  BUF U6818 ( .I(n28776), .Z(n28774) );
  BUF U6819 ( .I(n28541), .Z(n28539) );
  BUF U6820 ( .I(n28306), .Z(n28304) );
  BUF U6821 ( .I(n28071), .Z(n28069) );
  BUF U6822 ( .I(n27836), .Z(n27834) );
  BUF U6823 ( .I(n27601), .Z(n27599) );
  BUF U6824 ( .I(n29246), .Z(n29245) );
  BUF U6825 ( .I(n29011), .Z(n29010) );
  BUF U6826 ( .I(n28776), .Z(n28775) );
  BUF U6827 ( .I(n28541), .Z(n28540) );
  BUF U6828 ( .I(n28306), .Z(n28305) );
  BUF U6829 ( .I(n28071), .Z(n28070) );
  BUF U6830 ( .I(n27836), .Z(n27835) );
  BUF U6831 ( .I(n27601), .Z(n27600) );
  BUF U6832 ( .I(n29579), .Z(n29576) );
  BUF U6833 ( .I(n29579), .Z(n29577) );
  BUF U6834 ( .I(n29580), .Z(n29575) );
  BUF U6835 ( .I(n29580), .Z(n29573) );
  BUF U6836 ( .I(n29580), .Z(n29574) );
  BUF U6837 ( .I(n29572), .Z(n29569) );
  BUF U6838 ( .I(n29572), .Z(n29570) );
  BUF U6839 ( .I(n29579), .Z(n29578) );
  BUF U6840 ( .I(n26882), .Z(n27023) );
  BUF U6841 ( .I(n26881), .Z(n26882) );
  BUF U6842 ( .I(n26867), .Z(n26878) );
  BUF U6843 ( .I(n26392), .Z(n26403) );
  BUF U6844 ( .I(n26867), .Z(n26877) );
  BUF U6845 ( .I(n26392), .Z(n26402) );
  BUF U6846 ( .I(n26868), .Z(n26875) );
  BUF U6847 ( .I(n26393), .Z(n26400) );
  BUF U6848 ( .I(n26868), .Z(n26874) );
  BUF U6849 ( .I(n26393), .Z(n26399) );
  BUF U6850 ( .I(n26869), .Z(n26871) );
  BUF U6851 ( .I(n26394), .Z(n26396) );
  BUF U6852 ( .I(n26881), .Z(n26883) );
  BUF U6853 ( .I(n26879), .Z(n26888) );
  BUF U6854 ( .I(n26880), .Z(n26887) );
  BUF U6855 ( .I(n26867), .Z(n26876) );
  BUF U6856 ( .I(n26392), .Z(n26401) );
  BUF U6857 ( .I(n26868), .Z(n26873) );
  BUF U6858 ( .I(n26393), .Z(n26398) );
  BUF U6859 ( .I(n26869), .Z(n26872) );
  BUF U6860 ( .I(n26394), .Z(n26397) );
  BUF U6861 ( .I(n26869), .Z(n26870) );
  BUF U6862 ( .I(n26394), .Z(n26395) );
  BUF U6863 ( .I(n26880), .Z(n26886) );
  BUF U6864 ( .I(n26405), .Z(n26411) );
  BUF U6865 ( .I(n26881), .Z(n26884) );
  BUF U6866 ( .I(n26880), .Z(n26885) );
  BUF U6867 ( .I(n26879), .Z(n26890) );
  BUF U6868 ( .I(n26404), .Z(n26415) );
  BUF U6869 ( .I(n26879), .Z(n26889) );
  BUF U6870 ( .I(n26167), .Z(n26272) );
  BUF U6871 ( .I(n26166), .Z(n26167) );
  BUF U6872 ( .I(n26285), .Z(n26390) );
  BUF U6873 ( .I(n26284), .Z(n26285) );
  BUF U6874 ( .I(n26407), .Z(n26548) );
  BUF U6875 ( .I(n26406), .Z(n26407) );
  BUF U6876 ( .I(n26406), .Z(n26408) );
  BUF U6877 ( .I(n26404), .Z(n26413) );
  BUF U6878 ( .I(n26405), .Z(n26412) );
  BUF U6879 ( .I(n26406), .Z(n26409) );
  BUF U6880 ( .I(n26405), .Z(n26410) );
  BUF U6881 ( .I(n26404), .Z(n26414) );
  BUF U6882 ( .I(n26158), .Z(n26193) );
  BUF U6883 ( .I(n26276), .Z(n26311) );
  BUF U6884 ( .I(n26159), .Z(n26190) );
  BUF U6885 ( .I(n26277), .Z(n26308) );
  BUF U6886 ( .I(n26160), .Z(n26186) );
  BUF U6887 ( .I(n26278), .Z(n26304) );
  BUF U6888 ( .I(n26160), .Z(n26187) );
  BUF U6889 ( .I(n26278), .Z(n26305) );
  BUF U6890 ( .I(n26161), .Z(n26183) );
  BUF U6891 ( .I(n26279), .Z(n26301) );
  BUF U6892 ( .I(n26162), .Z(n26180) );
  BUF U6893 ( .I(n26280), .Z(n26298) );
  BUF U6894 ( .I(n26163), .Z(n26177) );
  BUF U6895 ( .I(n26281), .Z(n26295) );
  BUF U6896 ( .I(n26164), .Z(n26173) );
  BUF U6897 ( .I(n26282), .Z(n26291) );
  BUF U6898 ( .I(n26165), .Z(n26170) );
  BUF U6899 ( .I(n26283), .Z(n26288) );
  BUF U6900 ( .I(n26158), .Z(n26191) );
  BUF U6901 ( .I(n26276), .Z(n26309) );
  BUF U6902 ( .I(n26158), .Z(n26192) );
  BUF U6903 ( .I(n26276), .Z(n26310) );
  BUF U6904 ( .I(n26159), .Z(n26189) );
  BUF U6905 ( .I(n26277), .Z(n26307) );
  BUF U6906 ( .I(n26159), .Z(n26188) );
  BUF U6907 ( .I(n26277), .Z(n26306) );
  BUF U6908 ( .I(n26161), .Z(n26184) );
  BUF U6909 ( .I(n26279), .Z(n26302) );
  BUF U6910 ( .I(n26160), .Z(n26185) );
  BUF U6911 ( .I(n26278), .Z(n26303) );
  BUF U6912 ( .I(n26162), .Z(n26181) );
  BUF U6913 ( .I(n26280), .Z(n26299) );
  BUF U6914 ( .I(n26161), .Z(n26182) );
  BUF U6915 ( .I(n26279), .Z(n26300) );
  BUF U6916 ( .I(n26163), .Z(n26178) );
  BUF U6917 ( .I(n26281), .Z(n26296) );
  BUF U6918 ( .I(n26162), .Z(n26179) );
  BUF U6919 ( .I(n26280), .Z(n26297) );
  BUF U6920 ( .I(n26164), .Z(n26174) );
  BUF U6921 ( .I(n26282), .Z(n26292) );
  BUF U6922 ( .I(n26163), .Z(n26176) );
  BUF U6923 ( .I(n26281), .Z(n26294) );
  BUF U6924 ( .I(n26164), .Z(n26175) );
  BUF U6925 ( .I(n26282), .Z(n26293) );
  BUF U6926 ( .I(n26165), .Z(n26171) );
  BUF U6927 ( .I(n26283), .Z(n26289) );
  BUF U6928 ( .I(n26165), .Z(n26172) );
  BUF U6929 ( .I(n26283), .Z(n26290) );
  BUF U6930 ( .I(n26166), .Z(n26168) );
  BUF U6931 ( .I(n26284), .Z(n26286) );
  BUF U6932 ( .I(n26166), .Z(n26169) );
  BUF U6933 ( .I(n26284), .Z(n26287) );
  AND2 U6934 ( .A1(n4099), .A2(n4100), .Z(n23) );
  BUF U6935 ( .I(n26103), .Z(n26108) );
  BUF U6936 ( .I(n26103), .Z(n26109) );
  BUF U6937 ( .I(n26103), .Z(n26110) );
  BUF U6938 ( .I(n26102), .Z(n26112) );
  BUF U6939 ( .I(n26102), .Z(n26111) );
  BUF U6940 ( .I(n26102), .Z(n26113) );
  BUF U6941 ( .I(n26101), .Z(n26114) );
  BUF U6942 ( .I(n26100), .Z(n26117) );
  BUF U6943 ( .I(n26101), .Z(n26115) );
  BUF U6944 ( .I(n26101), .Z(n26116) );
  BUF U6945 ( .I(n26100), .Z(n26119) );
  BUF U6946 ( .I(n26100), .Z(n26118) );
  BUF U6947 ( .I(n26099), .Z(n26122) );
  BUF U6948 ( .I(n26099), .Z(n26120) );
  BUF U6949 ( .I(n26099), .Z(n26121) );
  BUF U6950 ( .I(n26098), .Z(n26124) );
  BUF U6951 ( .I(n26098), .Z(n26123) );
  BUF U6952 ( .I(n26128), .Z(n26154) );
  BUF U6953 ( .I(n26128), .Z(n26153) );
  BUF U6954 ( .I(n26133), .Z(n26138) );
  BUF U6955 ( .I(n26133), .Z(n26139) );
  BUF U6956 ( .I(n26133), .Z(n26140) );
  BUF U6957 ( .I(n26132), .Z(n26142) );
  BUF U6958 ( .I(n26132), .Z(n26141) );
  BUF U6959 ( .I(n26132), .Z(n26143) );
  BUF U6960 ( .I(n26131), .Z(n26144) );
  BUF U6961 ( .I(n26130), .Z(n26147) );
  BUF U6962 ( .I(n26131), .Z(n26145) );
  BUF U6963 ( .I(n26131), .Z(n26146) );
  BUF U6964 ( .I(n26130), .Z(n26149) );
  BUF U6965 ( .I(n26130), .Z(n26148) );
  BUF U6966 ( .I(n26129), .Z(n26152) );
  BUF U6967 ( .I(n26129), .Z(n26150) );
  BUF U6968 ( .I(n26129), .Z(n26151) );
  BUF U6969 ( .I(n29316), .Z(n29247) );
  BUF U6970 ( .I(n29081), .Z(n29012) );
  BUF U6971 ( .I(n28846), .Z(n28777) );
  BUF U6972 ( .I(n28611), .Z(n28542) );
  BUF U6973 ( .I(n28376), .Z(n28307) );
  BUF U6974 ( .I(n28141), .Z(n28072) );
  BUF U6975 ( .I(n27906), .Z(n27837) );
  BUF U6976 ( .I(n27671), .Z(n27602) );
  BUF U6977 ( .I(n29316), .Z(n29246) );
  BUF U6978 ( .I(n29081), .Z(n29011) );
  BUF U6979 ( .I(n28846), .Z(n28776) );
  BUF U6980 ( .I(n28611), .Z(n28541) );
  BUF U6981 ( .I(n28376), .Z(n28306) );
  BUF U6982 ( .I(n28141), .Z(n28071) );
  BUF U6983 ( .I(n27906), .Z(n27836) );
  BUF U6984 ( .I(n27671), .Z(n27601) );
  BUF U6985 ( .I(n29299), .Z(n29297) );
  BUF U6986 ( .I(n29064), .Z(n29062) );
  BUF U6987 ( .I(n28829), .Z(n28827) );
  BUF U6988 ( .I(n28594), .Z(n28592) );
  BUF U6989 ( .I(n28359), .Z(n28357) );
  BUF U6990 ( .I(n28124), .Z(n28122) );
  BUF U6991 ( .I(n27889), .Z(n27887) );
  BUF U6992 ( .I(n27654), .Z(n27652) );
  BUF U6993 ( .I(n29299), .Z(n29296) );
  BUF U6994 ( .I(n29064), .Z(n29061) );
  BUF U6995 ( .I(n28829), .Z(n28826) );
  BUF U6996 ( .I(n28594), .Z(n28591) );
  BUF U6997 ( .I(n28359), .Z(n28356) );
  BUF U6998 ( .I(n28124), .Z(n28121) );
  BUF U6999 ( .I(n27889), .Z(n27886) );
  BUF U7000 ( .I(n27654), .Z(n27651) );
  BUF U7001 ( .I(n29300), .Z(n29295) );
  BUF U7002 ( .I(n29065), .Z(n29060) );
  BUF U7003 ( .I(n28830), .Z(n28825) );
  BUF U7004 ( .I(n28595), .Z(n28590) );
  BUF U7005 ( .I(n28360), .Z(n28355) );
  BUF U7006 ( .I(n28125), .Z(n28120) );
  BUF U7007 ( .I(n27890), .Z(n27885) );
  BUF U7008 ( .I(n27655), .Z(n27650) );
  BUF U7009 ( .I(n29300), .Z(n29294) );
  BUF U7010 ( .I(n29065), .Z(n29059) );
  BUF U7011 ( .I(n28830), .Z(n28824) );
  BUF U7012 ( .I(n28595), .Z(n28589) );
  BUF U7013 ( .I(n28360), .Z(n28354) );
  BUF U7014 ( .I(n28125), .Z(n28119) );
  BUF U7015 ( .I(n27890), .Z(n27884) );
  BUF U7016 ( .I(n27655), .Z(n27649) );
  BUF U7017 ( .I(n29300), .Z(n29293) );
  BUF U7018 ( .I(n29065), .Z(n29058) );
  BUF U7019 ( .I(n28830), .Z(n28823) );
  BUF U7020 ( .I(n28595), .Z(n28588) );
  BUF U7021 ( .I(n28360), .Z(n28353) );
  BUF U7022 ( .I(n28125), .Z(n28118) );
  BUF U7023 ( .I(n27890), .Z(n27883) );
  BUF U7024 ( .I(n27655), .Z(n27648) );
  BUF U7025 ( .I(n29301), .Z(n29292) );
  BUF U7026 ( .I(n29066), .Z(n29057) );
  BUF U7027 ( .I(n28831), .Z(n28822) );
  BUF U7028 ( .I(n28596), .Z(n28587) );
  BUF U7029 ( .I(n28361), .Z(n28352) );
  BUF U7030 ( .I(n28126), .Z(n28117) );
  BUF U7031 ( .I(n27891), .Z(n27882) );
  BUF U7032 ( .I(n27656), .Z(n27647) );
  BUF U7033 ( .I(n29301), .Z(n29291) );
  BUF U7034 ( .I(n29066), .Z(n29056) );
  BUF U7035 ( .I(n28831), .Z(n28821) );
  BUF U7036 ( .I(n28596), .Z(n28586) );
  BUF U7037 ( .I(n28361), .Z(n28351) );
  BUF U7038 ( .I(n28126), .Z(n28116) );
  BUF U7039 ( .I(n27891), .Z(n27881) );
  BUF U7040 ( .I(n27656), .Z(n27646) );
  BUF U7041 ( .I(n29301), .Z(n29290) );
  BUF U7042 ( .I(n29066), .Z(n29055) );
  BUF U7043 ( .I(n28831), .Z(n28820) );
  BUF U7044 ( .I(n28596), .Z(n28585) );
  BUF U7045 ( .I(n28361), .Z(n28350) );
  BUF U7046 ( .I(n28126), .Z(n28115) );
  BUF U7047 ( .I(n27891), .Z(n27880) );
  BUF U7048 ( .I(n27656), .Z(n27645) );
  BUF U7049 ( .I(n29302), .Z(n29289) );
  BUF U7050 ( .I(n29067), .Z(n29054) );
  BUF U7051 ( .I(n28832), .Z(n28819) );
  BUF U7052 ( .I(n28597), .Z(n28584) );
  BUF U7053 ( .I(n28362), .Z(n28349) );
  BUF U7054 ( .I(n28127), .Z(n28114) );
  BUF U7055 ( .I(n27892), .Z(n27879) );
  BUF U7056 ( .I(n27657), .Z(n27644) );
  BUF U7057 ( .I(n29302), .Z(n29288) );
  BUF U7058 ( .I(n29067), .Z(n29053) );
  BUF U7059 ( .I(n28832), .Z(n28818) );
  BUF U7060 ( .I(n28597), .Z(n28583) );
  BUF U7061 ( .I(n28362), .Z(n28348) );
  BUF U7062 ( .I(n28127), .Z(n28113) );
  BUF U7063 ( .I(n27892), .Z(n27878) );
  BUF U7064 ( .I(n27657), .Z(n27643) );
  BUF U7065 ( .I(n29302), .Z(n29287) );
  BUF U7066 ( .I(n29067), .Z(n29052) );
  BUF U7067 ( .I(n28832), .Z(n28817) );
  BUF U7068 ( .I(n28597), .Z(n28582) );
  BUF U7069 ( .I(n28362), .Z(n28347) );
  BUF U7070 ( .I(n28127), .Z(n28112) );
  BUF U7071 ( .I(n27892), .Z(n27877) );
  BUF U7072 ( .I(n27657), .Z(n27642) );
  BUF U7073 ( .I(n29303), .Z(n29286) );
  BUF U7074 ( .I(n29068), .Z(n29051) );
  BUF U7075 ( .I(n28833), .Z(n28816) );
  BUF U7076 ( .I(n28598), .Z(n28581) );
  BUF U7077 ( .I(n28363), .Z(n28346) );
  BUF U7078 ( .I(n28128), .Z(n28111) );
  BUF U7079 ( .I(n27893), .Z(n27876) );
  BUF U7080 ( .I(n27658), .Z(n27641) );
  BUF U7081 ( .I(n29303), .Z(n29285) );
  BUF U7082 ( .I(n29068), .Z(n29050) );
  BUF U7083 ( .I(n28833), .Z(n28815) );
  BUF U7084 ( .I(n28598), .Z(n28580) );
  BUF U7085 ( .I(n28363), .Z(n28345) );
  BUF U7086 ( .I(n28128), .Z(n28110) );
  BUF U7087 ( .I(n27893), .Z(n27875) );
  BUF U7088 ( .I(n27658), .Z(n27640) );
  BUF U7089 ( .I(n29303), .Z(n29284) );
  BUF U7090 ( .I(n29068), .Z(n29049) );
  BUF U7091 ( .I(n28833), .Z(n28814) );
  BUF U7092 ( .I(n28598), .Z(n28579) );
  BUF U7093 ( .I(n28363), .Z(n28344) );
  BUF U7094 ( .I(n28128), .Z(n28109) );
  BUF U7095 ( .I(n27893), .Z(n27874) );
  BUF U7096 ( .I(n27658), .Z(n27639) );
  BUF U7097 ( .I(n29304), .Z(n29283) );
  BUF U7098 ( .I(n29069), .Z(n29048) );
  BUF U7099 ( .I(n28834), .Z(n28813) );
  BUF U7100 ( .I(n28599), .Z(n28578) );
  BUF U7101 ( .I(n28364), .Z(n28343) );
  BUF U7102 ( .I(n28129), .Z(n28108) );
  BUF U7103 ( .I(n27894), .Z(n27873) );
  BUF U7104 ( .I(n27659), .Z(n27638) );
  BUF U7105 ( .I(n29304), .Z(n29282) );
  BUF U7106 ( .I(n29069), .Z(n29047) );
  BUF U7107 ( .I(n28834), .Z(n28812) );
  BUF U7108 ( .I(n28599), .Z(n28577) );
  BUF U7109 ( .I(n28364), .Z(n28342) );
  BUF U7110 ( .I(n28129), .Z(n28107) );
  BUF U7111 ( .I(n27894), .Z(n27872) );
  BUF U7112 ( .I(n27659), .Z(n27637) );
  BUF U7113 ( .I(n29304), .Z(n29281) );
  BUF U7114 ( .I(n29069), .Z(n29046) );
  BUF U7115 ( .I(n28834), .Z(n28811) );
  BUF U7116 ( .I(n28599), .Z(n28576) );
  BUF U7117 ( .I(n28364), .Z(n28341) );
  BUF U7118 ( .I(n28129), .Z(n28106) );
  BUF U7119 ( .I(n27894), .Z(n27871) );
  BUF U7120 ( .I(n27659), .Z(n27636) );
  BUF U7121 ( .I(n29305), .Z(n29280) );
  BUF U7122 ( .I(n29070), .Z(n29045) );
  BUF U7123 ( .I(n28835), .Z(n28810) );
  BUF U7124 ( .I(n28600), .Z(n28575) );
  BUF U7125 ( .I(n28365), .Z(n28340) );
  BUF U7126 ( .I(n28130), .Z(n28105) );
  BUF U7127 ( .I(n27895), .Z(n27870) );
  BUF U7128 ( .I(n27660), .Z(n27635) );
  BUF U7129 ( .I(n29305), .Z(n29279) );
  BUF U7130 ( .I(n29070), .Z(n29044) );
  BUF U7131 ( .I(n28835), .Z(n28809) );
  BUF U7132 ( .I(n28600), .Z(n28574) );
  BUF U7133 ( .I(n28365), .Z(n28339) );
  BUF U7134 ( .I(n28130), .Z(n28104) );
  BUF U7135 ( .I(n27895), .Z(n27869) );
  BUF U7136 ( .I(n27660), .Z(n27634) );
  BUF U7137 ( .I(n29305), .Z(n29278) );
  BUF U7138 ( .I(n29070), .Z(n29043) );
  BUF U7139 ( .I(n28835), .Z(n28808) );
  BUF U7140 ( .I(n28600), .Z(n28573) );
  BUF U7141 ( .I(n28365), .Z(n28338) );
  BUF U7142 ( .I(n28130), .Z(n28103) );
  BUF U7143 ( .I(n27895), .Z(n27868) );
  BUF U7144 ( .I(n27660), .Z(n27633) );
  BUF U7145 ( .I(n29306), .Z(n29277) );
  BUF U7146 ( .I(n29071), .Z(n29042) );
  BUF U7147 ( .I(n28836), .Z(n28807) );
  BUF U7148 ( .I(n28601), .Z(n28572) );
  BUF U7149 ( .I(n28366), .Z(n28337) );
  BUF U7150 ( .I(n28131), .Z(n28102) );
  BUF U7151 ( .I(n27896), .Z(n27867) );
  BUF U7152 ( .I(n27661), .Z(n27632) );
  BUF U7153 ( .I(n29306), .Z(n29276) );
  BUF U7154 ( .I(n29071), .Z(n29041) );
  BUF U7155 ( .I(n28836), .Z(n28806) );
  BUF U7156 ( .I(n28601), .Z(n28571) );
  BUF U7157 ( .I(n28366), .Z(n28336) );
  BUF U7158 ( .I(n28131), .Z(n28101) );
  BUF U7159 ( .I(n27896), .Z(n27866) );
  BUF U7160 ( .I(n27661), .Z(n27631) );
  BUF U7161 ( .I(n29306), .Z(n29275) );
  BUF U7162 ( .I(n29071), .Z(n29040) );
  BUF U7163 ( .I(n28836), .Z(n28805) );
  BUF U7164 ( .I(n28601), .Z(n28570) );
  BUF U7165 ( .I(n28366), .Z(n28335) );
  BUF U7166 ( .I(n28131), .Z(n28100) );
  BUF U7167 ( .I(n27896), .Z(n27865) );
  BUF U7168 ( .I(n27661), .Z(n27630) );
  BUF U7169 ( .I(n29307), .Z(n29274) );
  BUF U7170 ( .I(n29072), .Z(n29039) );
  BUF U7171 ( .I(n28837), .Z(n28804) );
  BUF U7172 ( .I(n28602), .Z(n28569) );
  BUF U7173 ( .I(n28367), .Z(n28334) );
  BUF U7174 ( .I(n28132), .Z(n28099) );
  BUF U7175 ( .I(n27897), .Z(n27864) );
  BUF U7176 ( .I(n27662), .Z(n27629) );
  BUF U7177 ( .I(n29307), .Z(n29273) );
  BUF U7178 ( .I(n29072), .Z(n29038) );
  BUF U7179 ( .I(n28837), .Z(n28803) );
  BUF U7180 ( .I(n28602), .Z(n28568) );
  BUF U7181 ( .I(n28367), .Z(n28333) );
  BUF U7182 ( .I(n28132), .Z(n28098) );
  BUF U7183 ( .I(n27897), .Z(n27863) );
  BUF U7184 ( .I(n27662), .Z(n27628) );
  BUF U7185 ( .I(n29307), .Z(n29272) );
  BUF U7186 ( .I(n29072), .Z(n29037) );
  BUF U7187 ( .I(n28837), .Z(n28802) );
  BUF U7188 ( .I(n28602), .Z(n28567) );
  BUF U7189 ( .I(n28367), .Z(n28332) );
  BUF U7190 ( .I(n28132), .Z(n28097) );
  BUF U7191 ( .I(n27897), .Z(n27862) );
  BUF U7192 ( .I(n27662), .Z(n27627) );
  BUF U7193 ( .I(n29308), .Z(n29271) );
  BUF U7194 ( .I(n29073), .Z(n29036) );
  BUF U7195 ( .I(n28838), .Z(n28801) );
  BUF U7196 ( .I(n28603), .Z(n28566) );
  BUF U7197 ( .I(n28368), .Z(n28331) );
  BUF U7198 ( .I(n28133), .Z(n28096) );
  BUF U7199 ( .I(n27898), .Z(n27861) );
  BUF U7200 ( .I(n27663), .Z(n27626) );
  BUF U7201 ( .I(n29308), .Z(n29270) );
  BUF U7202 ( .I(n29073), .Z(n29035) );
  BUF U7203 ( .I(n28838), .Z(n28800) );
  BUF U7204 ( .I(n28603), .Z(n28565) );
  BUF U7205 ( .I(n28368), .Z(n28330) );
  BUF U7206 ( .I(n28133), .Z(n28095) );
  BUF U7207 ( .I(n27898), .Z(n27860) );
  BUF U7208 ( .I(n27663), .Z(n27625) );
  BUF U7209 ( .I(n29308), .Z(n29269) );
  BUF U7210 ( .I(n29073), .Z(n29034) );
  BUF U7211 ( .I(n28838), .Z(n28799) );
  BUF U7212 ( .I(n28603), .Z(n28564) );
  BUF U7213 ( .I(n28368), .Z(n28329) );
  BUF U7214 ( .I(n28133), .Z(n28094) );
  BUF U7215 ( .I(n27898), .Z(n27859) );
  BUF U7216 ( .I(n27663), .Z(n27624) );
  BUF U7217 ( .I(n29309), .Z(n29268) );
  BUF U7218 ( .I(n29074), .Z(n29033) );
  BUF U7219 ( .I(n28839), .Z(n28798) );
  BUF U7220 ( .I(n28604), .Z(n28563) );
  BUF U7221 ( .I(n28369), .Z(n28328) );
  BUF U7222 ( .I(n28134), .Z(n28093) );
  BUF U7223 ( .I(n27899), .Z(n27858) );
  BUF U7224 ( .I(n27664), .Z(n27623) );
  BUF U7225 ( .I(n29309), .Z(n29267) );
  BUF U7226 ( .I(n29074), .Z(n29032) );
  BUF U7227 ( .I(n28839), .Z(n28797) );
  BUF U7228 ( .I(n28604), .Z(n28562) );
  BUF U7229 ( .I(n28369), .Z(n28327) );
  BUF U7230 ( .I(n28134), .Z(n28092) );
  BUF U7231 ( .I(n27899), .Z(n27857) );
  BUF U7232 ( .I(n27664), .Z(n27622) );
  BUF U7233 ( .I(n29309), .Z(n29266) );
  BUF U7234 ( .I(n29074), .Z(n29031) );
  BUF U7235 ( .I(n28839), .Z(n28796) );
  BUF U7236 ( .I(n28604), .Z(n28561) );
  BUF U7237 ( .I(n28369), .Z(n28326) );
  BUF U7238 ( .I(n28134), .Z(n28091) );
  BUF U7239 ( .I(n27899), .Z(n27856) );
  BUF U7240 ( .I(n27664), .Z(n27621) );
  BUF U7241 ( .I(n29310), .Z(n29265) );
  BUF U7242 ( .I(n29075), .Z(n29030) );
  BUF U7243 ( .I(n28840), .Z(n28795) );
  BUF U7244 ( .I(n28605), .Z(n28560) );
  BUF U7245 ( .I(n28370), .Z(n28325) );
  BUF U7246 ( .I(n28135), .Z(n28090) );
  BUF U7247 ( .I(n27900), .Z(n27855) );
  BUF U7248 ( .I(n27665), .Z(n27620) );
  BUF U7249 ( .I(n29310), .Z(n29264) );
  BUF U7250 ( .I(n29075), .Z(n29029) );
  BUF U7251 ( .I(n28840), .Z(n28794) );
  BUF U7252 ( .I(n28605), .Z(n28559) );
  BUF U7253 ( .I(n28370), .Z(n28324) );
  BUF U7254 ( .I(n28135), .Z(n28089) );
  BUF U7255 ( .I(n27900), .Z(n27854) );
  BUF U7256 ( .I(n27665), .Z(n27619) );
  BUF U7257 ( .I(n29310), .Z(n29263) );
  BUF U7258 ( .I(n29075), .Z(n29028) );
  BUF U7259 ( .I(n28840), .Z(n28793) );
  BUF U7260 ( .I(n28605), .Z(n28558) );
  BUF U7261 ( .I(n28370), .Z(n28323) );
  BUF U7262 ( .I(n28135), .Z(n28088) );
  BUF U7263 ( .I(n27900), .Z(n27853) );
  BUF U7264 ( .I(n27665), .Z(n27618) );
  BUF U7265 ( .I(n29311), .Z(n29262) );
  BUF U7266 ( .I(n29076), .Z(n29027) );
  BUF U7267 ( .I(n28841), .Z(n28792) );
  BUF U7268 ( .I(n28606), .Z(n28557) );
  BUF U7269 ( .I(n28371), .Z(n28322) );
  BUF U7270 ( .I(n28136), .Z(n28087) );
  BUF U7271 ( .I(n27901), .Z(n27852) );
  BUF U7272 ( .I(n27666), .Z(n27617) );
  BUF U7273 ( .I(n29311), .Z(n29261) );
  BUF U7274 ( .I(n29076), .Z(n29026) );
  BUF U7275 ( .I(n28841), .Z(n28791) );
  BUF U7276 ( .I(n28606), .Z(n28556) );
  BUF U7277 ( .I(n28371), .Z(n28321) );
  BUF U7278 ( .I(n28136), .Z(n28086) );
  BUF U7279 ( .I(n27901), .Z(n27851) );
  BUF U7280 ( .I(n27666), .Z(n27616) );
  BUF U7281 ( .I(n29311), .Z(n29260) );
  BUF U7282 ( .I(n29076), .Z(n29025) );
  BUF U7283 ( .I(n28841), .Z(n28790) );
  BUF U7284 ( .I(n28606), .Z(n28555) );
  BUF U7285 ( .I(n28371), .Z(n28320) );
  BUF U7286 ( .I(n28136), .Z(n28085) );
  BUF U7287 ( .I(n27901), .Z(n27850) );
  BUF U7288 ( .I(n27666), .Z(n27615) );
  BUF U7289 ( .I(n29312), .Z(n29259) );
  BUF U7290 ( .I(n29077), .Z(n29024) );
  BUF U7291 ( .I(n28842), .Z(n28789) );
  BUF U7292 ( .I(n28607), .Z(n28554) );
  BUF U7293 ( .I(n28372), .Z(n28319) );
  BUF U7294 ( .I(n28137), .Z(n28084) );
  BUF U7295 ( .I(n27902), .Z(n27849) );
  BUF U7296 ( .I(n27667), .Z(n27614) );
  BUF U7297 ( .I(n29312), .Z(n29258) );
  BUF U7298 ( .I(n29077), .Z(n29023) );
  BUF U7299 ( .I(n28842), .Z(n28788) );
  BUF U7300 ( .I(n28607), .Z(n28553) );
  BUF U7301 ( .I(n28372), .Z(n28318) );
  BUF U7302 ( .I(n28137), .Z(n28083) );
  BUF U7303 ( .I(n27902), .Z(n27848) );
  BUF U7304 ( .I(n27667), .Z(n27613) );
  BUF U7305 ( .I(n29312), .Z(n29257) );
  BUF U7306 ( .I(n29077), .Z(n29022) );
  BUF U7307 ( .I(n28842), .Z(n28787) );
  BUF U7308 ( .I(n28607), .Z(n28552) );
  BUF U7309 ( .I(n28372), .Z(n28317) );
  BUF U7310 ( .I(n28137), .Z(n28082) );
  BUF U7311 ( .I(n27902), .Z(n27847) );
  BUF U7312 ( .I(n27667), .Z(n27612) );
  BUF U7313 ( .I(n29313), .Z(n29256) );
  BUF U7314 ( .I(n29078), .Z(n29021) );
  BUF U7315 ( .I(n28843), .Z(n28786) );
  BUF U7316 ( .I(n28608), .Z(n28551) );
  BUF U7317 ( .I(n28373), .Z(n28316) );
  BUF U7318 ( .I(n28138), .Z(n28081) );
  BUF U7319 ( .I(n27903), .Z(n27846) );
  BUF U7320 ( .I(n27668), .Z(n27611) );
  BUF U7321 ( .I(n29313), .Z(n29255) );
  BUF U7322 ( .I(n29078), .Z(n29020) );
  BUF U7323 ( .I(n28843), .Z(n28785) );
  BUF U7324 ( .I(n28608), .Z(n28550) );
  BUF U7325 ( .I(n28373), .Z(n28315) );
  BUF U7326 ( .I(n28138), .Z(n28080) );
  BUF U7327 ( .I(n27903), .Z(n27845) );
  BUF U7328 ( .I(n27668), .Z(n27610) );
  BUF U7329 ( .I(n29313), .Z(n29254) );
  BUF U7330 ( .I(n29078), .Z(n29019) );
  BUF U7331 ( .I(n28843), .Z(n28784) );
  BUF U7332 ( .I(n28608), .Z(n28549) );
  BUF U7333 ( .I(n28373), .Z(n28314) );
  BUF U7334 ( .I(n28138), .Z(n28079) );
  BUF U7335 ( .I(n27903), .Z(n27844) );
  BUF U7336 ( .I(n27668), .Z(n27609) );
  BUF U7337 ( .I(n29314), .Z(n29253) );
  BUF U7338 ( .I(n29079), .Z(n29018) );
  BUF U7339 ( .I(n28844), .Z(n28783) );
  BUF U7340 ( .I(n28609), .Z(n28548) );
  BUF U7341 ( .I(n28374), .Z(n28313) );
  BUF U7342 ( .I(n28139), .Z(n28078) );
  BUF U7343 ( .I(n27904), .Z(n27843) );
  BUF U7344 ( .I(n27669), .Z(n27608) );
  BUF U7345 ( .I(n29314), .Z(n29252) );
  BUF U7346 ( .I(n29079), .Z(n29017) );
  BUF U7347 ( .I(n28844), .Z(n28782) );
  BUF U7348 ( .I(n28609), .Z(n28547) );
  BUF U7349 ( .I(n28374), .Z(n28312) );
  BUF U7350 ( .I(n28139), .Z(n28077) );
  BUF U7351 ( .I(n27904), .Z(n27842) );
  BUF U7352 ( .I(n27669), .Z(n27607) );
  BUF U7353 ( .I(n29314), .Z(n29251) );
  BUF U7354 ( .I(n29079), .Z(n29016) );
  BUF U7355 ( .I(n28844), .Z(n28781) );
  BUF U7356 ( .I(n28609), .Z(n28546) );
  BUF U7357 ( .I(n28374), .Z(n28311) );
  BUF U7358 ( .I(n28139), .Z(n28076) );
  BUF U7359 ( .I(n27904), .Z(n27841) );
  BUF U7360 ( .I(n27669), .Z(n27606) );
  BUF U7361 ( .I(n29315), .Z(n29250) );
  BUF U7362 ( .I(n29080), .Z(n29015) );
  BUF U7363 ( .I(n28845), .Z(n28780) );
  BUF U7364 ( .I(n28610), .Z(n28545) );
  BUF U7365 ( .I(n28375), .Z(n28310) );
  BUF U7366 ( .I(n28140), .Z(n28075) );
  BUF U7367 ( .I(n27905), .Z(n27840) );
  BUF U7368 ( .I(n27670), .Z(n27605) );
  BUF U7369 ( .I(n29315), .Z(n29249) );
  BUF U7370 ( .I(n29080), .Z(n29014) );
  BUF U7371 ( .I(n28845), .Z(n28779) );
  BUF U7372 ( .I(n28610), .Z(n28544) );
  BUF U7373 ( .I(n28375), .Z(n28309) );
  BUF U7374 ( .I(n28140), .Z(n28074) );
  BUF U7375 ( .I(n27905), .Z(n27839) );
  BUF U7376 ( .I(n27670), .Z(n27604) );
  BUF U7377 ( .I(n29315), .Z(n29248) );
  BUF U7378 ( .I(n29080), .Z(n29013) );
  BUF U7379 ( .I(n28845), .Z(n28778) );
  BUF U7380 ( .I(n28610), .Z(n28543) );
  BUF U7381 ( .I(n28375), .Z(n28308) );
  BUF U7382 ( .I(n28140), .Z(n28073) );
  BUF U7383 ( .I(n27905), .Z(n27838) );
  BUF U7384 ( .I(n27670), .Z(n27603) );
  BUF U7385 ( .I(n29299), .Z(n29298) );
  BUF U7386 ( .I(n29064), .Z(n29063) );
  BUF U7387 ( .I(n28829), .Z(n28828) );
  BUF U7388 ( .I(n28594), .Z(n28593) );
  BUF U7389 ( .I(n28359), .Z(n28358) );
  BUF U7390 ( .I(n28124), .Z(n28123) );
  BUF U7391 ( .I(n27889), .Z(n27888) );
  BUF U7392 ( .I(n27654), .Z(n27653) );
  BUF U7393 ( .I(n29581), .Z(n29572) );
  BUF U7394 ( .I(we), .Z(n29581) );
  BUF U7395 ( .I(we), .Z(n29579) );
  BUF U7396 ( .I(we), .Z(n29580) );
  BUF U7397 ( .I(n27340), .Z(n26867) );
  BUF U7398 ( .I(n26865), .Z(n26392) );
  BUF U7399 ( .I(n27340), .Z(n26868) );
  BUF U7400 ( .I(n26865), .Z(n26393) );
  BUF U7401 ( .I(n26866), .Z(n26881) );
  BUF U7402 ( .I(n26866), .Z(n26880) );
  BUF U7403 ( .I(n26391), .Z(n26405) );
  BUF U7404 ( .I(n27340), .Z(n26869) );
  BUF U7405 ( .I(n26865), .Z(n26394) );
  BUF U7406 ( .I(n26866), .Z(n26879) );
  BUF U7407 ( .I(n26391), .Z(n26404) );
  BUF U7408 ( .I(n26391), .Z(n26406) );
  BUF U7409 ( .I(n26157), .Z(n26158) );
  BUF U7410 ( .I(n26275), .Z(n26276) );
  BUF U7411 ( .I(n26157), .Z(n26159) );
  BUF U7412 ( .I(n26275), .Z(n26277) );
  BUF U7413 ( .I(n26157), .Z(n26160) );
  BUF U7414 ( .I(n26275), .Z(n26278) );
  BUF U7415 ( .I(n26156), .Z(n26161) );
  BUF U7416 ( .I(n26274), .Z(n26279) );
  BUF U7417 ( .I(n26156), .Z(n26162) );
  BUF U7418 ( .I(n26274), .Z(n26280) );
  BUF U7419 ( .I(n26156), .Z(n26163) );
  BUF U7420 ( .I(n26274), .Z(n26281) );
  BUF U7421 ( .I(n26155), .Z(n26164) );
  BUF U7422 ( .I(n26273), .Z(n26282) );
  BUF U7423 ( .I(n26155), .Z(n26165) );
  BUF U7424 ( .I(n26273), .Z(n26283) );
  BUF U7425 ( .I(n26155), .Z(n26166) );
  BUF U7426 ( .I(n26273), .Z(n26284) );
  NOR3 U7427 ( .A1(n29586), .A2(n29585), .A3(n29587), .ZN(n4100) );
  NOR3 U7428 ( .A1(n29583), .A2(n29582), .A3(n29584), .ZN(n4099) );
  NOR3 U7429 ( .A1(n29589), .A2(n29588), .A3(n29590), .ZN(n214) );
  AND2 U7430 ( .A1(n4118), .A2(n4100), .Z(n42) );
  AND2 U7431 ( .A1(n4121), .A2(n4100), .Z(n45) );
  AND2 U7432 ( .A1(n4158), .A2(n4099), .Z(n96) );
  AND2 U7433 ( .A1(n4158), .A2(n4103), .Z(n99) );
  AND2 U7434 ( .A1(n4158), .A2(n4106), .Z(n102) );
  AND2 U7435 ( .A1(n4158), .A2(n4109), .Z(n105) );
  AND2 U7436 ( .A1(n4158), .A2(n4112), .Z(n108) );
  AND2 U7437 ( .A1(n4158), .A2(n4115), .Z(n111) );
  AND2 U7438 ( .A1(n4158), .A2(n4118), .Z(n114) );
  AND2 U7439 ( .A1(n4158), .A2(n4121), .Z(n117) );
  AND2 U7440 ( .A1(n4192), .A2(n4099), .Z(n144) );
  AND2 U7441 ( .A1(n4192), .A2(n4103), .Z(n147) );
  AND2 U7442 ( .A1(n4192), .A2(n4106), .Z(n150) );
  AND2 U7443 ( .A1(n4192), .A2(n4109), .Z(n153) );
  AND2 U7444 ( .A1(n4192), .A2(n4112), .Z(n156) );
  AND2 U7445 ( .A1(n4192), .A2(n4115), .Z(n159) );
  AND2 U7446 ( .A1(n4192), .A2(n4118), .Z(n162) );
  AND2 U7447 ( .A1(n4192), .A2(n4121), .Z(n165) );
  AND2 U7448 ( .A1(n4124), .A2(n4099), .Z(n48) );
  AND2 U7449 ( .A1(n4124), .A2(n4103), .Z(n51) );
  AND2 U7450 ( .A1(n4124), .A2(n4106), .Z(n54) );
  AND2 U7451 ( .A1(n4124), .A2(n4109), .Z(n57) );
  AND2 U7452 ( .A1(n4124), .A2(n4112), .Z(n60) );
  AND2 U7453 ( .A1(n4124), .A2(n4115), .Z(n63) );
  AND2 U7454 ( .A1(n4124), .A2(n4118), .Z(n66) );
  AND2 U7455 ( .A1(n4124), .A2(n4121), .Z(n69) );
  AND2 U7456 ( .A1(n4141), .A2(n4099), .Z(n72) );
  AND2 U7457 ( .A1(n4141), .A2(n4103), .Z(n75) );
  AND2 U7458 ( .A1(n4141), .A2(n4106), .Z(n78) );
  AND2 U7459 ( .A1(n4141), .A2(n4109), .Z(n81) );
  AND2 U7460 ( .A1(n4141), .A2(n4112), .Z(n84) );
  AND2 U7461 ( .A1(n4141), .A2(n4115), .Z(n87) );
  AND2 U7462 ( .A1(n4141), .A2(n4118), .Z(n90) );
  AND2 U7463 ( .A1(n4141), .A2(n4121), .Z(n93) );
  AND2 U7464 ( .A1(n4175), .A2(n4099), .Z(n120) );
  AND2 U7465 ( .A1(n4175), .A2(n4103), .Z(n123) );
  AND2 U7466 ( .A1(n4175), .A2(n4106), .Z(n126) );
  AND2 U7467 ( .A1(n4175), .A2(n4109), .Z(n129) );
  AND2 U7468 ( .A1(n4175), .A2(n4112), .Z(n132) );
  AND2 U7469 ( .A1(n4175), .A2(n4115), .Z(n135) );
  AND2 U7470 ( .A1(n4175), .A2(n4118), .Z(n138) );
  AND2 U7471 ( .A1(n4175), .A2(n4121), .Z(n141) );
  BUF U7472 ( .I(n26104), .Z(n26107) );
  BUF U7473 ( .I(n26104), .Z(n26106) );
  BUF U7474 ( .I(n26104), .Z(n26105) );
  INV U7475 ( .I(n26087), .ZN(n26089) );
  INV U7476 ( .I(n26086), .ZN(n26090) );
  BUF U7477 ( .I(n26134), .Z(n26137) );
  BUF U7478 ( .I(n26134), .Z(n26136) );
  INV U7479 ( .I(n26087), .ZN(n26088) );
  BUF U7480 ( .I(n26134), .Z(n26135) );
  BUF U7481 ( .I(n26096), .Z(n26103) );
  BUF U7482 ( .I(n26126), .Z(n26133) );
  BUF U7483 ( .I(n26096), .Z(n26102) );
  BUF U7484 ( .I(n26126), .Z(n26132) );
  BUF U7485 ( .I(n26096), .Z(n26101) );
  BUF U7486 ( .I(n26126), .Z(n26131) );
  BUF U7487 ( .I(n26097), .Z(n26100) );
  BUF U7488 ( .I(n26127), .Z(n26130) );
  BUF U7489 ( .I(n26097), .Z(n26099) );
  BUF U7490 ( .I(n26127), .Z(n26129) );
  BUF U7491 ( .I(n26097), .Z(n26098) );
  BUF U7492 ( .I(n26127), .Z(n26128) );
  INV U7493 ( .I(n26092), .ZN(n26093) );
  NOR2 U7494 ( .A1(n29591), .A2(n29592), .ZN(n215) );
  BUF U7495 ( .I(n29082), .Z(n29299) );
  BUF U7496 ( .I(n28847), .Z(n29064) );
  BUF U7497 ( .I(n28612), .Z(n28829) );
  BUF U7498 ( .I(n28377), .Z(n28594) );
  BUF U7499 ( .I(n28142), .Z(n28359) );
  BUF U7500 ( .I(n27907), .Z(n28124) );
  BUF U7501 ( .I(n27672), .Z(n27889) );
  BUF U7502 ( .I(n27437), .Z(n27654) );
  BUF U7503 ( .I(n29082), .Z(n29300) );
  BUF U7504 ( .I(n28847), .Z(n29065) );
  BUF U7505 ( .I(n28612), .Z(n28830) );
  BUF U7506 ( .I(n28377), .Z(n28595) );
  BUF U7507 ( .I(n28142), .Z(n28360) );
  BUF U7508 ( .I(n27907), .Z(n28125) );
  BUF U7509 ( .I(n27672), .Z(n27890) );
  BUF U7510 ( .I(n27437), .Z(n27655) );
  BUF U7511 ( .I(n29082), .Z(n29301) );
  BUF U7512 ( .I(n28847), .Z(n29066) );
  BUF U7513 ( .I(n28612), .Z(n28831) );
  BUF U7514 ( .I(n28377), .Z(n28596) );
  BUF U7515 ( .I(n28142), .Z(n28361) );
  BUF U7516 ( .I(n27907), .Z(n28126) );
  BUF U7517 ( .I(n27672), .Z(n27891) );
  BUF U7518 ( .I(n27437), .Z(n27656) );
  BUF U7519 ( .I(n29083), .Z(n29302) );
  BUF U7520 ( .I(n28848), .Z(n29067) );
  BUF U7521 ( .I(n28613), .Z(n28832) );
  BUF U7522 ( .I(n28378), .Z(n28597) );
  BUF U7523 ( .I(n28143), .Z(n28362) );
  BUF U7524 ( .I(n27908), .Z(n28127) );
  BUF U7525 ( .I(n27673), .Z(n27892) );
  BUF U7526 ( .I(n27438), .Z(n27657) );
  BUF U7527 ( .I(n29083), .Z(n29303) );
  BUF U7528 ( .I(n28848), .Z(n29068) );
  BUF U7529 ( .I(n28613), .Z(n28833) );
  BUF U7530 ( .I(n28378), .Z(n28598) );
  BUF U7531 ( .I(n28143), .Z(n28363) );
  BUF U7532 ( .I(n27908), .Z(n28128) );
  BUF U7533 ( .I(n27673), .Z(n27893) );
  BUF U7534 ( .I(n27438), .Z(n27658) );
  BUF U7535 ( .I(n29083), .Z(n29304) );
  BUF U7536 ( .I(n28848), .Z(n29069) );
  BUF U7537 ( .I(n28613), .Z(n28834) );
  BUF U7538 ( .I(n28378), .Z(n28599) );
  BUF U7539 ( .I(n28143), .Z(n28364) );
  BUF U7540 ( .I(n27908), .Z(n28129) );
  BUF U7541 ( .I(n27673), .Z(n27894) );
  BUF U7542 ( .I(n27438), .Z(n27659) );
  BUF U7543 ( .I(n29084), .Z(n29305) );
  BUF U7544 ( .I(n28849), .Z(n29070) );
  BUF U7545 ( .I(n28614), .Z(n28835) );
  BUF U7546 ( .I(n28379), .Z(n28600) );
  BUF U7547 ( .I(n28144), .Z(n28365) );
  BUF U7548 ( .I(n27909), .Z(n28130) );
  BUF U7549 ( .I(n27674), .Z(n27895) );
  BUF U7550 ( .I(n27439), .Z(n27660) );
  BUF U7551 ( .I(n29084), .Z(n29306) );
  BUF U7552 ( .I(n28849), .Z(n29071) );
  BUF U7553 ( .I(n28614), .Z(n28836) );
  BUF U7554 ( .I(n28379), .Z(n28601) );
  BUF U7555 ( .I(n28144), .Z(n28366) );
  BUF U7556 ( .I(n27909), .Z(n28131) );
  BUF U7557 ( .I(n27674), .Z(n27896) );
  BUF U7558 ( .I(n27439), .Z(n27661) );
  BUF U7559 ( .I(n29084), .Z(n29307) );
  BUF U7560 ( .I(n28849), .Z(n29072) );
  BUF U7561 ( .I(n28614), .Z(n28837) );
  BUF U7562 ( .I(n28379), .Z(n28602) );
  BUF U7563 ( .I(n28144), .Z(n28367) );
  BUF U7564 ( .I(n27909), .Z(n28132) );
  BUF U7565 ( .I(n27674), .Z(n27897) );
  BUF U7566 ( .I(n27439), .Z(n27662) );
  BUF U7567 ( .I(n29085), .Z(n29308) );
  BUF U7568 ( .I(n28850), .Z(n29073) );
  BUF U7569 ( .I(n28615), .Z(n28838) );
  BUF U7570 ( .I(n28380), .Z(n28603) );
  BUF U7571 ( .I(n28145), .Z(n28368) );
  BUF U7572 ( .I(n27910), .Z(n28133) );
  BUF U7573 ( .I(n27675), .Z(n27898) );
  BUF U7574 ( .I(n27440), .Z(n27663) );
  BUF U7575 ( .I(n29085), .Z(n29309) );
  BUF U7576 ( .I(n28850), .Z(n29074) );
  BUF U7577 ( .I(n28615), .Z(n28839) );
  BUF U7578 ( .I(n28380), .Z(n28604) );
  BUF U7579 ( .I(n28145), .Z(n28369) );
  BUF U7580 ( .I(n27910), .Z(n28134) );
  BUF U7581 ( .I(n27675), .Z(n27899) );
  BUF U7582 ( .I(n27440), .Z(n27664) );
  BUF U7583 ( .I(n29085), .Z(n29310) );
  BUF U7584 ( .I(n28850), .Z(n29075) );
  BUF U7585 ( .I(n28615), .Z(n28840) );
  BUF U7586 ( .I(n28380), .Z(n28605) );
  BUF U7587 ( .I(n28145), .Z(n28370) );
  BUF U7588 ( .I(n27910), .Z(n28135) );
  BUF U7589 ( .I(n27675), .Z(n27900) );
  BUF U7590 ( .I(n27440), .Z(n27665) );
  BUF U7591 ( .I(n29086), .Z(n29311) );
  BUF U7592 ( .I(n28851), .Z(n29076) );
  BUF U7593 ( .I(n28616), .Z(n28841) );
  BUF U7594 ( .I(n28381), .Z(n28606) );
  BUF U7595 ( .I(n28146), .Z(n28371) );
  BUF U7596 ( .I(n27911), .Z(n28136) );
  BUF U7597 ( .I(n27676), .Z(n27901) );
  BUF U7598 ( .I(n27441), .Z(n27666) );
  BUF U7599 ( .I(n29086), .Z(n29312) );
  BUF U7600 ( .I(n28851), .Z(n29077) );
  BUF U7601 ( .I(n28616), .Z(n28842) );
  BUF U7602 ( .I(n28381), .Z(n28607) );
  BUF U7603 ( .I(n28146), .Z(n28372) );
  BUF U7604 ( .I(n27911), .Z(n28137) );
  BUF U7605 ( .I(n27676), .Z(n27902) );
  BUF U7606 ( .I(n27441), .Z(n27667) );
  BUF U7607 ( .I(n29086), .Z(n29313) );
  BUF U7608 ( .I(n28851), .Z(n29078) );
  BUF U7609 ( .I(n28616), .Z(n28843) );
  BUF U7610 ( .I(n28381), .Z(n28608) );
  BUF U7611 ( .I(n28146), .Z(n28373) );
  BUF U7612 ( .I(n27911), .Z(n28138) );
  BUF U7613 ( .I(n27676), .Z(n27903) );
  BUF U7614 ( .I(n27441), .Z(n27668) );
  BUF U7615 ( .I(n29087), .Z(n29314) );
  BUF U7616 ( .I(n28852), .Z(n29079) );
  BUF U7617 ( .I(n28617), .Z(n28844) );
  BUF U7618 ( .I(n28382), .Z(n28609) );
  BUF U7619 ( .I(n28147), .Z(n28374) );
  BUF U7620 ( .I(n27912), .Z(n28139) );
  BUF U7621 ( .I(n27677), .Z(n27904) );
  BUF U7622 ( .I(n27442), .Z(n27669) );
  BUF U7623 ( .I(n29087), .Z(n29315) );
  BUF U7624 ( .I(n28852), .Z(n29080) );
  BUF U7625 ( .I(n28617), .Z(n28845) );
  BUF U7626 ( .I(n28382), .Z(n28610) );
  BUF U7627 ( .I(n28147), .Z(n28375) );
  BUF U7628 ( .I(n27912), .Z(n28140) );
  BUF U7629 ( .I(n27677), .Z(n27905) );
  BUF U7630 ( .I(n27442), .Z(n27670) );
  BUF U7631 ( .I(n29087), .Z(n29316) );
  BUF U7632 ( .I(n28852), .Z(n29081) );
  BUF U7633 ( .I(n28617), .Z(n28846) );
  BUF U7634 ( .I(n28382), .Z(n28611) );
  BUF U7635 ( .I(n28147), .Z(n28376) );
  BUF U7636 ( .I(n27912), .Z(n28141) );
  BUF U7637 ( .I(n27677), .Z(n27906) );
  BUF U7638 ( .I(n27442), .Z(n27671) );
  MUX41 U7639 ( .I0(n20694), .I1(n20695), .I2(n20696), .I3(n20697), .S0(
        n26088), .S1(n26094), .ZN(n20693) );
  MUX41 U7640 ( .I0(n20779), .I1(n20780), .I2(n20781), .I3(n20782), .S0(
        n26088), .S1(n26094), .ZN(n20778) );
  MUX41 U7641 ( .I0(n20648), .I1(n20638), .I2(n20643), .I3(n20633), .S0(
        n26105), .S1(n26135), .ZN(n20695) );
  MUX41 U7642 ( .I0(n21378), .I1(n21379), .I2(n21380), .I3(n21381), .S0(
        n26088), .S1(n26094), .ZN(n21377) );
  MUX41 U7643 ( .I0(n21463), .I1(n21464), .I2(n21465), .I3(n21466), .S0(
        n26088), .S1(n26094), .ZN(n21462) );
  MUX41 U7644 ( .I0(n21332), .I1(n21322), .I2(n21327), .I3(n21317), .S0(
        n26107), .S1(n26137), .ZN(n21379) );
  MUX41 U7645 ( .I0(n22062), .I1(n22063), .I2(n22064), .I3(n22065), .S0(
        n26089), .S1(n26094), .ZN(n22061) );
  MUX41 U7646 ( .I0(n22147), .I1(n22148), .I2(n22149), .I3(n22150), .S0(
        n26089), .S1(n26093), .ZN(n22146) );
  MUX41 U7647 ( .I0(n22016), .I1(n22006), .I2(n22011), .I3(n22001), .S0(
        n26110), .S1(n26140), .ZN(n22063) );
  MUX41 U7648 ( .I0(n22746), .I1(n22747), .I2(n22748), .I3(n22749), .S0(
        n26089), .S1(n26094), .ZN(n22745) );
  MUX41 U7649 ( .I0(n22831), .I1(n22832), .I2(n22833), .I3(n22834), .S0(
        n26090), .S1(n26093), .ZN(n22830) );
  MUX41 U7650 ( .I0(n22700), .I1(n22690), .I2(n22695), .I3(n22685), .S0(
        n26112), .S1(n26142), .ZN(n22747) );
  MUX41 U7651 ( .I0(n23430), .I1(n23431), .I2(n23432), .I3(n23433), .S0(
        n26090), .S1(n26093), .ZN(n23429) );
  MUX41 U7652 ( .I0(n23515), .I1(n23516), .I2(n23517), .I3(n23518), .S0(
        n26090), .S1(n26093), .ZN(n23514) );
  MUX41 U7653 ( .I0(n23384), .I1(n23374), .I2(n23379), .I3(n23369), .S0(
        n26115), .S1(n26145), .ZN(n23431) );
  MUX41 U7654 ( .I0(n24114), .I1(n24115), .I2(n24116), .I3(n24117), .S0(
        n26090), .S1(n26093), .ZN(n24113) );
  MUX41 U7655 ( .I0(n24199), .I1(n24200), .I2(n24201), .I3(n24202), .S0(
        n26089), .S1(n26093), .ZN(n24198) );
  MUX41 U7656 ( .I0(n24068), .I1(n24058), .I2(n24063), .I3(n24053), .S0(
        n26117), .S1(n26147), .ZN(n24115) );
  MUX41 U7657 ( .I0(n24798), .I1(n24799), .I2(n24800), .I3(n24801), .S0(
        n26088), .S1(n26093), .ZN(n24797) );
  MUX41 U7658 ( .I0(n24883), .I1(n24884), .I2(n24885), .I3(n24886), .S0(
        n26088), .S1(n26093), .ZN(n24882) );
  MUX41 U7659 ( .I0(n24752), .I1(n24742), .I2(n24747), .I3(n24737), .S0(
        n26120), .S1(n26150), .ZN(n24799) );
  MUX41 U7660 ( .I0(n25482), .I1(n25483), .I2(n25484), .I3(n25485), .S0(
        n26090), .S1(n26094), .ZN(n25481) );
  MUX41 U7661 ( .I0(n25567), .I1(n25568), .I2(n25569), .I3(n25570), .S0(
        n26089), .S1(n26094), .ZN(n25566) );
  MUX41 U7662 ( .I0(n25436), .I1(n25426), .I2(n25431), .I3(n25421), .S0(
        n26122), .S1(n26152), .ZN(n25483) );
  MUX41 U7663 ( .I0(n20713), .I1(n20703), .I2(n20708), .I3(n20698), .S0(
        n26105), .S1(n26135), .ZN(n20782) );
  MUX41 U7664 ( .I0(n20699), .I1(n20700), .I2(n20701), .I3(n20702), .S0(
        n26195), .S1(n26313), .ZN(n20698) );
  MUX41 U7665 ( .I0(n20704), .I1(n20705), .I2(n20706), .I3(n20707), .S0(
        n26195), .S1(n26313), .ZN(n20703) );
  MUX41 U7666 ( .I0(n20714), .I1(n20715), .I2(n20716), .I3(n20717), .S0(
        n26195), .S1(n26313), .ZN(n20713) );
  MUX41 U7667 ( .I0(n20628), .I1(n3324), .I2(n3969), .I3(n2678), .S0(
        n26105), .S1(n26135), .ZN(n20697) );
  MUX41 U7668 ( .I0(n2807), .I1(n2936), .I2(n3065), .I3(n3194), .S0(
        n26194), .S1(n26312), .ZN(n2678) );
  MUX41 U7669 ( .I0(n3453), .I1(n3582), .I2(n3711), .I3(n3840), .S0(
        n26194), .S1(n26312), .ZN(n3324) );
  MUX41 U7670 ( .I0(n20629), .I1(n20630), .I2(n20631), .I3(n20632), .S0(
        n26194), .S1(n26312), .ZN(n20628) );
  MUX41 U7671 ( .I0(n21397), .I1(n21387), .I2(n21392), .I3(n21382), .S0(
        n26108), .S1(n26138), .ZN(n21466) );
  MUX41 U7672 ( .I0(n21383), .I1(n21384), .I2(n21385), .I3(n21386), .S0(
        n26205), .S1(n26323), .ZN(n21382) );
  MUX41 U7673 ( .I0(n21388), .I1(n21389), .I2(n21390), .I3(n21391), .S0(
        n26205), .S1(n26323), .ZN(n21387) );
  MUX41 U7674 ( .I0(n21398), .I1(n21399), .I2(n21400), .I3(n21401), .S0(
        n26205), .S1(n26323), .ZN(n21397) );
  MUX41 U7675 ( .I0(n21312), .I1(n21302), .I2(n21307), .I3(n21297), .S0(
        n26107), .S1(n26137), .ZN(n21381) );
  MUX41 U7676 ( .I0(n21298), .I1(n21299), .I2(n21300), .I3(n21301), .S0(
        n26204), .S1(n26322), .ZN(n21297) );
  MUX41 U7677 ( .I0(n21303), .I1(n21304), .I2(n21305), .I3(n21306), .S0(
        n26204), .S1(n26322), .ZN(n21302) );
  MUX41 U7678 ( .I0(n21313), .I1(n21314), .I2(n21315), .I3(n21316), .S0(
        n26204), .S1(n26322), .ZN(n21312) );
  MUX41 U7679 ( .I0(n22081), .I1(n22071), .I2(n22076), .I3(n22066), .S0(
        n26110), .S1(n26140), .ZN(n22150) );
  MUX41 U7680 ( .I0(n22067), .I1(n22068), .I2(n22069), .I3(n22070), .S0(
        n26215), .S1(n26333), .ZN(n22066) );
  MUX41 U7681 ( .I0(n22072), .I1(n22073), .I2(n22074), .I3(n22075), .S0(
        n26215), .S1(n26333), .ZN(n22071) );
  MUX41 U7682 ( .I0(n22082), .I1(n22083), .I2(n22084), .I3(n22085), .S0(
        n26215), .S1(n26333), .ZN(n22081) );
  MUX41 U7683 ( .I0(n21996), .I1(n21986), .I2(n21991), .I3(n21981), .S0(
        n26110), .S1(n26140), .ZN(n22065) );
  MUX41 U7684 ( .I0(n21982), .I1(n21983), .I2(n21984), .I3(n21985), .S0(
        n26213), .S1(n26331), .ZN(n21981) );
  MUX41 U7685 ( .I0(n21987), .I1(n21988), .I2(n21989), .I3(n21990), .S0(
        n26214), .S1(n26332), .ZN(n21986) );
  MUX41 U7686 ( .I0(n21997), .I1(n21998), .I2(n21999), .I3(n22000), .S0(
        n26214), .S1(n26332), .ZN(n21996) );
  MUX41 U7687 ( .I0(n22765), .I1(n22755), .I2(n22760), .I3(n22750), .S0(
        n26113), .S1(n26143), .ZN(n22834) );
  MUX41 U7688 ( .I0(n22751), .I1(n22752), .I2(n22753), .I3(n22754), .S0(
        n26225), .S1(n26343), .ZN(n22750) );
  MUX41 U7689 ( .I0(n22756), .I1(n22757), .I2(n22758), .I3(n22759), .S0(
        n26225), .S1(n26343), .ZN(n22755) );
  MUX41 U7690 ( .I0(n22766), .I1(n22767), .I2(n22768), .I3(n22769), .S0(
        n26225), .S1(n26343), .ZN(n22765) );
  MUX41 U7691 ( .I0(n22680), .I1(n22670), .I2(n22675), .I3(n22665), .S0(
        n26112), .S1(n26142), .ZN(n22749) );
  MUX41 U7692 ( .I0(n22666), .I1(n22667), .I2(n22668), .I3(n22669), .S0(
        n26223), .S1(n26341), .ZN(n22665) );
  MUX41 U7693 ( .I0(n22671), .I1(n22672), .I2(n22673), .I3(n22674), .S0(
        n26223), .S1(n26341), .ZN(n22670) );
  MUX41 U7694 ( .I0(n22681), .I1(n22682), .I2(n22683), .I3(n22684), .S0(
        n26224), .S1(n26342), .ZN(n22680) );
  MUX41 U7695 ( .I0(n23449), .I1(n23439), .I2(n23444), .I3(n23434), .S0(
        n26115), .S1(n26145), .ZN(n23518) );
  MUX41 U7696 ( .I0(n23435), .I1(n23436), .I2(n23437), .I3(n23438), .S0(
        n26234), .S1(n26352), .ZN(n23434) );
  MUX41 U7697 ( .I0(n23440), .I1(n23441), .I2(n23442), .I3(n23443), .S0(
        n26234), .S1(n26352), .ZN(n23439) );
  MUX41 U7698 ( .I0(n23450), .I1(n23451), .I2(n23452), .I3(n23453), .S0(
        n26235), .S1(n26353), .ZN(n23449) );
  MUX41 U7699 ( .I0(n23364), .I1(n23354), .I2(n23359), .I3(n23349), .S0(
        n26115), .S1(n26145), .ZN(n23433) );
  MUX41 U7700 ( .I0(n23350), .I1(n23351), .I2(n23352), .I3(n23353), .S0(
        n26233), .S1(n26351), .ZN(n23349) );
  MUX41 U7701 ( .I0(n23355), .I1(n23356), .I2(n23357), .I3(n23358), .S0(
        n26233), .S1(n26351), .ZN(n23354) );
  MUX41 U7702 ( .I0(n23365), .I1(n23366), .I2(n23367), .I3(n23368), .S0(
        n26233), .S1(n26351), .ZN(n23364) );
  MUX41 U7703 ( .I0(n24133), .I1(n24123), .I2(n24128), .I3(n24118), .S0(
        n26117), .S1(n26147), .ZN(n24202) );
  MUX41 U7704 ( .I0(n24119), .I1(n24120), .I2(n24121), .I3(n24122), .S0(
        n26244), .S1(n26362), .ZN(n24118) );
  MUX41 U7705 ( .I0(n24124), .I1(n24125), .I2(n24126), .I3(n24127), .S0(
        n26244), .S1(n26362), .ZN(n24123) );
  MUX41 U7706 ( .I0(n24134), .I1(n24135), .I2(n24136), .I3(n24137), .S0(
        n26244), .S1(n26362), .ZN(n24133) );
  MUX41 U7707 ( .I0(n24048), .I1(n24038), .I2(n24043), .I3(n24033), .S0(
        n26117), .S1(n26147), .ZN(n24117) );
  MUX41 U7708 ( .I0(n24034), .I1(n24035), .I2(n24036), .I3(n24037), .S0(
        n26243), .S1(n26361), .ZN(n24033) );
  MUX41 U7709 ( .I0(n24039), .I1(n24040), .I2(n24041), .I3(n24042), .S0(
        n26243), .S1(n26361), .ZN(n24038) );
  MUX41 U7710 ( .I0(n24049), .I1(n24050), .I2(n24051), .I3(n24052), .S0(
        n26243), .S1(n26361), .ZN(n24048) );
  MUX41 U7711 ( .I0(n24817), .I1(n24807), .I2(n24812), .I3(n24802), .S0(
        n26120), .S1(n26150), .ZN(n24886) );
  MUX41 U7712 ( .I0(n24803), .I1(n24804), .I2(n24805), .I3(n24806), .S0(
        n26254), .S1(n26372), .ZN(n24802) );
  MUX41 U7713 ( .I0(n24808), .I1(n24809), .I2(n24810), .I3(n24811), .S0(
        n26254), .S1(n26372), .ZN(n24807) );
  MUX41 U7714 ( .I0(n24818), .I1(n24819), .I2(n24820), .I3(n24821), .S0(
        n26254), .S1(n26372), .ZN(n24817) );
  MUX41 U7715 ( .I0(n24732), .I1(n24722), .I2(n24727), .I3(n24717), .S0(
        n26120), .S1(n26150), .ZN(n24801) );
  MUX41 U7716 ( .I0(n24718), .I1(n24719), .I2(n24720), .I3(n24721), .S0(
        n26253), .S1(n26371), .ZN(n24717) );
  MUX41 U7717 ( .I0(n24723), .I1(n24724), .I2(n24725), .I3(n24726), .S0(
        n26253), .S1(n26371), .ZN(n24722) );
  MUX41 U7718 ( .I0(n24733), .I1(n24734), .I2(n24735), .I3(n24736), .S0(
        n26253), .S1(n26371), .ZN(n24732) );
  MUX41 U7719 ( .I0(n25501), .I1(n25491), .I2(n25496), .I3(n25486), .S0(
        n26122), .S1(n26152), .ZN(n25570) );
  MUX41 U7720 ( .I0(n25487), .I1(n25488), .I2(n25489), .I3(n25490), .S0(
        n26264), .S1(n26382), .ZN(n25486) );
  MUX41 U7721 ( .I0(n25492), .I1(n25493), .I2(n25494), .I3(n25495), .S0(
        n26264), .S1(n26382), .ZN(n25491) );
  MUX41 U7722 ( .I0(n25502), .I1(n25503), .I2(n25504), .I3(n25505), .S0(
        n26264), .S1(n26382), .ZN(n25501) );
  MUX41 U7723 ( .I0(n25416), .I1(n25406), .I2(n25411), .I3(n25401), .S0(
        n26122), .S1(n26152), .ZN(n25485) );
  MUX41 U7724 ( .I0(n25402), .I1(n25403), .I2(n25404), .I3(n25405), .S0(
        n26263), .S1(n26381), .ZN(n25401) );
  MUX41 U7725 ( .I0(n25407), .I1(n25408), .I2(n25409), .I3(n25410), .S0(
        n26263), .S1(n26381), .ZN(n25406) );
  MUX41 U7726 ( .I0(n25417), .I1(n25418), .I2(n25419), .I3(n25420), .S0(
        n26263), .S1(n26381), .ZN(n25416) );
  MUX41 U7727 ( .I0(n20733), .I1(n20723), .I2(n20728), .I3(n20718), .S0(
        n26105), .S1(n26135), .ZN(n20780) );
  MUX41 U7728 ( .I0(n20719), .I1(n20720), .I2(n20721), .I3(n20722), .S0(
        n26195), .S1(n26313), .ZN(n20718) );
  MUX41 U7729 ( .I0(n20724), .I1(n20725), .I2(n20726), .I3(n20727), .S0(
        n26195), .S1(n26313), .ZN(n20723) );
  MUX41 U7730 ( .I0(n20734), .I1(n20735), .I2(n20736), .I3(n20737), .S0(
        n26196), .S1(n26314), .ZN(n20733) );
  MUX41 U7731 ( .I0(n21417), .I1(n21407), .I2(n21412), .I3(n21402), .S0(
        n26108), .S1(n26138), .ZN(n21464) );
  MUX41 U7732 ( .I0(n21403), .I1(n21404), .I2(n21405), .I3(n21406), .S0(
        n26205), .S1(n26323), .ZN(n21402) );
  MUX41 U7733 ( .I0(n21408), .I1(n21409), .I2(n21410), .I3(n21411), .S0(
        n26205), .S1(n26323), .ZN(n21407) );
  MUX41 U7734 ( .I0(n21418), .I1(n21419), .I2(n21420), .I3(n21421), .S0(
        n26205), .S1(n26323), .ZN(n21417) );
  MUX41 U7735 ( .I0(n22101), .I1(n22091), .I2(n22096), .I3(n22086), .S0(
        n26110), .S1(n26140), .ZN(n22148) );
  MUX41 U7736 ( .I0(n22087), .I1(n22088), .I2(n22089), .I3(n22090), .S0(
        n26215), .S1(n26333), .ZN(n22086) );
  MUX41 U7737 ( .I0(n22092), .I1(n22093), .I2(n22094), .I3(n22095), .S0(
        n26215), .S1(n26333), .ZN(n22091) );
  MUX41 U7738 ( .I0(n22102), .I1(n22103), .I2(n22104), .I3(n22105), .S0(
        n26215), .S1(n26333), .ZN(n22101) );
  MUX41 U7739 ( .I0(n22785), .I1(n22775), .I2(n22780), .I3(n22770), .S0(
        n26113), .S1(n26143), .ZN(n22832) );
  MUX41 U7740 ( .I0(n22771), .I1(n22772), .I2(n22773), .I3(n22774), .S0(
        n26225), .S1(n26343), .ZN(n22770) );
  MUX41 U7741 ( .I0(n22776), .I1(n22777), .I2(n22778), .I3(n22779), .S0(
        n26225), .S1(n26343), .ZN(n22775) );
  MUX41 U7742 ( .I0(n22786), .I1(n22787), .I2(n22788), .I3(n22789), .S0(
        n26225), .S1(n26343), .ZN(n22785) );
  MUX41 U7743 ( .I0(n23469), .I1(n23459), .I2(n23464), .I3(n23454), .S0(
        n26115), .S1(n26145), .ZN(n23516) );
  MUX41 U7744 ( .I0(n23455), .I1(n23456), .I2(n23457), .I3(n23458), .S0(
        n26235), .S1(n26353), .ZN(n23454) );
  MUX41 U7745 ( .I0(n23460), .I1(n23461), .I2(n23462), .I3(n23463), .S0(
        n26235), .S1(n26353), .ZN(n23459) );
  MUX41 U7746 ( .I0(n23470), .I1(n23471), .I2(n23472), .I3(n23473), .S0(
        n26235), .S1(n26353), .ZN(n23469) );
  MUX41 U7747 ( .I0(n24153), .I1(n24143), .I2(n24148), .I3(n24138), .S0(
        n26118), .S1(n26148), .ZN(n24200) );
  MUX41 U7748 ( .I0(n24139), .I1(n24140), .I2(n24141), .I3(n24142), .S0(
        n26245), .S1(n26363), .ZN(n24138) );
  MUX41 U7749 ( .I0(n24144), .I1(n24145), .I2(n24146), .I3(n24147), .S0(
        n26245), .S1(n26363), .ZN(n24143) );
  MUX41 U7750 ( .I0(n24154), .I1(n24155), .I2(n24156), .I3(n24157), .S0(
        n26245), .S1(n26363), .ZN(n24153) );
  MUX41 U7751 ( .I0(n24837), .I1(n24827), .I2(n24832), .I3(n24822), .S0(
        n26120), .S1(n26150), .ZN(n24884) );
  MUX41 U7752 ( .I0(n24823), .I1(n24824), .I2(n24825), .I3(n24826), .S0(
        n26254), .S1(n26372), .ZN(n24822) );
  MUX41 U7753 ( .I0(n24828), .I1(n24829), .I2(n24830), .I3(n24831), .S0(
        n26254), .S1(n26372), .ZN(n24827) );
  MUX41 U7754 ( .I0(n24838), .I1(n24839), .I2(n24840), .I3(n24841), .S0(
        n26255), .S1(n26373), .ZN(n24837) );
  MUX41 U7755 ( .I0(n25521), .I1(n25511), .I2(n25516), .I3(n25506), .S0(
        n26122), .S1(n26152), .ZN(n25568) );
  MUX41 U7756 ( .I0(n25507), .I1(n25508), .I2(n25509), .I3(n25510), .S0(
        n26264), .S1(n26382), .ZN(n25506) );
  MUX41 U7757 ( .I0(n25512), .I1(n25513), .I2(n25514), .I3(n25515), .S0(
        n26264), .S1(n26382), .ZN(n25511) );
  MUX41 U7758 ( .I0(n25522), .I1(n25523), .I2(n25524), .I3(n25525), .S0(
        n26264), .S1(n26382), .ZN(n25521) );
  MUX41 U7759 ( .I0(n22233), .I1(n22234), .I2(n22235), .I3(n22236), .S0(
        n26089), .S1(n26093), .ZN(n22232) );
  MUX41 U7760 ( .I0(n22187), .I1(n22177), .I2(n22182), .I3(n22172), .S0(
        n26110), .S1(n26140), .ZN(n22234) );
  MUX41 U7761 ( .I0(n22167), .I1(n22157), .I2(n22162), .I3(n22152), .S0(
        n26110), .S1(n26140), .ZN(n22236) );
  MUX41 U7762 ( .I0(n22227), .I1(n22217), .I2(n22222), .I3(n22212), .S0(
        n26111), .S1(n26141), .ZN(n22233) );
  MUX41 U7763 ( .I0(n22917), .I1(n22918), .I2(n22919), .I3(n22920), .S0(
        n26090), .S1(n26093), .ZN(n22916) );
  MUX41 U7764 ( .I0(n22871), .I1(n22861), .I2(n22866), .I3(n22856), .S0(
        n26113), .S1(n26143), .ZN(n22918) );
  MUX41 U7765 ( .I0(n22851), .I1(n22841), .I2(n22846), .I3(n22836), .S0(
        n26113), .S1(n26143), .ZN(n22920) );
  MUX41 U7766 ( .I0(n22911), .I1(n22901), .I2(n22906), .I3(n22896), .S0(
        n26113), .S1(n26143), .ZN(n22917) );
  MUX41 U7767 ( .I0(n23601), .I1(n23602), .I2(n23603), .I3(n23604), .S0(
        n26090), .S1(n26093), .ZN(n23600) );
  MUX41 U7768 ( .I0(n23555), .I1(n23545), .I2(n23550), .I3(n23540), .S0(
        n26115), .S1(n26145), .ZN(n23602) );
  MUX41 U7769 ( .I0(n23535), .I1(n23525), .I2(n23530), .I3(n23520), .S0(
        n26115), .S1(n26145), .ZN(n23604) );
  MUX41 U7770 ( .I0(n23595), .I1(n23585), .I2(n23590), .I3(n23580), .S0(
        n26116), .S1(n26146), .ZN(n23601) );
  MUX41 U7771 ( .I0(n24285), .I1(n24286), .I2(n24287), .I3(n24288), .S0(
        n26088), .S1(n26093), .ZN(n24284) );
  MUX41 U7772 ( .I0(n24239), .I1(n24229), .I2(n24234), .I3(n24224), .S0(
        n26118), .S1(n26148), .ZN(n24286) );
  MUX41 U7773 ( .I0(n24219), .I1(n24209), .I2(n24214), .I3(n24204), .S0(
        n26118), .S1(n26148), .ZN(n24288) );
  MUX41 U7774 ( .I0(n24279), .I1(n24269), .I2(n24274), .I3(n24264), .S0(
        n26118), .S1(n26148), .ZN(n24285) );
  MUX41 U7775 ( .I0(n24969), .I1(n24970), .I2(n24971), .I3(n24972), .S0(
        n26090), .S1(n26094), .ZN(n24968) );
  MUX41 U7776 ( .I0(n24923), .I1(n24913), .I2(n24918), .I3(n24908), .S0(
        n26120), .S1(n26150), .ZN(n24970) );
  MUX41 U7777 ( .I0(n24903), .I1(n24893), .I2(n24898), .I3(n24888), .S0(
        n26120), .S1(n26150), .ZN(n24972) );
  MUX41 U7778 ( .I0(n24963), .I1(n24953), .I2(n24958), .I3(n24948), .S0(
        n26120), .S1(n26150), .ZN(n24969) );
  MUX41 U7779 ( .I0(n25653), .I1(n25654), .I2(n25655), .I3(n25656), .S0(
        n26090), .S1(n26094), .ZN(n25652) );
  MUX41 U7780 ( .I0(n25607), .I1(n25597), .I2(n25602), .I3(n25592), .S0(
        n26123), .S1(n26153), .ZN(n25654) );
  MUX41 U7781 ( .I0(n25587), .I1(n25577), .I2(n25582), .I3(n25572), .S0(
        n26123), .S1(n26153), .ZN(n25656) );
  MUX41 U7782 ( .I0(n25647), .I1(n25637), .I2(n25642), .I3(n25632), .S0(
        n26123), .S1(n26153), .ZN(n25653) );
  MUX41 U7783 ( .I0(n20865), .I1(n20866), .I2(n20867), .I3(n20868), .S0(
        n26088), .S1(n26093), .ZN(n20864) );
  MUX41 U7784 ( .I0(n20819), .I1(n20809), .I2(n20814), .I3(n20804), .S0(
        n26106), .S1(n26136), .ZN(n20866) );
  MUX41 U7785 ( .I0(n20799), .I1(n20789), .I2(n20794), .I3(n20784), .S0(
        n26105), .S1(n26135), .ZN(n20868) );
  MUX41 U7786 ( .I0(n20859), .I1(n20849), .I2(n20854), .I3(n20844), .S0(
        n26106), .S1(n26136), .ZN(n20865) );
  MUX41 U7787 ( .I0(n21549), .I1(n21550), .I2(n21551), .I3(n21552), .S0(
        n26088), .S1(n26094), .ZN(n21548) );
  MUX41 U7788 ( .I0(n21503), .I1(n21493), .I2(n21498), .I3(n21488), .S0(
        n26108), .S1(n26138), .ZN(n21550) );
  MUX41 U7789 ( .I0(n21483), .I1(n21473), .I2(n21478), .I3(n21468), .S0(
        n26108), .S1(n26138), .ZN(n21552) );
  MUX41 U7790 ( .I0(n21543), .I1(n21533), .I2(n21538), .I3(n21528), .S0(
        n26108), .S1(n26138), .ZN(n21549) );
  MUX41 U7791 ( .I0(n21891), .I1(n21892), .I2(n21893), .I3(n21894), .S0(
        n26089), .S1(n26093), .ZN(n21890) );
  MUX41 U7792 ( .I0(n21825), .I1(n21815), .I2(n21820), .I3(n21810), .S0(
        n26109), .S1(n26139), .ZN(n21894) );
  MUX41 U7793 ( .I0(n21845), .I1(n21835), .I2(n21840), .I3(n21830), .S0(
        n26109), .S1(n26139), .ZN(n21892) );
  MUX41 U7794 ( .I0(n21885), .I1(n21875), .I2(n21880), .I3(n21870), .S0(
        n26109), .S1(n26139), .ZN(n21891) );
  MUX41 U7795 ( .I0(n21720), .I1(n21721), .I2(n21722), .I3(n21723), .S0(
        n26089), .S1(n26094), .ZN(n21719) );
  MUX41 U7796 ( .I0(n21674), .I1(n21664), .I2(n21669), .I3(n21659), .S0(
        n26109), .S1(n26139), .ZN(n21721) );
  MUX41 U7797 ( .I0(n21654), .I1(n21644), .I2(n21649), .I3(n21639), .S0(
        n26109), .S1(n26139), .ZN(n21723) );
  MUX41 U7798 ( .I0(n21714), .I1(n21704), .I2(n21709), .I3(n21699), .S0(
        n26109), .S1(n26139), .ZN(n21720) );
  MUX41 U7799 ( .I0(n22575), .I1(n22576), .I2(n22577), .I3(n22578), .S0(
        n26089), .S1(n26093), .ZN(n22574) );
  MUX41 U7800 ( .I0(n22509), .I1(n22499), .I2(n22504), .I3(n22494), .S0(
        n26112), .S1(n26142), .ZN(n22578) );
  MUX41 U7801 ( .I0(n22529), .I1(n22519), .I2(n22524), .I3(n22514), .S0(
        n26112), .S1(n26142), .ZN(n22576) );
  MUX41 U7802 ( .I0(n22569), .I1(n22559), .I2(n22564), .I3(n22554), .S0(
        n26112), .S1(n26142), .ZN(n22575) );
  MUX41 U7803 ( .I0(n22404), .I1(n22405), .I2(n22406), .I3(n22407), .S0(
        n26089), .S1(n26094), .ZN(n22403) );
  MUX41 U7804 ( .I0(n22358), .I1(n22348), .I2(n22353), .I3(n22343), .S0(
        n26111), .S1(n26141), .ZN(n22405) );
  MUX41 U7805 ( .I0(n22338), .I1(n22328), .I2(n22333), .I3(n22323), .S0(
        n26111), .S1(n26141), .ZN(n22407) );
  MUX41 U7806 ( .I0(n22398), .I1(n22388), .I2(n22393), .I3(n22383), .S0(
        n26111), .S1(n26141), .ZN(n22404) );
  MUX41 U7807 ( .I0(n23259), .I1(n23260), .I2(n23261), .I3(n23262), .S0(
        n26090), .S1(n26093), .ZN(n23258) );
  MUX41 U7808 ( .I0(n23193), .I1(n23183), .I2(n23188), .I3(n23178), .S0(
        n26114), .S1(n26144), .ZN(n23262) );
  MUX41 U7809 ( .I0(n23213), .I1(n23203), .I2(n23208), .I3(n23198), .S0(
        n26114), .S1(n26144), .ZN(n23260) );
  MUX41 U7810 ( .I0(n23253), .I1(n23243), .I2(n23248), .I3(n23238), .S0(
        n26114), .S1(n26144), .ZN(n23259) );
  MUX41 U7811 ( .I0(n23088), .I1(n23089), .I2(n23090), .I3(n23091), .S0(
        n26090), .S1(n26093), .ZN(n23087) );
  MUX41 U7812 ( .I0(n23042), .I1(n23032), .I2(n23037), .I3(n23027), .S0(
        n26114), .S1(n26144), .ZN(n23089) );
  MUX41 U7813 ( .I0(n23022), .I1(n23012), .I2(n23017), .I3(n23007), .S0(
        n26113), .S1(n26143), .ZN(n23091) );
  MUX41 U7814 ( .I0(n23082), .I1(n23072), .I2(n23077), .I3(n23067), .S0(
        n26114), .S1(n26144), .ZN(n23088) );
  MUX41 U7815 ( .I0(n23943), .I1(n23944), .I2(n23945), .I3(n23946), .S0(
        n26090), .S1(raddr[6]), .ZN(n23942) );
  MUX41 U7816 ( .I0(n23877), .I1(n23867), .I2(n23872), .I3(n23862), .S0(
        n26117), .S1(n26147), .ZN(n23946) );
  MUX41 U7817 ( .I0(n23897), .I1(n23887), .I2(n23892), .I3(n23882), .S0(
        n26117), .S1(n26147), .ZN(n23944) );
  MUX41 U7818 ( .I0(n23937), .I1(n23927), .I2(n23932), .I3(n23922), .S0(
        n26117), .S1(n26147), .ZN(n23943) );
  MUX41 U7819 ( .I0(n23772), .I1(n23773), .I2(n23774), .I3(n23775), .S0(
        n26090), .S1(n26093), .ZN(n23771) );
  MUX41 U7820 ( .I0(n23726), .I1(n23716), .I2(n23721), .I3(n23711), .S0(
        n26116), .S1(n26146), .ZN(n23773) );
  MUX41 U7821 ( .I0(n23706), .I1(n23696), .I2(n23701), .I3(n23691), .S0(
        n26116), .S1(n26146), .ZN(n23775) );
  MUX41 U7822 ( .I0(n23766), .I1(n23756), .I2(n23761), .I3(n23751), .S0(
        n26116), .S1(n26146), .ZN(n23772) );
  MUX41 U7823 ( .I0(n24627), .I1(n24628), .I2(n24629), .I3(n24630), .S0(
        n26088), .S1(raddr[6]), .ZN(n24626) );
  MUX41 U7824 ( .I0(n24561), .I1(n24551), .I2(n24556), .I3(n24546), .S0(
        n26119), .S1(n26149), .ZN(n24630) );
  MUX41 U7825 ( .I0(n24581), .I1(n24571), .I2(n24576), .I3(n24566), .S0(
        n26119), .S1(n26149), .ZN(n24628) );
  MUX41 U7826 ( .I0(n24621), .I1(n24611), .I2(n24616), .I3(n24606), .S0(
        n26119), .S1(n26149), .ZN(n24627) );
  MUX41 U7827 ( .I0(n24456), .I1(n24457), .I2(n24458), .I3(n24459), .S0(
        n26089), .S1(raddr[6]), .ZN(n24455) );
  MUX41 U7828 ( .I0(n24410), .I1(n24400), .I2(n24405), .I3(n24395), .S0(
        n26118), .S1(n26148), .ZN(n24457) );
  MUX41 U7829 ( .I0(n24390), .I1(n24380), .I2(n24385), .I3(n24375), .S0(
        n26118), .S1(n26148), .ZN(n24459) );
  MUX41 U7830 ( .I0(n24450), .I1(n24440), .I2(n24445), .I3(n24435), .S0(
        n26119), .S1(n26149), .ZN(n24456) );
  MUX41 U7831 ( .I0(n25311), .I1(n25312), .I2(n25313), .I3(n25314), .S0(
        n26088), .S1(n26094), .ZN(n25310) );
  MUX41 U7832 ( .I0(n25245), .I1(n25235), .I2(n25240), .I3(n25230), .S0(
        n26121), .S1(n26151), .ZN(n25314) );
  MUX41 U7833 ( .I0(n25265), .I1(n25255), .I2(n25260), .I3(n25250), .S0(
        n26122), .S1(n26152), .ZN(n25312) );
  MUX41 U7834 ( .I0(n25305), .I1(n25295), .I2(n25300), .I3(n25290), .S0(
        n26122), .S1(n26152), .ZN(n25311) );
  MUX41 U7835 ( .I0(n25140), .I1(n25141), .I2(n25142), .I3(n25143), .S0(
        n26089), .S1(n26094), .ZN(n25139) );
  MUX41 U7836 ( .I0(n25094), .I1(n25084), .I2(n25089), .I3(n25079), .S0(
        n26121), .S1(n26151), .ZN(n25141) );
  MUX41 U7837 ( .I0(n25074), .I1(n25064), .I2(n25069), .I3(n25059), .S0(
        n26121), .S1(n26151), .ZN(n25143) );
  MUX41 U7838 ( .I0(n25134), .I1(n25124), .I2(n25129), .I3(n25119), .S0(
        n26121), .S1(n26151), .ZN(n25140) );
  MUX41 U7839 ( .I0(n25995), .I1(n25996), .I2(n25997), .I3(n25998), .S0(
        n26088), .S1(n26094), .ZN(n25994) );
  MUX41 U7840 ( .I0(n25929), .I1(n25919), .I2(n25924), .I3(n25914), .S0(
        n26124), .S1(n26154), .ZN(n25998) );
  MUX41 U7841 ( .I0(n25949), .I1(n25939), .I2(n25944), .I3(n25934), .S0(
        n26124), .S1(n26154), .ZN(n25996) );
  MUX41 U7842 ( .I0(n25989), .I1(n25979), .I2(n25984), .I3(n25974), .S0(
        n26124), .S1(n26154), .ZN(n25995) );
  MUX41 U7843 ( .I0(n25824), .I1(n25825), .I2(n25826), .I3(n25827), .S0(
        n26090), .S1(n26094), .ZN(n25823) );
  MUX41 U7844 ( .I0(n25778), .I1(n25768), .I2(n25773), .I3(n25763), .S0(
        n26123), .S1(n26153), .ZN(n25825) );
  MUX41 U7845 ( .I0(n25758), .I1(n25748), .I2(n25753), .I3(n25743), .S0(
        n26123), .S1(n26153), .ZN(n25827) );
  MUX41 U7846 ( .I0(n25818), .I1(n25808), .I2(n25813), .I3(n25803), .S0(
        n26124), .S1(n26154), .ZN(n25824) );
  MUX41 U7847 ( .I0(n21207), .I1(n21208), .I2(n21209), .I3(n21210), .S0(
        n26088), .S1(raddr[6]), .ZN(n21206) );
  MUX41 U7848 ( .I0(n21141), .I1(n21131), .I2(n21136), .I3(n21126), .S0(
        n26107), .S1(n26137), .ZN(n21210) );
  MUX41 U7849 ( .I0(n21161), .I1(n21151), .I2(n21156), .I3(n21146), .S0(
        n26107), .S1(n26137), .ZN(n21208) );
  MUX41 U7850 ( .I0(n21201), .I1(n21191), .I2(n21196), .I3(n21186), .S0(
        n26107), .S1(n26137), .ZN(n21207) );
  MUX41 U7851 ( .I0(n21036), .I1(n21037), .I2(n21038), .I3(n21039), .S0(
        n26088), .S1(n26093), .ZN(n21035) );
  MUX41 U7852 ( .I0(n20990), .I1(n20980), .I2(n20985), .I3(n20975), .S0(
        n26106), .S1(n26136), .ZN(n21037) );
  MUX41 U7853 ( .I0(n20970), .I1(n20960), .I2(n20965), .I3(n20955), .S0(
        n26106), .S1(n26136), .ZN(n21039) );
  MUX41 U7854 ( .I0(n21030), .I1(n21020), .I2(n21025), .I3(n21015), .S0(
        n26106), .S1(n26136), .ZN(n21036) );
  MUX41 U7855 ( .I0(n20753), .I1(n20743), .I2(n20748), .I3(n20738), .S0(
        n26105), .S1(n26135), .ZN(n20781) );
  MUX41 U7856 ( .I0(n20739), .I1(n20740), .I2(n20741), .I3(n20742), .S0(
        n26196), .S1(n26314), .ZN(n20738) );
  MUX41 U7857 ( .I0(n20744), .I1(n20745), .I2(n20746), .I3(n20747), .S0(
        n26196), .S1(n26314), .ZN(n20743) );
  MUX41 U7858 ( .I0(n20754), .I1(n20755), .I2(n20756), .I3(n20757), .S0(
        n26196), .S1(n26314), .ZN(n20753) );
  MUX41 U7859 ( .I0(n20668), .I1(n20658), .I2(n20663), .I3(n20653), .S0(
        n26105), .S1(n26135), .ZN(n20696) );
  MUX41 U7860 ( .I0(n20654), .I1(n20655), .I2(n20656), .I3(n20657), .S0(
        n26194), .S1(n26312), .ZN(n20653) );
  MUX41 U7861 ( .I0(n20659), .I1(n20660), .I2(n20661), .I3(n20662), .S0(
        n26194), .S1(n26312), .ZN(n20658) );
  MUX41 U7862 ( .I0(n20669), .I1(n20670), .I2(n20671), .I3(n20672), .S0(
        n26195), .S1(n26313), .ZN(n20668) );
  MUX41 U7863 ( .I0(n21437), .I1(n21427), .I2(n21432), .I3(n21422), .S0(
        n26108), .S1(n26138), .ZN(n21465) );
  MUX41 U7864 ( .I0(n21423), .I1(n21424), .I2(n21425), .I3(n21426), .S0(
        n26205), .S1(n26323), .ZN(n21422) );
  MUX41 U7865 ( .I0(n21428), .I1(n21429), .I2(n21430), .I3(n21431), .S0(
        n26206), .S1(n26324), .ZN(n21427) );
  MUX41 U7866 ( .I0(n21438), .I1(n21439), .I2(n21440), .I3(n21441), .S0(
        n26206), .S1(n26324), .ZN(n21437) );
  MUX41 U7867 ( .I0(n21352), .I1(n21342), .I2(n21347), .I3(n21337), .S0(
        n26107), .S1(n26137), .ZN(n21380) );
  MUX41 U7868 ( .I0(n21338), .I1(n21339), .I2(n21340), .I3(n21341), .S0(
        n26204), .S1(n26322), .ZN(n21337) );
  MUX41 U7869 ( .I0(n21343), .I1(n21344), .I2(n21345), .I3(n21346), .S0(
        n26204), .S1(n26322), .ZN(n21342) );
  MUX41 U7870 ( .I0(n21353), .I1(n21354), .I2(n21355), .I3(n21356), .S0(
        n26204), .S1(n26322), .ZN(n21352) );
  MUX41 U7871 ( .I0(n22121), .I1(n22111), .I2(n22116), .I3(n22106), .S0(
        n26110), .S1(n26140), .ZN(n22149) );
  MUX41 U7872 ( .I0(n22107), .I1(n22108), .I2(n22109), .I3(n22110), .S0(
        n26215), .S1(n26333), .ZN(n22106) );
  MUX41 U7873 ( .I0(n22112), .I1(n22113), .I2(n22114), .I3(n22115), .S0(
        n26215), .S1(n26333), .ZN(n22111) );
  MUX41 U7874 ( .I0(n22122), .I1(n22123), .I2(n22124), .I3(n22125), .S0(
        n26216), .S1(n26334), .ZN(n22121) );
  MUX41 U7875 ( .I0(n22036), .I1(n22026), .I2(n22031), .I3(n22021), .S0(
        n26110), .S1(n26140), .ZN(n22064) );
  MUX41 U7876 ( .I0(n22022), .I1(n22023), .I2(n22024), .I3(n22025), .S0(
        n26214), .S1(n26332), .ZN(n22021) );
  MUX41 U7877 ( .I0(n22027), .I1(n22028), .I2(n22029), .I3(n22030), .S0(
        n26214), .S1(n26332), .ZN(n22026) );
  MUX41 U7878 ( .I0(n22037), .I1(n22038), .I2(n22039), .I3(n22040), .S0(
        n26214), .S1(n26332), .ZN(n22036) );
  MUX41 U7879 ( .I0(n22805), .I1(n22795), .I2(n22800), .I3(n22790), .S0(
        n26113), .S1(n26143), .ZN(n22833) );
  MUX41 U7880 ( .I0(n22791), .I1(n22792), .I2(n22793), .I3(n22794), .S0(
        n26225), .S1(n26343), .ZN(n22790) );
  MUX41 U7881 ( .I0(n22796), .I1(n22797), .I2(n22798), .I3(n22799), .S0(
        n26225), .S1(n26343), .ZN(n22795) );
  MUX41 U7882 ( .I0(n22806), .I1(n22807), .I2(n22808), .I3(n22809), .S0(
        n26225), .S1(n26343), .ZN(n22805) );
  MUX41 U7883 ( .I0(n22720), .I1(n22710), .I2(n22715), .I3(n22705), .S0(
        n26112), .S1(n26142), .ZN(n22748) );
  MUX41 U7884 ( .I0(n22706), .I1(n22707), .I2(n22708), .I3(n22709), .S0(
        n26224), .S1(n26342), .ZN(n22705) );
  MUX41 U7885 ( .I0(n22711), .I1(n22712), .I2(n22713), .I3(n22714), .S0(
        n26224), .S1(n26342), .ZN(n22710) );
  MUX41 U7886 ( .I0(n22721), .I1(n22722), .I2(n22723), .I3(n22724), .S0(
        n26224), .S1(n26342), .ZN(n22720) );
  MUX41 U7887 ( .I0(n23489), .I1(n23479), .I2(n23484), .I3(n23474), .S0(
        n26115), .S1(n26145), .ZN(n23517) );
  MUX41 U7888 ( .I0(n23475), .I1(n23476), .I2(n23477), .I3(n23478), .S0(
        n26235), .S1(n26353), .ZN(n23474) );
  MUX41 U7889 ( .I0(n23480), .I1(n23481), .I2(n23482), .I3(n23483), .S0(
        n26235), .S1(n26353), .ZN(n23479) );
  MUX41 U7890 ( .I0(n23490), .I1(n23491), .I2(n23492), .I3(n23493), .S0(
        n26235), .S1(n26353), .ZN(n23489) );
  MUX41 U7891 ( .I0(n23404), .I1(n23394), .I2(n23399), .I3(n23389), .S0(
        n26115), .S1(n26145), .ZN(n23432) );
  MUX41 U7892 ( .I0(n23390), .I1(n23391), .I2(n23392), .I3(n23393), .S0(
        n26234), .S1(n26352), .ZN(n23389) );
  MUX41 U7893 ( .I0(n23395), .I1(n23396), .I2(n23397), .I3(n23398), .S0(
        n26234), .S1(n26352), .ZN(n23394) );
  MUX41 U7894 ( .I0(n23405), .I1(n23406), .I2(n23407), .I3(n23408), .S0(
        n26234), .S1(n26352), .ZN(n23404) );
  MUX41 U7895 ( .I0(n24173), .I1(n24163), .I2(n24168), .I3(n24158), .S0(
        n26118), .S1(n26148), .ZN(n24201) );
  MUX41 U7896 ( .I0(n24159), .I1(n24160), .I2(n24161), .I3(n24162), .S0(
        n26245), .S1(n26363), .ZN(n24158) );
  MUX41 U7897 ( .I0(n24164), .I1(n24165), .I2(n24166), .I3(n24167), .S0(
        n26245), .S1(n26363), .ZN(n24163) );
  MUX41 U7898 ( .I0(n24174), .I1(n24175), .I2(n24176), .I3(n24177), .S0(
        n26245), .S1(n26363), .ZN(n24173) );
  MUX41 U7899 ( .I0(n24088), .I1(n24078), .I2(n24083), .I3(n24073), .S0(
        n26117), .S1(n26147), .ZN(n24116) );
  MUX41 U7900 ( .I0(n24074), .I1(n24075), .I2(n24076), .I3(n24077), .S0(
        n26244), .S1(n26362), .ZN(n24073) );
  MUX41 U7901 ( .I0(n24079), .I1(n24080), .I2(n24081), .I3(n24082), .S0(
        n26244), .S1(n26362), .ZN(n24078) );
  MUX41 U7902 ( .I0(n24089), .I1(n24090), .I2(n24091), .I3(n24092), .S0(
        n26244), .S1(n26362), .ZN(n24088) );
  MUX41 U7903 ( .I0(n24857), .I1(n24847), .I2(n24852), .I3(n24842), .S0(
        n26120), .S1(n26150), .ZN(n24885) );
  MUX41 U7904 ( .I0(n24843), .I1(n24844), .I2(n24845), .I3(n24846), .S0(
        n26255), .S1(n26373), .ZN(n24842) );
  MUX41 U7905 ( .I0(n24848), .I1(n24849), .I2(n24850), .I3(n24851), .S0(
        n26255), .S1(n26373), .ZN(n24847) );
  MUX41 U7906 ( .I0(n24858), .I1(n24859), .I2(n24860), .I3(n24861), .S0(
        n26255), .S1(n26373), .ZN(n24857) );
  MUX41 U7907 ( .I0(n24772), .I1(n24762), .I2(n24767), .I3(n24757), .S0(
        n26120), .S1(n26150), .ZN(n24800) );
  MUX41 U7908 ( .I0(n24758), .I1(n24759), .I2(n24760), .I3(n24761), .S0(
        n26253), .S1(n26371), .ZN(n24757) );
  MUX41 U7909 ( .I0(n24763), .I1(n24764), .I2(n24765), .I3(n24766), .S0(
        n26254), .S1(n26372), .ZN(n24762) );
  MUX41 U7910 ( .I0(n24773), .I1(n24774), .I2(n24775), .I3(n24776), .S0(
        n26254), .S1(n26372), .ZN(n24772) );
  MUX41 U7911 ( .I0(n25541), .I1(n25531), .I2(n25536), .I3(n25526), .S0(
        n26123), .S1(n26153), .ZN(n25569) );
  MUX41 U7912 ( .I0(n25527), .I1(n25528), .I2(n25529), .I3(n25530), .S0(
        n26265), .S1(n26383), .ZN(n25526) );
  MUX41 U7913 ( .I0(n25532), .I1(n25533), .I2(n25534), .I3(n25535), .S0(
        n26265), .S1(n26383), .ZN(n25531) );
  MUX41 U7914 ( .I0(n25542), .I1(n25543), .I2(n25544), .I3(n25545), .S0(
        n26265), .S1(n26383), .ZN(n25541) );
  MUX41 U7915 ( .I0(n25456), .I1(n25446), .I2(n25451), .I3(n25441), .S0(
        n26122), .S1(n26152), .ZN(n25484) );
  MUX41 U7916 ( .I0(n25442), .I1(n25443), .I2(n25444), .I3(n25445), .S0(
        n26263), .S1(n26381), .ZN(n25441) );
  MUX41 U7917 ( .I0(n25447), .I1(n25448), .I2(n25449), .I3(n25450), .S0(
        n26263), .S1(n26381), .ZN(n25446) );
  MUX41 U7918 ( .I0(n25457), .I1(n25458), .I2(n25459), .I3(n25460), .S0(
        n26264), .S1(n26382), .ZN(n25456) );
  MUX41 U7919 ( .I0(n21266), .I1(n21256), .I2(n21261), .I3(n21251), .S0(
        n26107), .S1(n26137), .ZN(n21294) );
  MUX41 U7920 ( .I0(n21252), .I1(n21253), .I2(n21254), .I3(n21255), .S0(
        n26203), .S1(n26321), .ZN(n21251) );
  MUX41 U7921 ( .I0(n21257), .I1(n21258), .I2(n21259), .I3(n21260), .S0(
        n26203), .S1(n26321), .ZN(n21256) );
  MUX41 U7922 ( .I0(n21267), .I1(n21268), .I2(n21269), .I3(n21270), .S0(
        n26203), .S1(n26321), .ZN(n21266) );
  MUX41 U7923 ( .I0(n21181), .I1(n21171), .I2(n21176), .I3(n21166), .S0(
        n26107), .S1(n26137), .ZN(n21209) );
  MUX41 U7924 ( .I0(n21167), .I1(n21168), .I2(n21169), .I3(n21170), .S0(
        n26202), .S1(n26320), .ZN(n21166) );
  MUX41 U7925 ( .I0(n21172), .I1(n21173), .I2(n21174), .I3(n21175), .S0(
        n26202), .S1(n26320), .ZN(n21171) );
  MUX41 U7926 ( .I0(n21182), .I1(n21183), .I2(n21184), .I3(n21185), .S0(
        n26202), .S1(n26320), .ZN(n21181) );
  MUX41 U7927 ( .I0(n20924), .I1(n20914), .I2(n20919), .I3(n20909), .S0(
        n26106), .S1(n26136), .ZN(n20952) );
  MUX41 U7928 ( .I0(n20910), .I1(n20911), .I2(n20912), .I3(n20913), .S0(
        n26198), .S1(n26316), .ZN(n20909) );
  MUX41 U7929 ( .I0(n20915), .I1(n20916), .I2(n20917), .I3(n20918), .S0(
        n26198), .S1(n26316), .ZN(n20914) );
  MUX41 U7930 ( .I0(n20925), .I1(n20926), .I2(n20927), .I3(n20928), .S0(
        n26198), .S1(n26316), .ZN(n20924) );
  MUX41 U7931 ( .I0(n20839), .I1(n20829), .I2(n20834), .I3(n20824), .S0(
        n26106), .S1(n26136), .ZN(n20867) );
  MUX41 U7932 ( .I0(n20825), .I1(n20826), .I2(n20827), .I3(n20828), .S0(
        n26197), .S1(n26315), .ZN(n20824) );
  MUX41 U7933 ( .I0(n20830), .I1(n20831), .I2(n20832), .I3(n20833), .S0(
        n26197), .S1(n26315), .ZN(n20829) );
  MUX41 U7934 ( .I0(n20840), .I1(n20841), .I2(n20842), .I3(n20843), .S0(
        n26197), .S1(n26315), .ZN(n20839) );
  MUX41 U7935 ( .I0(n21095), .I1(n21085), .I2(n21090), .I3(n21080), .S0(
        n26107), .S1(n26137), .ZN(n21123) );
  MUX41 U7936 ( .I0(n21081), .I1(n21082), .I2(n21083), .I3(n21084), .S0(
        n26201), .S1(n26319), .ZN(n21080) );
  MUX41 U7937 ( .I0(n21086), .I1(n21087), .I2(n21088), .I3(n21089), .S0(
        n26201), .S1(n26319), .ZN(n21085) );
  MUX41 U7938 ( .I0(n21096), .I1(n21097), .I2(n21098), .I3(n21099), .S0(
        n26201), .S1(n26319), .ZN(n21095) );
  MUX41 U7939 ( .I0(n21010), .I1(n21000), .I2(n21005), .I3(n20995), .S0(
        n26106), .S1(n26136), .ZN(n21038) );
  MUX41 U7940 ( .I0(n20996), .I1(n20997), .I2(n20998), .I3(n20999), .S0(
        n26199), .S1(n26317), .ZN(n20995) );
  MUX41 U7941 ( .I0(n21001), .I1(n21002), .I2(n21003), .I3(n21004), .S0(
        n26199), .S1(n26317), .ZN(n21000) );
  MUX41 U7942 ( .I0(n21011), .I1(n21012), .I2(n21013), .I3(n21014), .S0(
        n26200), .S1(n26318), .ZN(n21010) );
  MUX41 U7943 ( .I0(n21950), .I1(n21940), .I2(n21945), .I3(n21935), .S0(
        n26110), .S1(n26140), .ZN(n21978) );
  MUX41 U7944 ( .I0(n21936), .I1(n21937), .I2(n21938), .I3(n21939), .S0(
        n26213), .S1(n26331), .ZN(n21935) );
  MUX41 U7945 ( .I0(n21941), .I1(n21942), .I2(n21943), .I3(n21944), .S0(
        n26213), .S1(n26331), .ZN(n21940) );
  MUX41 U7946 ( .I0(n21951), .I1(n21952), .I2(n21953), .I3(n21954), .S0(
        n26213), .S1(n26331), .ZN(n21950) );
  MUX41 U7947 ( .I0(n21865), .I1(n21855), .I2(n21860), .I3(n21850), .S0(
        n26109), .S1(n26139), .ZN(n21893) );
  MUX41 U7948 ( .I0(n21851), .I1(n21852), .I2(n21853), .I3(n21854), .S0(
        n26212), .S1(n26330), .ZN(n21850) );
  MUX41 U7949 ( .I0(n21856), .I1(n21857), .I2(n21858), .I3(n21859), .S0(
        n26212), .S1(n26330), .ZN(n21855) );
  MUX41 U7950 ( .I0(n21866), .I1(n21867), .I2(n21868), .I3(n21869), .S0(
        n26212), .S1(n26330), .ZN(n21865) );
  MUX41 U7951 ( .I0(n21608), .I1(n21598), .I2(n21603), .I3(n21593), .S0(
        n26108), .S1(n26138), .ZN(n21636) );
  MUX41 U7952 ( .I0(n21594), .I1(n21595), .I2(n21596), .I3(n21597), .S0(
        n26208), .S1(n26326), .ZN(n21593) );
  MUX41 U7953 ( .I0(n21599), .I1(n21600), .I2(n21601), .I3(n21602), .S0(
        n26208), .S1(n26326), .ZN(n21598) );
  MUX41 U7954 ( .I0(n21609), .I1(n21610), .I2(n21611), .I3(n21612), .S0(
        n26208), .S1(n26326), .ZN(n21608) );
  MUX41 U7955 ( .I0(n21523), .I1(n21513), .I2(n21518), .I3(n21508), .S0(
        n26108), .S1(n26138), .ZN(n21551) );
  MUX41 U7956 ( .I0(n21509), .I1(n21510), .I2(n21511), .I3(n21512), .S0(
        n26207), .S1(n26325), .ZN(n21508) );
  MUX41 U7957 ( .I0(n21514), .I1(n21515), .I2(n21516), .I3(n21517), .S0(
        n26207), .S1(n26325), .ZN(n21513) );
  MUX41 U7958 ( .I0(n21524), .I1(n21525), .I2(n21526), .I3(n21527), .S0(
        n26207), .S1(n26325), .ZN(n21523) );
  MUX41 U7959 ( .I0(n21779), .I1(n21769), .I2(n21774), .I3(n21764), .S0(
        n26109), .S1(n26139), .ZN(n21807) );
  MUX41 U7960 ( .I0(n21765), .I1(n21766), .I2(n21767), .I3(n21768), .S0(
        n26210), .S1(n26328), .ZN(n21764) );
  MUX41 U7961 ( .I0(n21770), .I1(n21771), .I2(n21772), .I3(n21773), .S0(
        n26210), .S1(n26328), .ZN(n21769) );
  MUX41 U7962 ( .I0(n21780), .I1(n21781), .I2(n21782), .I3(n21783), .S0(
        n26211), .S1(n26329), .ZN(n21779) );
  MUX41 U7963 ( .I0(n21694), .I1(n21684), .I2(n21689), .I3(n21679), .S0(
        n26109), .S1(n26139), .ZN(n21722) );
  MUX41 U7964 ( .I0(n21680), .I1(n21681), .I2(n21682), .I3(n21683), .S0(
        n26209), .S1(n26327), .ZN(n21679) );
  MUX41 U7965 ( .I0(n21685), .I1(n21686), .I2(n21687), .I3(n21688), .S0(
        n26209), .S1(n26327), .ZN(n21684) );
  MUX41 U7966 ( .I0(n21695), .I1(n21696), .I2(n21697), .I3(n21698), .S0(
        n26209), .S1(n26327), .ZN(n21694) );
  MUX41 U7967 ( .I0(n22634), .I1(n22624), .I2(n22629), .I3(n22619), .S0(
        n26112), .S1(n26142), .ZN(n22662) );
  MUX41 U7968 ( .I0(n22620), .I1(n22621), .I2(n22622), .I3(n22623), .S0(
        n26223), .S1(n26341), .ZN(n22619) );
  MUX41 U7969 ( .I0(n22625), .I1(n22626), .I2(n22627), .I3(n22628), .S0(
        n26223), .S1(n26341), .ZN(n22624) );
  MUX41 U7970 ( .I0(n22635), .I1(n22636), .I2(n22637), .I3(n22638), .S0(
        n26223), .S1(n26341), .ZN(n22634) );
  MUX41 U7971 ( .I0(n22549), .I1(n22539), .I2(n22544), .I3(n22534), .S0(
        n26112), .S1(n26142), .ZN(n22577) );
  MUX41 U7972 ( .I0(n22535), .I1(n22536), .I2(n22537), .I3(n22538), .S0(
        n26221), .S1(n26339), .ZN(n22534) );
  MUX41 U7973 ( .I0(n22540), .I1(n22541), .I2(n22542), .I3(n22543), .S0(
        n26222), .S1(n26340), .ZN(n22539) );
  MUX41 U7974 ( .I0(n22550), .I1(n22551), .I2(n22552), .I3(n22553), .S0(
        n26222), .S1(n26340), .ZN(n22549) );
  MUX41 U7975 ( .I0(n22292), .I1(n22282), .I2(n22287), .I3(n22277), .S0(
        n26111), .S1(n26141), .ZN(n22320) );
  MUX41 U7976 ( .I0(n22278), .I1(n22279), .I2(n22280), .I3(n22281), .S0(
        n26218), .S1(n26336), .ZN(n22277) );
  MUX41 U7977 ( .I0(n22283), .I1(n22284), .I2(n22285), .I3(n22286), .S0(
        n26218), .S1(n26336), .ZN(n22282) );
  MUX41 U7978 ( .I0(n22293), .I1(n22294), .I2(n22295), .I3(n22296), .S0(
        n26218), .S1(n26336), .ZN(n22292) );
  MUX41 U7979 ( .I0(n22207), .I1(n22197), .I2(n22202), .I3(n22192), .S0(
        n26111), .S1(n26141), .ZN(n22235) );
  MUX41 U7980 ( .I0(n22193), .I1(n22194), .I2(n22195), .I3(n22196), .S0(
        n26217), .S1(n26335), .ZN(n22192) );
  MUX41 U7981 ( .I0(n22198), .I1(n22199), .I2(n22200), .I3(n22201), .S0(
        n26217), .S1(n26335), .ZN(n22197) );
  MUX41 U7982 ( .I0(n22208), .I1(n22209), .I2(n22210), .I3(n22211), .S0(
        n26217), .S1(n26335), .ZN(n22207) );
  MUX41 U7983 ( .I0(n22463), .I1(n22453), .I2(n22458), .I3(n22448), .S0(
        n26111), .S1(n26141), .ZN(n22491) );
  MUX41 U7984 ( .I0(n22449), .I1(n22450), .I2(n22451), .I3(n22452), .S0(
        n26220), .S1(n26338), .ZN(n22448) );
  MUX41 U7985 ( .I0(n22454), .I1(n22455), .I2(n22456), .I3(n22457), .S0(
        n26220), .S1(n26338), .ZN(n22453) );
  MUX41 U7986 ( .I0(n22464), .I1(n22465), .I2(n22466), .I3(n22467), .S0(
        n26220), .S1(n26338), .ZN(n22463) );
  MUX41 U7987 ( .I0(n22378), .I1(n22368), .I2(n22373), .I3(n22363), .S0(
        n26111), .S1(n26141), .ZN(n22406) );
  MUX41 U7988 ( .I0(n22364), .I1(n22365), .I2(n22366), .I3(n22367), .S0(
        n26219), .S1(n26337), .ZN(n22363) );
  MUX41 U7989 ( .I0(n22369), .I1(n22370), .I2(n22371), .I3(n22372), .S0(
        n26219), .S1(n26337), .ZN(n22368) );
  MUX41 U7990 ( .I0(n22379), .I1(n22380), .I2(n22381), .I3(n22382), .S0(
        n26219), .S1(n26337), .ZN(n22378) );
  MUX41 U7991 ( .I0(n23318), .I1(n23308), .I2(n23313), .I3(n23303), .S0(
        n26115), .S1(n26145), .ZN(n23346) );
  MUX41 U7992 ( .I0(n23304), .I1(n23305), .I2(n23306), .I3(n23307), .S0(
        n26233), .S1(n26351), .ZN(n23303) );
  MUX41 U7993 ( .I0(n23309), .I1(n23310), .I2(n23311), .I3(n23312), .S0(
        n26233), .S1(n26351), .ZN(n23308) );
  MUX41 U7994 ( .I0(n23319), .I1(n23320), .I2(n23321), .I3(n23322), .S0(
        n26233), .S1(n26351), .ZN(n23318) );
  MUX41 U7995 ( .I0(n23233), .I1(n23223), .I2(n23228), .I3(n23218), .S0(
        n26114), .S1(n26144), .ZN(n23261) );
  MUX41 U7996 ( .I0(n23219), .I1(n23220), .I2(n23221), .I3(n23222), .S0(
        n26231), .S1(n26349), .ZN(n23218) );
  MUX41 U7997 ( .I0(n23224), .I1(n23225), .I2(n23226), .I3(n23227), .S0(
        n26231), .S1(n26349), .ZN(n23223) );
  MUX41 U7998 ( .I0(n23234), .I1(n23235), .I2(n23236), .I3(n23237), .S0(
        n26232), .S1(n26350), .ZN(n23233) );
  MUX41 U7999 ( .I0(n22976), .I1(n22966), .I2(n22971), .I3(n22961), .S0(
        n26113), .S1(n26143), .ZN(n23004) );
  MUX41 U8000 ( .I0(n22962), .I1(n22963), .I2(n22964), .I3(n22965), .S0(
        n26228), .S1(n26346), .ZN(n22961) );
  MUX41 U8001 ( .I0(n22967), .I1(n22968), .I2(n22969), .I3(n22970), .S0(
        n26228), .S1(n26346), .ZN(n22966) );
  MUX41 U8002 ( .I0(n22977), .I1(n22978), .I2(n22979), .I3(n22980), .S0(
        n26228), .S1(n26346), .ZN(n22976) );
  MUX41 U8003 ( .I0(n22891), .I1(n22881), .I2(n22886), .I3(n22876), .S0(
        n26113), .S1(n26143), .ZN(n22919) );
  MUX41 U8004 ( .I0(n22877), .I1(n22878), .I2(n22879), .I3(n22880), .S0(
        n26226), .S1(n26344), .ZN(n22876) );
  MUX41 U8005 ( .I0(n22882), .I1(n22883), .I2(n22884), .I3(n22885), .S0(
        n26226), .S1(n26344), .ZN(n22881) );
  MUX41 U8006 ( .I0(n22892), .I1(n22893), .I2(n22894), .I3(n22895), .S0(
        n26227), .S1(n26345), .ZN(n22891) );
  MUX41 U8007 ( .I0(n23147), .I1(n23137), .I2(n23142), .I3(n23132), .S0(
        n26114), .S1(n26144), .ZN(n23175) );
  MUX41 U8008 ( .I0(n23133), .I1(n23134), .I2(n23135), .I3(n23136), .S0(
        n26230), .S1(n26348), .ZN(n23132) );
  MUX41 U8009 ( .I0(n23138), .I1(n23139), .I2(n23140), .I3(n23141), .S0(
        n26230), .S1(n26348), .ZN(n23137) );
  MUX41 U8010 ( .I0(n23148), .I1(n23149), .I2(n23150), .I3(n23151), .S0(
        n26230), .S1(n26348), .ZN(n23147) );
  MUX41 U8011 ( .I0(n23062), .I1(n23052), .I2(n23057), .I3(n23047), .S0(
        n26114), .S1(n26144), .ZN(n23090) );
  MUX41 U8012 ( .I0(n23048), .I1(n23049), .I2(n23050), .I3(n23051), .S0(
        n26229), .S1(n26347), .ZN(n23047) );
  MUX41 U8013 ( .I0(n23053), .I1(n23054), .I2(n23055), .I3(n23056), .S0(
        n26229), .S1(n26347), .ZN(n23052) );
  MUX41 U8014 ( .I0(n23063), .I1(n23064), .I2(n23065), .I3(n23066), .S0(
        n26229), .S1(n26347), .ZN(n23062) );
  MUX41 U8015 ( .I0(n24002), .I1(n23992), .I2(n23997), .I3(n23987), .S0(
        n26117), .S1(n26147), .ZN(n24030) );
  MUX41 U8016 ( .I0(n23988), .I1(n23989), .I2(n23990), .I3(n23991), .S0(
        n26242), .S1(n26360), .ZN(n23987) );
  MUX41 U8017 ( .I0(n23993), .I1(n23994), .I2(n23995), .I3(n23996), .S0(
        n26242), .S1(n26360), .ZN(n23992) );
  MUX41 U8018 ( .I0(n24003), .I1(n24004), .I2(n24005), .I3(n24006), .S0(
        n26243), .S1(n26361), .ZN(n24002) );
  MUX41 U8019 ( .I0(n23917), .I1(n23907), .I2(n23912), .I3(n23902), .S0(
        n26117), .S1(n26147), .ZN(n23945) );
  MUX41 U8020 ( .I0(n23903), .I1(n23904), .I2(n23905), .I3(n23906), .S0(
        n26241), .S1(n26359), .ZN(n23902) );
  MUX41 U8021 ( .I0(n23908), .I1(n23909), .I2(n23910), .I3(n23911), .S0(
        n26241), .S1(n26359), .ZN(n23907) );
  MUX41 U8022 ( .I0(n23918), .I1(n23919), .I2(n23920), .I3(n23921), .S0(
        n26241), .S1(n26359), .ZN(n23917) );
  MUX41 U8023 ( .I0(n23660), .I1(n23650), .I2(n23655), .I3(n23645), .S0(
        n26116), .S1(n26146), .ZN(n23688) );
  MUX41 U8024 ( .I0(n23646), .I1(n23647), .I2(n23648), .I3(n23649), .S0(
        n26237), .S1(n26355), .ZN(n23645) );
  MUX41 U8025 ( .I0(n23651), .I1(n23652), .I2(n23653), .I3(n23654), .S0(
        n26238), .S1(n26356), .ZN(n23650) );
  MUX41 U8026 ( .I0(n23661), .I1(n23662), .I2(n23663), .I3(n23664), .S0(
        n26238), .S1(n26356), .ZN(n23660) );
  MUX41 U8027 ( .I0(n23575), .I1(n23565), .I2(n23570), .I3(n23560), .S0(
        n26115), .S1(n26145), .ZN(n23603) );
  MUX41 U8028 ( .I0(n23561), .I1(n23562), .I2(n23563), .I3(n23564), .S0(
        n26236), .S1(n26354), .ZN(n23560) );
  MUX41 U8029 ( .I0(n23566), .I1(n23567), .I2(n23568), .I3(n23569), .S0(
        n26236), .S1(n26354), .ZN(n23565) );
  MUX41 U8030 ( .I0(n23576), .I1(n23577), .I2(n23578), .I3(n23579), .S0(
        n26236), .S1(n26354), .ZN(n23575) );
  MUX41 U8031 ( .I0(n23831), .I1(n23821), .I2(n23826), .I3(n23816), .S0(
        n26116), .S1(n26146), .ZN(n23859) );
  MUX41 U8032 ( .I0(n23817), .I1(n23818), .I2(n23819), .I3(n23820), .S0(
        n26240), .S1(n26358), .ZN(n23816) );
  MUX41 U8033 ( .I0(n23822), .I1(n23823), .I2(n23824), .I3(n23825), .S0(
        n26240), .S1(n26358), .ZN(n23821) );
  MUX41 U8034 ( .I0(n23832), .I1(n23833), .I2(n23834), .I3(n23835), .S0(
        n26240), .S1(n26358), .ZN(n23831) );
  MUX41 U8035 ( .I0(n23746), .I1(n23736), .I2(n23741), .I3(n23731), .S0(
        n26116), .S1(n26146), .ZN(n23774) );
  MUX41 U8036 ( .I0(n23732), .I1(n23733), .I2(n23734), .I3(n23735), .S0(
        n26239), .S1(n26357), .ZN(n23731) );
  MUX41 U8037 ( .I0(n23737), .I1(n23738), .I2(n23739), .I3(n23740), .S0(
        n26239), .S1(n26357), .ZN(n23736) );
  MUX41 U8038 ( .I0(n23747), .I1(n23748), .I2(n23749), .I3(n23750), .S0(
        n26239), .S1(n26357), .ZN(n23746) );
  MUX41 U8039 ( .I0(n24686), .I1(n24676), .I2(n24681), .I3(n24671), .S0(
        n26119), .S1(n26149), .ZN(n24714) );
  MUX41 U8040 ( .I0(n24672), .I1(n24673), .I2(n24674), .I3(n24675), .S0(
        n26252), .S1(n26370), .ZN(n24671) );
  MUX41 U8041 ( .I0(n24677), .I1(n24678), .I2(n24679), .I3(n24680), .S0(
        n26252), .S1(n26370), .ZN(n24676) );
  MUX41 U8042 ( .I0(n24687), .I1(n24688), .I2(n24689), .I3(n24690), .S0(
        n26252), .S1(n26370), .ZN(n24686) );
  MUX41 U8043 ( .I0(n24601), .I1(n24591), .I2(n24596), .I3(n24586), .S0(
        n26119), .S1(n26149), .ZN(n24629) );
  MUX41 U8044 ( .I0(n24587), .I1(n24588), .I2(n24589), .I3(n24590), .S0(
        n26251), .S1(n26369), .ZN(n24586) );
  MUX41 U8045 ( .I0(n24592), .I1(n24593), .I2(n24594), .I3(n24595), .S0(
        n26251), .S1(n26369), .ZN(n24591) );
  MUX41 U8046 ( .I0(n24602), .I1(n24603), .I2(n24604), .I3(n24605), .S0(
        n26251), .S1(n26369), .ZN(n24601) );
  MUX41 U8047 ( .I0(n24344), .I1(n24334), .I2(n24339), .I3(n24329), .S0(
        n26118), .S1(n26148), .ZN(n24372) );
  MUX41 U8048 ( .I0(n24330), .I1(n24331), .I2(n24332), .I3(n24333), .S0(
        n26247), .S1(n26365), .ZN(n24329) );
  MUX41 U8049 ( .I0(n24335), .I1(n24336), .I2(n24337), .I3(n24338), .S0(
        n26247), .S1(n26365), .ZN(n24334) );
  MUX41 U8050 ( .I0(n24345), .I1(n24346), .I2(n24347), .I3(n24348), .S0(
        n26248), .S1(n26366), .ZN(n24344) );
  MUX41 U8051 ( .I0(n24259), .I1(n24249), .I2(n24254), .I3(n24244), .S0(
        n26118), .S1(n26148), .ZN(n24287) );
  MUX41 U8052 ( .I0(n24245), .I1(n24246), .I2(n24247), .I3(n24248), .S0(
        n26246), .S1(n26364), .ZN(n24244) );
  MUX41 U8053 ( .I0(n24250), .I1(n24251), .I2(n24252), .I3(n24253), .S0(
        n26246), .S1(n26364), .ZN(n24249) );
  MUX41 U8054 ( .I0(n24260), .I1(n24261), .I2(n24262), .I3(n24263), .S0(
        n26246), .S1(n26364), .ZN(n24259) );
  MUX41 U8055 ( .I0(n24515), .I1(n24505), .I2(n24510), .I3(n24500), .S0(
        n26119), .S1(n26149), .ZN(n24543) );
  MUX41 U8056 ( .I0(n24501), .I1(n24502), .I2(n24503), .I3(n24504), .S0(
        n26250), .S1(n26368), .ZN(n24500) );
  MUX41 U8057 ( .I0(n24506), .I1(n24507), .I2(n24508), .I3(n24509), .S0(
        n26250), .S1(n26368), .ZN(n24505) );
  MUX41 U8058 ( .I0(n24516), .I1(n24517), .I2(n24518), .I3(n24519), .S0(
        n26250), .S1(n26368), .ZN(n24515) );
  MUX41 U8059 ( .I0(n24430), .I1(n24420), .I2(n24425), .I3(n24415), .S0(
        n26119), .S1(n26149), .ZN(n24458) );
  MUX41 U8060 ( .I0(n24416), .I1(n24417), .I2(n24418), .I3(n24419), .S0(
        n26249), .S1(n26367), .ZN(n24415) );
  MUX41 U8061 ( .I0(n24421), .I1(n24422), .I2(n24423), .I3(n24424), .S0(
        n26249), .S1(n26367), .ZN(n24420) );
  MUX41 U8062 ( .I0(n24431), .I1(n24432), .I2(n24433), .I3(n24434), .S0(
        n26249), .S1(n26367), .ZN(n24430) );
  MUX41 U8063 ( .I0(n25370), .I1(n25360), .I2(n25365), .I3(n25355), .S0(
        n26122), .S1(n26152), .ZN(n25398) );
  MUX41 U8064 ( .I0(n25356), .I1(n25357), .I2(n25358), .I3(n25359), .S0(
        n26262), .S1(n26380), .ZN(n25355) );
  MUX41 U8065 ( .I0(n25361), .I1(n25362), .I2(n25363), .I3(n25364), .S0(
        n26262), .S1(n26380), .ZN(n25360) );
  MUX41 U8066 ( .I0(n25371), .I1(n25372), .I2(n25373), .I3(n25374), .S0(
        n26262), .S1(n26380), .ZN(n25370) );
  MUX41 U8067 ( .I0(n25285), .I1(n25275), .I2(n25280), .I3(n25270), .S0(
        n26122), .S1(n26152), .ZN(n25313) );
  MUX41 U8068 ( .I0(n25271), .I1(n25272), .I2(n25273), .I3(n25274), .S0(
        n26261), .S1(n26379), .ZN(n25270) );
  MUX41 U8069 ( .I0(n25276), .I1(n25277), .I2(n25278), .I3(n25279), .S0(
        n26261), .S1(n26379), .ZN(n25275) );
  MUX41 U8070 ( .I0(n25286), .I1(n25287), .I2(n25288), .I3(n25289), .S0(
        n26261), .S1(n26379), .ZN(n25285) );
  MUX41 U8071 ( .I0(n25028), .I1(n25018), .I2(n25023), .I3(n25013), .S0(
        n26121), .S1(n26151), .ZN(n25056) );
  MUX41 U8072 ( .I0(n25014), .I1(n25015), .I2(n25016), .I3(n25017), .S0(
        n26257), .S1(n26375), .ZN(n25013) );
  MUX41 U8073 ( .I0(n25019), .I1(n25020), .I2(n25021), .I3(n25022), .S0(
        n26257), .S1(n26375), .ZN(n25018) );
  MUX41 U8074 ( .I0(n25029), .I1(n25030), .I2(n25031), .I3(n25032), .S0(
        n26257), .S1(n26375), .ZN(n25028) );
  MUX41 U8075 ( .I0(n24943), .I1(n24933), .I2(n24938), .I3(n24928), .S0(
        n26120), .S1(n26150), .ZN(n24971) );
  MUX41 U8076 ( .I0(n24929), .I1(n24930), .I2(n24931), .I3(n24932), .S0(
        n26256), .S1(n26374), .ZN(n24928) );
  MUX41 U8077 ( .I0(n24934), .I1(n24935), .I2(n24936), .I3(n24937), .S0(
        n26256), .S1(n26374), .ZN(n24933) );
  MUX41 U8078 ( .I0(n24944), .I1(n24945), .I2(n24946), .I3(n24947), .S0(
        n26256), .S1(n26374), .ZN(n24943) );
  MUX41 U8079 ( .I0(n25199), .I1(n25189), .I2(n25194), .I3(n25184), .S0(
        n26121), .S1(n26151), .ZN(n25227) );
  MUX41 U8080 ( .I0(n25185), .I1(n25186), .I2(n25187), .I3(n25188), .S0(
        n26260), .S1(n26378), .ZN(n25184) );
  MUX41 U8081 ( .I0(n25190), .I1(n25191), .I2(n25192), .I3(n25193), .S0(
        n26260), .S1(n26378), .ZN(n25189) );
  MUX41 U8082 ( .I0(n25200), .I1(n25201), .I2(n25202), .I3(n25203), .S0(
        n26260), .S1(n26378), .ZN(n25199) );
  MUX41 U8083 ( .I0(n25114), .I1(n25104), .I2(n25109), .I3(n25099), .S0(
        n26121), .S1(n26151), .ZN(n25142) );
  MUX41 U8084 ( .I0(n25100), .I1(n25101), .I2(n25102), .I3(n25103), .S0(
        n26258), .S1(n26376), .ZN(n25099) );
  MUX41 U8085 ( .I0(n25105), .I1(n25106), .I2(n25107), .I3(n25108), .S0(
        n26258), .S1(n26376), .ZN(n25104) );
  MUX41 U8086 ( .I0(n25115), .I1(n25116), .I2(n25117), .I3(n25118), .S0(
        n26259), .S1(n26377), .ZN(n25114) );
  MUX41 U8087 ( .I0(n26054), .I1(n26044), .I2(n26049), .I3(n26039), .S0(
        n26124), .S1(n26154), .ZN(n26082) );
  MUX41 U8088 ( .I0(n26040), .I1(n26041), .I2(n26042), .I3(n26043), .S0(
        n26272), .S1(n26390), .ZN(n26039) );
  MUX41 U8089 ( .I0(n26045), .I1(n26046), .I2(n26047), .I3(n26048), .S0(
        n26272), .S1(n26390), .ZN(n26044) );
  MUX41 U8090 ( .I0(n26055), .I1(n26056), .I2(n26057), .I3(n26058), .S0(
        n26272), .S1(n26390), .ZN(n26054) );
  MUX41 U8091 ( .I0(n25969), .I1(n25959), .I2(n25964), .I3(n25954), .S0(
        n26124), .S1(n26154), .ZN(n25997) );
  MUX41 U8092 ( .I0(n25955), .I1(n25956), .I2(n25957), .I3(n25958), .S0(
        n26271), .S1(n26389), .ZN(n25954) );
  MUX41 U8093 ( .I0(n25960), .I1(n25961), .I2(n25962), .I3(n25963), .S0(
        n26271), .S1(n26389), .ZN(n25959) );
  MUX41 U8094 ( .I0(n25970), .I1(n25971), .I2(n25972), .I3(n25973), .S0(
        n26271), .S1(n26389), .ZN(n25969) );
  MUX41 U8095 ( .I0(n25712), .I1(n25702), .I2(n25707), .I3(n25697), .S0(
        n26123), .S1(n26153), .ZN(n25740) );
  MUX41 U8096 ( .I0(n25698), .I1(n25699), .I2(n25700), .I3(n25701), .S0(
        n26267), .S1(n26385), .ZN(n25697) );
  MUX41 U8097 ( .I0(n25703), .I1(n25704), .I2(n25705), .I3(n25706), .S0(
        n26267), .S1(n26385), .ZN(n25702) );
  MUX41 U8098 ( .I0(n25713), .I1(n25714), .I2(n25715), .I3(n25716), .S0(
        n26267), .S1(n26385), .ZN(n25712) );
  MUX41 U8099 ( .I0(n25627), .I1(n25617), .I2(n25622), .I3(n25612), .S0(
        n26123), .S1(n26153), .ZN(n25655) );
  MUX41 U8100 ( .I0(n25613), .I1(n25614), .I2(n25615), .I3(n25616), .S0(
        n26266), .S1(n26384), .ZN(n25612) );
  MUX41 U8101 ( .I0(n25618), .I1(n25619), .I2(n25620), .I3(n25621), .S0(
        n26266), .S1(n26384), .ZN(n25617) );
  MUX41 U8102 ( .I0(n25628), .I1(n25629), .I2(n25630), .I3(n25631), .S0(
        n26266), .S1(n26384), .ZN(n25627) );
  MUX41 U8103 ( .I0(n25883), .I1(n25873), .I2(n25878), .I3(n25868), .S0(
        n26124), .S1(n26154), .ZN(n25911) );
  MUX41 U8104 ( .I0(n25869), .I1(n25870), .I2(n25871), .I3(n25872), .S0(
        n26269), .S1(n26387), .ZN(n25868) );
  MUX41 U8105 ( .I0(n25874), .I1(n25875), .I2(n25876), .I3(n25877), .S0(
        n26270), .S1(n26388), .ZN(n25873) );
  MUX41 U8106 ( .I0(n25884), .I1(n25885), .I2(n25886), .I3(n25887), .S0(
        n26270), .S1(n26388), .ZN(n25883) );
  MUX41 U8107 ( .I0(n25798), .I1(n25788), .I2(n25793), .I3(n25783), .S0(
        n26123), .S1(n26153), .ZN(n25826) );
  MUX41 U8108 ( .I0(n25784), .I1(n25785), .I2(n25786), .I3(n25787), .S0(
        n26268), .S1(n26386), .ZN(n25783) );
  MUX41 U8109 ( .I0(n25789), .I1(n25790), .I2(n25791), .I3(n25792), .S0(
        n26268), .S1(n26386), .ZN(n25788) );
  MUX41 U8110 ( .I0(n25799), .I1(n25800), .I2(n25801), .I3(n25802), .S0(
        n26268), .S1(n26386), .ZN(n25798) );
  MUX41 U8111 ( .I0(n22318), .I1(n22319), .I2(n22320), .I3(n22321), .S0(
        n26089), .S1(n26093), .ZN(n22317) );
  MUX41 U8112 ( .I0(n22272), .I1(n22262), .I2(n22267), .I3(n22257), .S0(
        n26111), .S1(n26141), .ZN(n22319) );
  MUX41 U8113 ( .I0(n22252), .I1(n22242), .I2(n22247), .I3(n22237), .S0(
        n26111), .S1(n26141), .ZN(n22321) );
  MUX41 U8114 ( .I0(n22312), .I1(n22302), .I2(n22307), .I3(n22297), .S0(
        n26111), .S1(n26141), .ZN(n22318) );
  MUX41 U8115 ( .I0(n23002), .I1(n23003), .I2(n23004), .I3(n23005), .S0(
        n26090), .S1(n26093), .ZN(n23001) );
  MUX41 U8116 ( .I0(n22956), .I1(n22946), .I2(n22951), .I3(n22941), .S0(
        n26113), .S1(n26143), .ZN(n23003) );
  MUX41 U8117 ( .I0(n22936), .I1(n22926), .I2(n22931), .I3(n22921), .S0(
        n26113), .S1(n26143), .ZN(n23005) );
  MUX41 U8118 ( .I0(n22996), .I1(n22986), .I2(n22991), .I3(n22981), .S0(
        n26113), .S1(n26143), .ZN(n23002) );
  MUX41 U8119 ( .I0(n23686), .I1(n23687), .I2(n23688), .I3(n23689), .S0(
        n26090), .S1(n26093), .ZN(n23685) );
  MUX41 U8120 ( .I0(n23640), .I1(n23630), .I2(n23635), .I3(n23625), .S0(
        n26116), .S1(n26146), .ZN(n23687) );
  MUX41 U8121 ( .I0(n23620), .I1(n23610), .I2(n23615), .I3(n23605), .S0(
        n26116), .S1(n26146), .ZN(n23689) );
  MUX41 U8122 ( .I0(n23680), .I1(n23670), .I2(n23675), .I3(n23665), .S0(
        n26116), .S1(n26146), .ZN(n23686) );
  MUX41 U8123 ( .I0(n24370), .I1(n24371), .I2(n24372), .I3(n24373), .S0(
        n26088), .S1(raddr[6]), .ZN(n24369) );
  MUX41 U8124 ( .I0(n24324), .I1(n24314), .I2(n24319), .I3(n24309), .S0(
        n26118), .S1(n26148), .ZN(n24371) );
  MUX41 U8125 ( .I0(n24304), .I1(n24294), .I2(n24299), .I3(n24289), .S0(
        n26118), .S1(n26148), .ZN(n24373) );
  MUX41 U8126 ( .I0(n24364), .I1(n24354), .I2(n24359), .I3(n24349), .S0(
        n26118), .S1(n26148), .ZN(n24370) );
  MUX41 U8127 ( .I0(n25054), .I1(n25055), .I2(n25056), .I3(n25057), .S0(
        n26089), .S1(n26094), .ZN(n25053) );
  MUX41 U8128 ( .I0(n25008), .I1(n24998), .I2(n25003), .I3(n24993), .S0(
        n26121), .S1(n26151), .ZN(n25055) );
  MUX41 U8129 ( .I0(n24988), .I1(n24978), .I2(n24983), .I3(n24973), .S0(
        n26121), .S1(n26151), .ZN(n25057) );
  MUX41 U8130 ( .I0(n25048), .I1(n25038), .I2(n25043), .I3(n25033), .S0(
        n26121), .S1(n26151), .ZN(n25054) );
  MUX41 U8131 ( .I0(n25738), .I1(n25739), .I2(n25740), .I3(n25741), .S0(
        n26090), .S1(n26094), .ZN(n25737) );
  MUX41 U8132 ( .I0(n25692), .I1(n25682), .I2(n25687), .I3(n25677), .S0(
        n26123), .S1(n26153), .ZN(n25739) );
  MUX41 U8133 ( .I0(n25672), .I1(n25662), .I2(n25667), .I3(n25657), .S0(
        n26123), .S1(n26153), .ZN(n25741) );
  MUX41 U8134 ( .I0(n25732), .I1(n25722), .I2(n25727), .I3(n25717), .S0(
        n26123), .S1(n26153), .ZN(n25738) );
  MUX41 U8135 ( .I0(n20950), .I1(n20951), .I2(n20952), .I3(n20953), .S0(
        n26088), .S1(n26094), .ZN(n20949) );
  MUX41 U8136 ( .I0(n20904), .I1(n20894), .I2(n20899), .I3(n20889), .S0(
        n26106), .S1(n26136), .ZN(n20951) );
  MUX41 U8137 ( .I0(n20884), .I1(n20874), .I2(n20879), .I3(n20869), .S0(
        n26106), .S1(n26136), .ZN(n20953) );
  MUX41 U8138 ( .I0(n20944), .I1(n20934), .I2(n20939), .I3(n20929), .S0(
        n26106), .S1(n26136), .ZN(n20950) );
  MUX41 U8139 ( .I0(n21634), .I1(n21635), .I2(n21636), .I3(n21637), .S0(
        n26088), .S1(n26094), .ZN(n21633) );
  MUX41 U8140 ( .I0(n21588), .I1(n21578), .I2(n21583), .I3(n21573), .S0(
        n26108), .S1(n26138), .ZN(n21635) );
  MUX41 U8141 ( .I0(n21568), .I1(n21558), .I2(n21563), .I3(n21553), .S0(
        n26108), .S1(n26138), .ZN(n21637) );
  MUX41 U8142 ( .I0(n21628), .I1(n21618), .I2(n21623), .I3(n21613), .S0(
        n26108), .S1(n26138), .ZN(n21634) );
  MUX41 U8143 ( .I0(n21976), .I1(n21977), .I2(n21978), .I3(n21979), .S0(
        n26089), .S1(n26094), .ZN(n21975) );
  MUX41 U8144 ( .I0(n21910), .I1(n21900), .I2(n21905), .I3(n21895), .S0(
        n26109), .S1(n26139), .ZN(n21979) );
  MUX41 U8145 ( .I0(n21930), .I1(n21920), .I2(n21925), .I3(n21915), .S0(
        n26110), .S1(n26140), .ZN(n21977) );
  MUX41 U8146 ( .I0(n21970), .I1(n21960), .I2(n21965), .I3(n21955), .S0(
        n26110), .S1(n26140), .ZN(n21976) );
  MUX41 U8147 ( .I0(n21805), .I1(n21806), .I2(n21807), .I3(n21808), .S0(
        n26089), .S1(n26094), .ZN(n21804) );
  MUX41 U8148 ( .I0(n21759), .I1(n21749), .I2(n21754), .I3(n21744), .S0(
        n26109), .S1(n26139), .ZN(n21806) );
  MUX41 U8149 ( .I0(n21739), .I1(n21729), .I2(n21734), .I3(n21724), .S0(
        n26109), .S1(n26139), .ZN(n21808) );
  MUX41 U8150 ( .I0(n21799), .I1(n21789), .I2(n21794), .I3(n21784), .S0(
        n26109), .S1(n26139), .ZN(n21805) );
  MUX41 U8151 ( .I0(n22660), .I1(n22661), .I2(n22662), .I3(n22663), .S0(
        n26089), .S1(n26094), .ZN(n22659) );
  MUX41 U8152 ( .I0(n22594), .I1(n22584), .I2(n22589), .I3(n22579), .S0(
        n26112), .S1(n26142), .ZN(n22663) );
  MUX41 U8153 ( .I0(n22614), .I1(n22604), .I2(n22609), .I3(n22599), .S0(
        n26112), .S1(n26142), .ZN(n22661) );
  MUX41 U8154 ( .I0(n22654), .I1(n22644), .I2(n22649), .I3(n22639), .S0(
        n26112), .S1(n26142), .ZN(n22660) );
  MUX41 U8155 ( .I0(n22489), .I1(n22490), .I2(n22491), .I3(n22492), .S0(
        n26089), .S1(n26093), .ZN(n22488) );
  MUX41 U8156 ( .I0(n22443), .I1(n22433), .I2(n22438), .I3(n22428), .S0(
        n26111), .S1(n26141), .ZN(n22490) );
  MUX41 U8157 ( .I0(n22423), .I1(n22413), .I2(n22418), .I3(n22408), .S0(
        n26111), .S1(n26141), .ZN(n22492) );
  MUX41 U8158 ( .I0(n22483), .I1(n22473), .I2(n22478), .I3(n22468), .S0(
        n26112), .S1(n26142), .ZN(n22489) );
  MUX41 U8159 ( .I0(n23344), .I1(n23345), .I2(n23346), .I3(n23347), .S0(
        n26090), .S1(n26093), .ZN(n23343) );
  MUX41 U8160 ( .I0(n23278), .I1(n23268), .I2(n23273), .I3(n23263), .S0(
        n26114), .S1(n26144), .ZN(n23347) );
  MUX41 U8161 ( .I0(n23298), .I1(n23288), .I2(n23293), .I3(n23283), .S0(
        n26114), .S1(n26144), .ZN(n23345) );
  MUX41 U8162 ( .I0(n23338), .I1(n23328), .I2(n23333), .I3(n23323), .S0(
        n26115), .S1(n26145), .ZN(n23344) );
  MUX41 U8163 ( .I0(n23173), .I1(n23174), .I2(n23175), .I3(n23176), .S0(
        n26090), .S1(n26093), .ZN(n23172) );
  MUX41 U8164 ( .I0(n23127), .I1(n23117), .I2(n23122), .I3(n23112), .S0(
        n26114), .S1(n26144), .ZN(n23174) );
  MUX41 U8165 ( .I0(n23107), .I1(n23097), .I2(n23102), .I3(n23092), .S0(
        n26114), .S1(n26144), .ZN(n23176) );
  MUX41 U8166 ( .I0(n23167), .I1(n23157), .I2(n23162), .I3(n23152), .S0(
        n26114), .S1(n26144), .ZN(n23173) );
  MUX41 U8167 ( .I0(n24028), .I1(n24029), .I2(n24030), .I3(n24031), .S0(
        raddr[7]), .S1(raddr[6]), .ZN(n24027) );
  MUX41 U8168 ( .I0(n23962), .I1(n23952), .I2(n23957), .I3(n23947), .S0(
        n26117), .S1(n26147), .ZN(n24031) );
  MUX41 U8169 ( .I0(n23982), .I1(n23972), .I2(n23977), .I3(n23967), .S0(
        n26117), .S1(n26147), .ZN(n24029) );
  MUX41 U8170 ( .I0(n24022), .I1(n24012), .I2(n24017), .I3(n24007), .S0(
        n26117), .S1(n26147), .ZN(n24028) );
  MUX41 U8171 ( .I0(n23857), .I1(n23858), .I2(n23859), .I3(n23860), .S0(
        n26090), .S1(n26093), .ZN(n23856) );
  MUX41 U8172 ( .I0(n23811), .I1(n23801), .I2(n23806), .I3(n23796), .S0(
        n26116), .S1(n26146), .ZN(n23858) );
  MUX41 U8173 ( .I0(n23791), .I1(n23781), .I2(n23786), .I3(n23776), .S0(
        n26116), .S1(n26146), .ZN(n23860) );
  MUX41 U8174 ( .I0(n23851), .I1(n23841), .I2(n23846), .I3(n23836), .S0(
        n26116), .S1(n26146), .ZN(n23857) );
  MUX41 U8175 ( .I0(n24712), .I1(n24713), .I2(n24714), .I3(n24715), .S0(
        raddr[7]), .S1(raddr[6]), .ZN(n24711) );
  MUX41 U8176 ( .I0(n24646), .I1(n24636), .I2(n24641), .I3(n24631), .S0(
        n26119), .S1(n26149), .ZN(n24715) );
  MUX41 U8177 ( .I0(n24666), .I1(n24656), .I2(n24661), .I3(n24651), .S0(
        n26119), .S1(n26149), .ZN(n24713) );
  MUX41 U8178 ( .I0(n24706), .I1(n24696), .I2(n24701), .I3(n24691), .S0(
        n26120), .S1(n26150), .ZN(n24712) );
  MUX41 U8179 ( .I0(n24541), .I1(n24542), .I2(n24543), .I3(n24544), .S0(
        n26090), .S1(raddr[6]), .ZN(n24540) );
  MUX41 U8180 ( .I0(n24495), .I1(n24485), .I2(n24490), .I3(n24480), .S0(
        n26119), .S1(n26149), .ZN(n24542) );
  MUX41 U8181 ( .I0(n24475), .I1(n24465), .I2(n24470), .I3(n24460), .S0(
        n26119), .S1(n26149), .ZN(n24544) );
  MUX41 U8182 ( .I0(n24535), .I1(n24525), .I2(n24530), .I3(n24520), .S0(
        n26119), .S1(n26149), .ZN(n24541) );
  MUX41 U8183 ( .I0(n25396), .I1(n25397), .I2(n25398), .I3(n25399), .S0(
        raddr[7]), .S1(n26094), .ZN(n25395) );
  MUX41 U8184 ( .I0(n25330), .I1(n25320), .I2(n25325), .I3(n25315), .S0(
        n26122), .S1(n26152), .ZN(n25399) );
  MUX41 U8185 ( .I0(n25350), .I1(n25340), .I2(n25345), .I3(n25335), .S0(
        n26122), .S1(n26152), .ZN(n25397) );
  MUX41 U8186 ( .I0(n25390), .I1(n25380), .I2(n25385), .I3(n25375), .S0(
        n26122), .S1(n26152), .ZN(n25396) );
  MUX41 U8187 ( .I0(n25225), .I1(n25226), .I2(n25227), .I3(n25228), .S0(
        raddr[7]), .S1(n26094), .ZN(n25224) );
  MUX41 U8188 ( .I0(n25179), .I1(n25169), .I2(n25174), .I3(n25164), .S0(
        n26121), .S1(n26151), .ZN(n25226) );
  MUX41 U8189 ( .I0(n25159), .I1(n25149), .I2(n25154), .I3(n25144), .S0(
        n26121), .S1(n26151), .ZN(n25228) );
  MUX41 U8190 ( .I0(n25219), .I1(n25209), .I2(n25214), .I3(n25204), .S0(
        n26121), .S1(n26151), .ZN(n25225) );
  MUX41 U8191 ( .I0(n26080), .I1(n26081), .I2(n26082), .I3(n26083), .S0(
        n26089), .S1(n26094), .ZN(n26079) );
  MUX41 U8192 ( .I0(n26014), .I1(n26004), .I2(n26009), .I3(n25999), .S0(
        n26124), .S1(n26154), .ZN(n26083) );
  MUX41 U8193 ( .I0(n26034), .I1(n26024), .I2(n26029), .I3(n26019), .S0(
        n26124), .S1(n26154), .ZN(n26081) );
  MUX41 U8194 ( .I0(n26074), .I1(n26064), .I2(n26069), .I3(n26059), .S0(
        n26124), .S1(n26154), .ZN(n26080) );
  MUX41 U8195 ( .I0(n25909), .I1(n25910), .I2(n25911), .I3(n25912), .S0(
        raddr[7]), .S1(n26094), .ZN(n25908) );
  MUX41 U8196 ( .I0(n25863), .I1(n25853), .I2(n25858), .I3(n25848), .S0(
        n26124), .S1(n26154), .ZN(n25910) );
  MUX41 U8197 ( .I0(n25843), .I1(n25833), .I2(n25838), .I3(n25828), .S0(
        n26124), .S1(n26154), .ZN(n25912) );
  MUX41 U8198 ( .I0(n25903), .I1(n25893), .I2(n25898), .I3(n25888), .S0(
        n26124), .S1(n26154), .ZN(n25909) );
  MUX41 U8199 ( .I0(n20773), .I1(n20763), .I2(n20768), .I3(n20758), .S0(
        n26105), .S1(n26135), .ZN(n20779) );
  MUX41 U8200 ( .I0(n20759), .I1(n20760), .I2(n20761), .I3(n20762), .S0(
        n26196), .S1(n26314), .ZN(n20758) );
  MUX41 U8201 ( .I0(n20764), .I1(n20765), .I2(n20766), .I3(n20767), .S0(
        n26196), .S1(n26314), .ZN(n20763) );
  MUX41 U8202 ( .I0(n20774), .I1(n20775), .I2(n20776), .I3(n20777), .S0(
        n26196), .S1(n26314), .ZN(n20773) );
  MUX41 U8203 ( .I0(n20688), .I1(n20678), .I2(n20683), .I3(n20673), .S0(
        n26105), .S1(n26135), .ZN(n20694) );
  MUX41 U8204 ( .I0(n20674), .I1(n20675), .I2(n20676), .I3(n20677), .S0(
        n26195), .S1(n26313), .ZN(n20673) );
  MUX41 U8205 ( .I0(n20679), .I1(n20680), .I2(n20681), .I3(n20682), .S0(
        n26195), .S1(n26313), .ZN(n20678) );
  MUX41 U8206 ( .I0(n20689), .I1(n20690), .I2(n20691), .I3(n20692), .S0(
        n26195), .S1(n26313), .ZN(n20688) );
  MUX41 U8207 ( .I0(n21292), .I1(n21293), .I2(n21294), .I3(n21295), .S0(
        n26088), .S1(n26093), .ZN(n21291) );
  MUX41 U8208 ( .I0(n21226), .I1(n21216), .I2(n21221), .I3(n21211), .S0(
        n26107), .S1(n26137), .ZN(n21295) );
  MUX41 U8209 ( .I0(n21246), .I1(n21236), .I2(n21241), .I3(n21231), .S0(
        n26107), .S1(n26137), .ZN(n21293) );
  MUX41 U8210 ( .I0(n21286), .I1(n21276), .I2(n21281), .I3(n21271), .S0(
        n26107), .S1(n26137), .ZN(n21292) );
  MUX41 U8211 ( .I0(n21121), .I1(n21122), .I2(n21123), .I3(n21124), .S0(
        n26088), .S1(n26094), .ZN(n21120) );
  MUX41 U8212 ( .I0(n21075), .I1(n21065), .I2(n21070), .I3(n21060), .S0(
        n26106), .S1(n26136), .ZN(n21122) );
  MUX41 U8213 ( .I0(n21055), .I1(n21045), .I2(n21050), .I3(n21040), .S0(
        n26106), .S1(n26136), .ZN(n21124) );
  MUX41 U8214 ( .I0(n21115), .I1(n21105), .I2(n21110), .I3(n21100), .S0(
        n26107), .S1(n26137), .ZN(n21121) );
  MUX41 U8215 ( .I0(n21457), .I1(n21447), .I2(n21452), .I3(n21442), .S0(
        n26108), .S1(n26138), .ZN(n21463) );
  MUX41 U8216 ( .I0(n21443), .I1(n21444), .I2(n21445), .I3(n21446), .S0(
        n26206), .S1(n26324), .ZN(n21442) );
  MUX41 U8217 ( .I0(n21448), .I1(n21449), .I2(n21450), .I3(n21451), .S0(
        n26206), .S1(n26324), .ZN(n21447) );
  MUX41 U8218 ( .I0(n21458), .I1(n21459), .I2(n21460), .I3(n21461), .S0(
        n26206), .S1(n26324), .ZN(n21457) );
  MUX41 U8219 ( .I0(n21372), .I1(n21362), .I2(n21367), .I3(n21357), .S0(
        n26108), .S1(n26138), .ZN(n21378) );
  MUX41 U8220 ( .I0(n21358), .I1(n21359), .I2(n21360), .I3(n21361), .S0(
        n26205), .S1(n26323), .ZN(n21357) );
  MUX41 U8221 ( .I0(n21363), .I1(n21364), .I2(n21365), .I3(n21366), .S0(
        n26205), .S1(n26323), .ZN(n21362) );
  MUX41 U8222 ( .I0(n21373), .I1(n21374), .I2(n21375), .I3(n21376), .S0(
        n26205), .S1(n26323), .ZN(n21372) );
  MUX41 U8223 ( .I0(n22141), .I1(n22131), .I2(n22136), .I3(n22126), .S0(
        n26110), .S1(n26140), .ZN(n22147) );
  MUX41 U8224 ( .I0(n22127), .I1(n22128), .I2(n22129), .I3(n22130), .S0(
        n26216), .S1(n26334), .ZN(n22126) );
  MUX41 U8225 ( .I0(n22132), .I1(n22133), .I2(n22134), .I3(n22135), .S0(
        n26216), .S1(n26334), .ZN(n22131) );
  MUX41 U8226 ( .I0(n22142), .I1(n22143), .I2(n22144), .I3(n22145), .S0(
        n26216), .S1(n26334), .ZN(n22141) );
  MUX41 U8227 ( .I0(n22056), .I1(n22046), .I2(n22051), .I3(n22041), .S0(
        n26110), .S1(n26140), .ZN(n22062) );
  MUX41 U8228 ( .I0(n22042), .I1(n22043), .I2(n22044), .I3(n22045), .S0(
        n26214), .S1(n26332), .ZN(n22041) );
  MUX41 U8229 ( .I0(n22047), .I1(n22048), .I2(n22049), .I3(n22050), .S0(
        n26214), .S1(n26332), .ZN(n22046) );
  MUX41 U8230 ( .I0(n22057), .I1(n22058), .I2(n22059), .I3(n22060), .S0(
        n26215), .S1(n26333), .ZN(n22056) );
  MUX41 U8231 ( .I0(n22825), .I1(n22815), .I2(n22820), .I3(n22810), .S0(
        n26113), .S1(n26143), .ZN(n22831) );
  MUX41 U8232 ( .I0(n22811), .I1(n22812), .I2(n22813), .I3(n22814), .S0(
        n26225), .S1(n26343), .ZN(n22810) );
  MUX41 U8233 ( .I0(n22816), .I1(n22817), .I2(n22818), .I3(n22819), .S0(
        n26226), .S1(n26344), .ZN(n22815) );
  MUX41 U8234 ( .I0(n22826), .I1(n22827), .I2(n22828), .I3(n22829), .S0(
        n26226), .S1(n26344), .ZN(n22825) );
  MUX41 U8235 ( .I0(n22740), .I1(n22730), .I2(n22735), .I3(n22725), .S0(
        n26112), .S1(n26142), .ZN(n22746) );
  MUX41 U8236 ( .I0(n22726), .I1(n22727), .I2(n22728), .I3(n22729), .S0(
        n26224), .S1(n26342), .ZN(n22725) );
  MUX41 U8237 ( .I0(n22731), .I1(n22732), .I2(n22733), .I3(n22734), .S0(
        n26224), .S1(n26342), .ZN(n22730) );
  MUX41 U8238 ( .I0(n22741), .I1(n22742), .I2(n22743), .I3(n22744), .S0(
        n26224), .S1(n26342), .ZN(n22740) );
  MUX41 U8239 ( .I0(n23509), .I1(n23499), .I2(n23504), .I3(n23494), .S0(
        n26115), .S1(n26145), .ZN(n23515) );
  MUX41 U8240 ( .I0(n23495), .I1(n23496), .I2(n23497), .I3(n23498), .S0(
        n26235), .S1(n26353), .ZN(n23494) );
  MUX41 U8241 ( .I0(n23500), .I1(n23501), .I2(n23502), .I3(n23503), .S0(
        n26235), .S1(n26353), .ZN(n23499) );
  MUX41 U8242 ( .I0(n23510), .I1(n23511), .I2(n23512), .I3(n23513), .S0(
        n26236), .S1(n26354), .ZN(n23509) );
  MUX41 U8243 ( .I0(n23424), .I1(n23414), .I2(n23419), .I3(n23409), .S0(
        n26115), .S1(n26145), .ZN(n23430) );
  MUX41 U8244 ( .I0(n23410), .I1(n23411), .I2(n23412), .I3(n23413), .S0(
        n26234), .S1(n26352), .ZN(n23409) );
  MUX41 U8245 ( .I0(n23415), .I1(n23416), .I2(n23417), .I3(n23418), .S0(
        n26234), .S1(n26352), .ZN(n23414) );
  MUX41 U8246 ( .I0(n23425), .I1(n23426), .I2(n23427), .I3(n23428), .S0(
        n26234), .S1(n26352), .ZN(n23424) );
  MUX41 U8247 ( .I0(n24193), .I1(n24183), .I2(n24188), .I3(n24178), .S0(
        n26118), .S1(n26148), .ZN(n24199) );
  MUX41 U8248 ( .I0(n24179), .I1(n24180), .I2(n24181), .I3(n24182), .S0(
        n26245), .S1(n26363), .ZN(n24178) );
  MUX41 U8249 ( .I0(n24184), .I1(n24185), .I2(n24186), .I3(n24187), .S0(
        n26245), .S1(n26363), .ZN(n24183) );
  MUX41 U8250 ( .I0(n24194), .I1(n24195), .I2(n24196), .I3(n24197), .S0(
        n26245), .S1(n26363), .ZN(n24193) );
  MUX41 U8251 ( .I0(n24108), .I1(n24098), .I2(n24103), .I3(n24093), .S0(
        n26117), .S1(n26147), .ZN(n24114) );
  MUX41 U8252 ( .I0(n24094), .I1(n24095), .I2(n24096), .I3(n24097), .S0(
        n26244), .S1(n26362), .ZN(n24093) );
  MUX41 U8253 ( .I0(n24099), .I1(n24100), .I2(n24101), .I3(n24102), .S0(
        n26244), .S1(n26362), .ZN(n24098) );
  MUX41 U8254 ( .I0(n24109), .I1(n24110), .I2(n24111), .I3(n24112), .S0(
        n26244), .S1(n26362), .ZN(n24108) );
  MUX41 U8255 ( .I0(n24877), .I1(n24867), .I2(n24872), .I3(n24862), .S0(
        n26120), .S1(n26150), .ZN(n24883) );
  MUX41 U8256 ( .I0(n24863), .I1(n24864), .I2(n24865), .I3(n24866), .S0(
        n26255), .S1(n26373), .ZN(n24862) );
  MUX41 U8257 ( .I0(n24868), .I1(n24869), .I2(n24870), .I3(n24871), .S0(
        n26255), .S1(n26373), .ZN(n24867) );
  MUX41 U8258 ( .I0(n24878), .I1(n24879), .I2(n24880), .I3(n24881), .S0(
        n26255), .S1(n26373), .ZN(n24877) );
  MUX41 U8259 ( .I0(n24792), .I1(n24782), .I2(n24787), .I3(n24777), .S0(
        n26120), .S1(n26150), .ZN(n24798) );
  MUX41 U8260 ( .I0(n24778), .I1(n24779), .I2(n24780), .I3(n24781), .S0(
        n26254), .S1(n26372), .ZN(n24777) );
  MUX41 U8261 ( .I0(n24783), .I1(n24784), .I2(n24785), .I3(n24786), .S0(
        n26254), .S1(n26372), .ZN(n24782) );
  MUX41 U8262 ( .I0(n24793), .I1(n24794), .I2(n24795), .I3(n24796), .S0(
        n26254), .S1(n26372), .ZN(n24792) );
  MUX41 U8263 ( .I0(n25561), .I1(n25551), .I2(n25556), .I3(n25546), .S0(
        n26123), .S1(n26153), .ZN(n25567) );
  MUX41 U8264 ( .I0(n25547), .I1(n25548), .I2(n25549), .I3(n25550), .S0(
        n26265), .S1(n26383), .ZN(n25546) );
  MUX41 U8265 ( .I0(n25552), .I1(n25553), .I2(n25554), .I3(n25555), .S0(
        n26265), .S1(n26383), .ZN(n25551) );
  MUX41 U8266 ( .I0(n25562), .I1(n25563), .I2(n25564), .I3(n25565), .S0(
        n26265), .S1(n26383), .ZN(n25561) );
  MUX41 U8267 ( .I0(n25476), .I1(n25466), .I2(n25471), .I3(n25461), .S0(
        n26122), .S1(n26152), .ZN(n25482) );
  MUX41 U8268 ( .I0(n25462), .I1(n25463), .I2(n25464), .I3(n25465), .S0(
        n26264), .S1(n26382), .ZN(n25461) );
  MUX41 U8269 ( .I0(n25467), .I1(n25468), .I2(n25469), .I3(n25470), .S0(
        n26264), .S1(n26382), .ZN(n25466) );
  MUX41 U8270 ( .I0(n25477), .I1(n25478), .I2(n25479), .I3(n25480), .S0(
        n26264), .S1(n26382), .ZN(n25476) );
  BUF U8271 ( .I(raddr[0]), .Z(n27340) );
  BUF U8272 ( .I(raddr[1]), .Z(n26865) );
  BUF U8273 ( .I(n27339), .Z(n26866) );
  BUF U8274 ( .I(raddr[0]), .Z(n27339) );
  BUF U8275 ( .I(n26864), .Z(n26391) );
  BUF U8276 ( .I(raddr[1]), .Z(n26864) );
  BUF U8277 ( .I(n29318), .Z(n26157) );
  BUF U8278 ( .I(n29317), .Z(n26275) );
  BUF U8279 ( .I(n29318), .Z(n26156) );
  BUF U8280 ( .I(n29317), .Z(n26274) );
  BUF U8281 ( .I(n29318), .Z(n26155) );
  BUF U8282 ( .I(n29317), .Z(n26273) );
  NOR3 U8283 ( .A1(waddr[3]), .A2(waddr[4]), .A3(n29587), .ZN(n4158) );
  NOR3 U8284 ( .A1(waddr[3]), .A2(waddr[5]), .A3(n29586), .ZN(n4192) );
  NOR3 U8285 ( .A1(waddr[4]), .A2(waddr[5]), .A3(n29585), .ZN(n4209) );
  NOR3 U8286 ( .A1(n29586), .A2(waddr[3]), .A3(n29587), .ZN(n4124) );
  NOR3 U8287 ( .A1(n29585), .A2(waddr[4]), .A3(n29587), .ZN(n4141) );
  NOR3 U8288 ( .A1(n29585), .A2(waddr[5]), .A3(n29586), .ZN(n4175) );
  NOR3 U8289 ( .A1(waddr[6]), .A2(waddr[7]), .A3(n29590), .ZN(n605) );
  NOR3 U8290 ( .A1(waddr[6]), .A2(waddr[8]), .A3(n29589), .ZN(n865) );
  NOR3 U8291 ( .A1(waddr[7]), .A2(waddr[8]), .A3(n29588), .ZN(n995) );
  NOR3 U8292 ( .A1(n29589), .A2(waddr[6]), .A3(n29590), .ZN(n345) );
  NOR3 U8293 ( .A1(n29588), .A2(waddr[7]), .A3(n29590), .ZN(n475) );
  NOR3 U8294 ( .A1(n29588), .A2(waddr[8]), .A3(n29589), .ZN(n735) );
  BUF U8295 ( .I(n26085), .Z(n26087) );
  BUF U8296 ( .I(n26085), .Z(n26086) );
  BUF U8297 ( .I(n26091), .Z(n26092) );
  INV U8298 ( .I(n26092), .ZN(n26094) );
  BUF U8299 ( .I(n26125), .Z(n26134) );
  BUF U8300 ( .I(n29319), .Z(n26125) );
  BUF U8301 ( .I(n29320), .Z(n26096) );
  BUF U8302 ( .I(n29319), .Z(n26126) );
  BUF U8303 ( .I(n29320), .Z(n26097) );
  BUF U8304 ( .I(n29319), .Z(n26127) );
  BUF U8305 ( .I(n26095), .Z(n26104) );
  BUF U8306 ( .I(n29320), .Z(n26095) );
  NOR3 U8307 ( .A1(waddr[4]), .A2(waddr[5]), .A3(waddr[3]), .ZN(n4226) );
  NOR3 U8308 ( .A1(waddr[7]), .A2(waddr[8]), .A3(waddr[6]), .ZN(n1125) );
  NOR2 U8309 ( .A1(waddr[10]), .A2(waddr[9]), .ZN(n3321) );
  NOR2 U8310 ( .A1(n29592), .A2(waddr[9]), .ZN(n1255) );
  NOR2 U8311 ( .A1(n29591), .A2(waddr[10]), .ZN(n2288) );
  BUF U8312 ( .I(n17), .Z(n28612) );
  BUF U8313 ( .I(n20), .Z(n27907) );
  BUF U8314 ( .I(n21), .Z(n27672) );
  BUF U8315 ( .I(n17), .Z(n28613) );
  BUF U8316 ( .I(n20), .Z(n27908) );
  BUF U8317 ( .I(n21), .Z(n27673) );
  BUF U8318 ( .I(n17), .Z(n28614) );
  BUF U8319 ( .I(n20), .Z(n27909) );
  BUF U8320 ( .I(n21), .Z(n27674) );
  BUF U8321 ( .I(n17), .Z(n28615) );
  BUF U8322 ( .I(n20), .Z(n27910) );
  BUF U8323 ( .I(n21), .Z(n27675) );
  BUF U8324 ( .I(n17), .Z(n28616) );
  BUF U8325 ( .I(n20), .Z(n27911) );
  BUF U8326 ( .I(n21), .Z(n27676) );
  BUF U8327 ( .I(n17), .Z(n28617) );
  BUF U8328 ( .I(n20), .Z(n27912) );
  BUF U8329 ( .I(n21), .Z(n27677) );
  BUF U8330 ( .I(n14), .Z(n29082) );
  BUF U8331 ( .I(n16), .Z(n28847) );
  BUF U8332 ( .I(n18), .Z(n28377) );
  BUF U8333 ( .I(n19), .Z(n28142) );
  BUF U8334 ( .I(n22), .Z(n27437) );
  BUF U8335 ( .I(n14), .Z(n29083) );
  BUF U8336 ( .I(n16), .Z(n28848) );
  BUF U8337 ( .I(n18), .Z(n28378) );
  BUF U8338 ( .I(n19), .Z(n28143) );
  BUF U8339 ( .I(n22), .Z(n27438) );
  BUF U8340 ( .I(n14), .Z(n29084) );
  BUF U8341 ( .I(n16), .Z(n28849) );
  BUF U8342 ( .I(n18), .Z(n28379) );
  BUF U8343 ( .I(n19), .Z(n28144) );
  BUF U8344 ( .I(n22), .Z(n27439) );
  BUF U8345 ( .I(n14), .Z(n29085) );
  BUF U8346 ( .I(n16), .Z(n28850) );
  BUF U8347 ( .I(n18), .Z(n28380) );
  BUF U8348 ( .I(n19), .Z(n28145) );
  BUF U8349 ( .I(n22), .Z(n27440) );
  BUF U8350 ( .I(n14), .Z(n29086) );
  BUF U8351 ( .I(n16), .Z(n28851) );
  BUF U8352 ( .I(n18), .Z(n28381) );
  BUF U8353 ( .I(n19), .Z(n28146) );
  BUF U8354 ( .I(n22), .Z(n27441) );
  BUF U8355 ( .I(n14), .Z(n29087) );
  BUF U8356 ( .I(n16), .Z(n28852) );
  BUF U8357 ( .I(n18), .Z(n28382) );
  BUF U8358 ( .I(n19), .Z(n28147) );
  BUF U8359 ( .I(n22), .Z(n27442) );
  MUX41 U8360 ( .I0(ram[3480]), .I1(ram[3472]), .I2(ram[3464]), .I3(
        ram[3456]), .S0(n27032), .S1(n26557), .ZN(n20757) );
  MUX41 U8361 ( .I0(ram[3224]), .I1(ram[3216]), .I2(ram[3208]), .I3(
        ram[3200]), .S0(n27031), .S1(n26556), .ZN(n20747) );
  MUX41 U8362 ( .I0(ram[3096]), .I1(ram[3088]), .I2(ram[3080]), .I3(
        ram[3072]), .S0(n27031), .S1(n26556), .ZN(n20742) );
  MUX41 U8363 ( .I0(ram[3992]), .I1(ram[3984]), .I2(ram[3976]), .I3(
        ram[3968]), .S0(n27033), .S1(n26558), .ZN(n20777) );
  MUX41 U8364 ( .I0(ram[1432]), .I1(ram[1424]), .I2(ram[1416]), .I3(
        ram[1408]), .S0(n27027), .S1(n26552), .ZN(n20672) );
  MUX41 U8365 ( .I0(ram[1176]), .I1(ram[1168]), .I2(ram[1160]), .I3(
        ram[1152]), .S0(n27026), .S1(n26551), .ZN(n20662) );
  MUX41 U8366 ( .I0(ram[1048]), .I1(ram[1040]), .I2(ram[1032]), .I3(
        ram[1024]), .S0(n27026), .S1(n26551), .ZN(n20657) );
  MUX41 U8367 ( .I0(ram[1944]), .I1(ram[1936]), .I2(ram[1928]), .I3(
        ram[1920]), .S0(n27028), .S1(n26553), .ZN(n20692) );
  MUX41 U8368 ( .I0(ram[3481]), .I1(ram[3473]), .I2(ram[3465]), .I3(
        ram[3457]), .S0(n27071), .S1(n26596), .ZN(n21441) );
  MUX41 U8369 ( .I0(ram[3225]), .I1(ram[3217]), .I2(ram[3209]), .I3(
        ram[3201]), .S0(n27071), .S1(n26596), .ZN(n21431) );
  MUX41 U8370 ( .I0(ram[3097]), .I1(ram[3089]), .I2(ram[3081]), .I3(
        ram[3073]), .S0(n27070), .S1(n26595), .ZN(n21426) );
  MUX41 U8371 ( .I0(ram[3993]), .I1(ram[3985]), .I2(ram[3977]), .I3(
        ram[3969]), .S0(n27072), .S1(n26597), .ZN(n21461) );
  MUX41 U8372 ( .I0(ram[1433]), .I1(ram[1425]), .I2(ram[1417]), .I3(
        ram[1409]), .S0(n27066), .S1(n26591), .ZN(n21356) );
  MUX41 U8373 ( .I0(ram[1177]), .I1(ram[1169]), .I2(ram[1161]), .I3(
        ram[1153]), .S0(n27066), .S1(n26591), .ZN(n21346) );
  MUX41 U8374 ( .I0(ram[1049]), .I1(ram[1041]), .I2(ram[1033]), .I3(
        ram[1025]), .S0(n27065), .S1(n26590), .ZN(n21341) );
  MUX41 U8375 ( .I0(ram[1945]), .I1(ram[1937]), .I2(ram[1929]), .I3(
        ram[1921]), .S0(n27067), .S1(n26592), .ZN(n21376) );
  MUX41 U8376 ( .I0(ram[3482]), .I1(ram[3474]), .I2(ram[3466]), .I3(
        ram[3458]), .S0(n27111), .S1(n26636), .ZN(n22125) );
  MUX41 U8377 ( .I0(ram[3226]), .I1(ram[3218]), .I2(ram[3210]), .I3(
        ram[3202]), .S0(n27110), .S1(n26635), .ZN(n22115) );
  MUX41 U8378 ( .I0(ram[3098]), .I1(ram[3090]), .I2(ram[3082]), .I3(
        ram[3074]), .S0(n27110), .S1(n26635), .ZN(n22110) );
  MUX41 U8379 ( .I0(ram[3994]), .I1(ram[3986]), .I2(ram[3978]), .I3(
        ram[3970]), .S0(n27112), .S1(n26637), .ZN(n22145) );
  MUX41 U8380 ( .I0(ram[1434]), .I1(ram[1426]), .I2(ram[1418]), .I3(
        ram[1410]), .S0(n27106), .S1(n26631), .ZN(n22040) );
  MUX41 U8381 ( .I0(ram[1178]), .I1(ram[1170]), .I2(ram[1162]), .I3(
        ram[1154]), .S0(n27105), .S1(n26630), .ZN(n22030) );
  MUX41 U8382 ( .I0(ram[1050]), .I1(ram[1042]), .I2(ram[1034]), .I3(
        ram[1026]), .S0(n27105), .S1(n26630), .ZN(n22025) );
  MUX41 U8383 ( .I0(ram[1946]), .I1(ram[1938]), .I2(ram[1930]), .I3(
        ram[1922]), .S0(n27107), .S1(n26632), .ZN(n22060) );
  MUX41 U8384 ( .I0(ram[3483]), .I1(ram[3475]), .I2(ram[3467]), .I3(
        ram[3459]), .S0(n27150), .S1(n26675), .ZN(n22809) );
  MUX41 U8385 ( .I0(ram[3227]), .I1(ram[3219]), .I2(ram[3211]), .I3(
        ram[3203]), .S0(n27149), .S1(n26674), .ZN(n22799) );
  MUX41 U8386 ( .I0(ram[3099]), .I1(ram[3091]), .I2(ram[3083]), .I3(
        ram[3075]), .S0(n27149), .S1(n26674), .ZN(n22794) );
  MUX41 U8387 ( .I0(ram[3995]), .I1(ram[3987]), .I2(ram[3979]), .I3(
        ram[3971]), .S0(n27151), .S1(n26676), .ZN(n22829) );
  MUX41 U8388 ( .I0(ram[1435]), .I1(ram[1427]), .I2(ram[1419]), .I3(
        ram[1411]), .S0(n27145), .S1(n26670), .ZN(n22724) );
  MUX41 U8389 ( .I0(ram[1179]), .I1(ram[1171]), .I2(ram[1163]), .I3(
        ram[1155]), .S0(n27144), .S1(n26669), .ZN(n22714) );
  MUX41 U8390 ( .I0(ram[1051]), .I1(ram[1043]), .I2(ram[1035]), .I3(
        ram[1027]), .S0(n27144), .S1(n26669), .ZN(n22709) );
  MUX41 U8391 ( .I0(ram[1947]), .I1(ram[1939]), .I2(ram[1931]), .I3(
        ram[1923]), .S0(n27146), .S1(n26671), .ZN(n22744) );
  MUX41 U8392 ( .I0(ram[3484]), .I1(ram[3476]), .I2(ram[3468]), .I3(
        ram[3460]), .S0(n27189), .S1(n26714), .ZN(n23493) );
  MUX41 U8393 ( .I0(ram[3228]), .I1(ram[3220]), .I2(ram[3212]), .I3(
        ram[3204]), .S0(n27189), .S1(n26714), .ZN(n23483) );
  MUX41 U8394 ( .I0(ram[3100]), .I1(ram[3092]), .I2(ram[3084]), .I3(
        ram[3076]), .S0(n27188), .S1(n26713), .ZN(n23478) );
  MUX41 U8395 ( .I0(ram[3996]), .I1(ram[3988]), .I2(ram[3980]), .I3(
        ram[3972]), .S0(n27191), .S1(n26716), .ZN(n23513) );
  MUX41 U8396 ( .I0(ram[1436]), .I1(ram[1428]), .I2(ram[1420]), .I3(
        ram[1412]), .S0(n27184), .S1(n26709), .ZN(n23408) );
  MUX41 U8397 ( .I0(ram[1180]), .I1(ram[1172]), .I2(ram[1164]), .I3(
        ram[1156]), .S0(n27184), .S1(n26709), .ZN(n23398) );
  MUX41 U8398 ( .I0(ram[1052]), .I1(ram[1044]), .I2(ram[1036]), .I3(
        ram[1028]), .S0(n27183), .S1(n26708), .ZN(n23393) );
  MUX41 U8399 ( .I0(ram[1948]), .I1(ram[1940]), .I2(ram[1932]), .I3(
        ram[1924]), .S0(n27186), .S1(n26711), .ZN(n23428) );
  MUX41 U8400 ( .I0(ram[3485]), .I1(ram[3477]), .I2(ram[3469]), .I3(
        ram[3461]), .S0(n27229), .S1(n26754), .ZN(n24177) );
  MUX41 U8401 ( .I0(ram[3229]), .I1(ram[3221]), .I2(ram[3213]), .I3(
        ram[3205]), .S0(n27228), .S1(n26753), .ZN(n24167) );
  MUX41 U8402 ( .I0(ram[3101]), .I1(ram[3093]), .I2(ram[3085]), .I3(
        ram[3077]), .S0(n27228), .S1(n26753), .ZN(n24162) );
  MUX41 U8403 ( .I0(ram[3997]), .I1(ram[3989]), .I2(ram[3981]), .I3(
        ram[3973]), .S0(n27230), .S1(n26755), .ZN(n24197) );
  MUX41 U8404 ( .I0(ram[1437]), .I1(ram[1429]), .I2(ram[1421]), .I3(
        ram[1413]), .S0(n27224), .S1(n26749), .ZN(n24092) );
  MUX41 U8405 ( .I0(ram[1181]), .I1(ram[1173]), .I2(ram[1165]), .I3(
        ram[1157]), .S0(n27223), .S1(n26748), .ZN(n24082) );
  MUX41 U8406 ( .I0(ram[1053]), .I1(ram[1045]), .I2(ram[1037]), .I3(
        ram[1029]), .S0(n27223), .S1(n26748), .ZN(n24077) );
  MUX41 U8407 ( .I0(ram[1949]), .I1(ram[1941]), .I2(ram[1933]), .I3(
        ram[1925]), .S0(n27225), .S1(n26750), .ZN(n24112) );
  MUX41 U8408 ( .I0(ram[3486]), .I1(ram[3478]), .I2(ram[3470]), .I3(
        ram[3462]), .S0(n27268), .S1(n26793), .ZN(n24861) );
  MUX41 U8409 ( .I0(ram[3230]), .I1(ram[3222]), .I2(ram[3214]), .I3(
        ram[3206]), .S0(n27267), .S1(n26792), .ZN(n24851) );
  MUX41 U8410 ( .I0(ram[3102]), .I1(ram[3094]), .I2(ram[3086]), .I3(
        ram[3078]), .S0(n27267), .S1(n26792), .ZN(n24846) );
  MUX41 U8411 ( .I0(ram[3998]), .I1(ram[3990]), .I2(ram[3982]), .I3(
        ram[3974]), .S0(n27269), .S1(n26794), .ZN(n24881) );
  MUX41 U8412 ( .I0(ram[1438]), .I1(ram[1430]), .I2(ram[1422]), .I3(
        ram[1414]), .S0(n27263), .S1(n26788), .ZN(n24776) );
  MUX41 U8413 ( .I0(ram[1182]), .I1(ram[1174]), .I2(ram[1166]), .I3(
        ram[1158]), .S0(n27263), .S1(n26788), .ZN(n24766) );
  MUX41 U8414 ( .I0(ram[1054]), .I1(ram[1046]), .I2(ram[1038]), .I3(
        ram[1030]), .S0(n27262), .S1(n26787), .ZN(n24761) );
  MUX41 U8415 ( .I0(ram[1950]), .I1(ram[1942]), .I2(ram[1934]), .I3(
        ram[1926]), .S0(n27264), .S1(n26789), .ZN(n24796) );
  MUX41 U8416 ( .I0(ram[3487]), .I1(ram[3479]), .I2(ram[3471]), .I3(
        ram[3463]), .S0(n27307), .S1(n26832), .ZN(n25545) );
  MUX41 U8417 ( .I0(ram[3231]), .I1(ram[3223]), .I2(ram[3215]), .I3(
        ram[3207]), .S0(n27307), .S1(n26832), .ZN(n25535) );
  MUX41 U8418 ( .I0(ram[3103]), .I1(ram[3095]), .I2(ram[3087]), .I3(
        ram[3079]), .S0(n27307), .S1(n26832), .ZN(n25530) );
  MUX41 U8419 ( .I0(ram[3999]), .I1(ram[3991]), .I2(ram[3983]), .I3(
        ram[3975]), .S0(n27309), .S1(n26834), .ZN(n25565) );
  MUX41 U8420 ( .I0(ram[1439]), .I1(ram[1431]), .I2(ram[1423]), .I3(
        ram[1415]), .S0(n27303), .S1(n26828), .ZN(n25460) );
  MUX41 U8421 ( .I0(ram[1183]), .I1(ram[1175]), .I2(ram[1167]), .I3(
        ram[1159]), .S0(n27302), .S1(n26827), .ZN(n25450) );
  MUX41 U8422 ( .I0(ram[1055]), .I1(ram[1047]), .I2(ram[1039]), .I3(
        ram[1031]), .S0(n27302), .S1(n26827), .ZN(n25445) );
  MUX41 U8423 ( .I0(ram[1951]), .I1(ram[1943]), .I2(ram[1935]), .I3(
        ram[1927]), .S0(n27304), .S1(n26829), .ZN(n25480) );
  MUX41 U8424 ( .I0(ram[15768]), .I1(ram[15760]), .I2(ram[15752]), .I3(
        ram[15744]), .S0(n27061), .S1(n26586), .ZN(n21270) );
  MUX41 U8425 ( .I0(ram[15512]), .I1(ram[15504]), .I2(ram[15496]), .I3(
        ram[15488]), .S0(n27061), .S1(n26586), .ZN(n21260) );
  MUX41 U8426 ( .I0(ram[15384]), .I1(ram[15376]), .I2(ram[15368]), .I3(
        ram[15360]), .S0(n27060), .S1(n26585), .ZN(n21255) );
  MUX41 U8427 ( .I0(ram[13720]), .I1(ram[13712]), .I2(ram[13704]), .I3(
        ram[13696]), .S0(n27056), .S1(n26581), .ZN(n21185) );
  MUX41 U8428 ( .I0(ram[13464]), .I1(ram[13456]), .I2(ram[13448]), .I3(
        ram[13440]), .S0(n27056), .S1(n26581), .ZN(n21175) );
  MUX41 U8429 ( .I0(ram[13336]), .I1(ram[13328]), .I2(ram[13320]), .I3(
        ram[13312]), .S0(n27055), .S1(n26580), .ZN(n21170) );
  MUX41 U8430 ( .I0(ram[7576]), .I1(ram[7568]), .I2(ram[7560]), .I3(
        ram[7552]), .S0(n27042), .S1(n26567), .ZN(n20928) );
  MUX41 U8431 ( .I0(ram[7320]), .I1(ram[7312]), .I2(ram[7304]), .I3(
        ram[7296]), .S0(n27041), .S1(n26566), .ZN(n20918) );
  MUX41 U8432 ( .I0(ram[7192]), .I1(ram[7184]), .I2(ram[7176]), .I3(
        ram[7168]), .S0(n27041), .S1(n26566), .ZN(n20913) );
  MUX41 U8433 ( .I0(ram[5528]), .I1(ram[5520]), .I2(ram[5512]), .I3(
        ram[5504]), .S0(n27037), .S1(n26562), .ZN(n20843) );
  MUX41 U8434 ( .I0(ram[11672]), .I1(ram[11664]), .I2(ram[11656]), .I3(
        ram[11648]), .S0(n27051), .S1(n26576), .ZN(n21099) );
  MUX41 U8435 ( .I0(ram[11416]), .I1(ram[11408]), .I2(ram[11400]), .I3(
        ram[11392]), .S0(n27051), .S1(n26576), .ZN(n21089) );
  MUX41 U8436 ( .I0(ram[11288]), .I1(ram[11280]), .I2(ram[11272]), .I3(
        ram[11264]), .S0(n27051), .S1(n26576), .ZN(n21084) );
  MUX41 U8437 ( .I0(ram[9624]), .I1(ram[9616]), .I2(ram[9608]), .I3(
        ram[9600]), .S0(n27047), .S1(n26572), .ZN(n21014) );
  MUX41 U8438 ( .I0(ram[9368]), .I1(ram[9360]), .I2(ram[9352]), .I3(
        ram[9344]), .S0(n27046), .S1(n26571), .ZN(n21004) );
  MUX41 U8439 ( .I0(ram[15769]), .I1(ram[15761]), .I2(ram[15753]), .I3(
        ram[15745]), .S0(n27101), .S1(n26626), .ZN(n21954) );
  MUX41 U8440 ( .I0(ram[15513]), .I1(ram[15505]), .I2(ram[15497]), .I3(
        ram[15489]), .S0(n27100), .S1(n26625), .ZN(n21944) );
  MUX41 U8441 ( .I0(ram[15385]), .I1(ram[15377]), .I2(ram[15369]), .I3(
        ram[15361]), .S0(n27100), .S1(n26625), .ZN(n21939) );
  MUX41 U8442 ( .I0(ram[13721]), .I1(ram[13713]), .I2(ram[13705]), .I3(
        ram[13697]), .S0(n27096), .S1(n26621), .ZN(n21869) );
  MUX41 U8443 ( .I0(ram[13465]), .I1(ram[13457]), .I2(ram[13449]), .I3(
        ram[13441]), .S0(n27095), .S1(n26620), .ZN(n21859) );
  MUX41 U8444 ( .I0(ram[13337]), .I1(ram[13329]), .I2(ram[13321]), .I3(
        ram[13313]), .S0(n27095), .S1(n26620), .ZN(n21854) );
  MUX41 U8445 ( .I0(ram[7577]), .I1(ram[7569]), .I2(ram[7561]), .I3(
        ram[7553]), .S0(n27081), .S1(n26606), .ZN(n21612) );
  MUX41 U8446 ( .I0(ram[7321]), .I1(ram[7313]), .I2(ram[7305]), .I3(
        ram[7297]), .S0(n27080), .S1(n26605), .ZN(n21602) );
  MUX41 U8447 ( .I0(ram[7193]), .I1(ram[7185]), .I2(ram[7177]), .I3(
        ram[7169]), .S0(n27080), .S1(n26605), .ZN(n21597) );
  MUX41 U8448 ( .I0(ram[5529]), .I1(ram[5521]), .I2(ram[5513]), .I3(
        ram[5505]), .S0(n27076), .S1(n26601), .ZN(n21527) );
  MUX41 U8449 ( .I0(ram[11673]), .I1(ram[11665]), .I2(ram[11657]), .I3(
        ram[11649]), .S0(n27091), .S1(n26616), .ZN(n21783) );
  MUX41 U8450 ( .I0(ram[11417]), .I1(ram[11409]), .I2(ram[11401]), .I3(
        ram[11393]), .S0(n27090), .S1(n26615), .ZN(n21773) );
  MUX41 U8451 ( .I0(ram[11289]), .I1(ram[11281]), .I2(ram[11273]), .I3(
        ram[11265]), .S0(n27090), .S1(n26615), .ZN(n21768) );
  MUX41 U8452 ( .I0(ram[9625]), .I1(ram[9617]), .I2(ram[9609]), .I3(
        ram[9601]), .S0(n27086), .S1(n26611), .ZN(n21698) );
  MUX41 U8453 ( .I0(ram[9369]), .I1(ram[9361]), .I2(ram[9353]), .I3(
        ram[9345]), .S0(n27085), .S1(n26610), .ZN(n21688) );
  MUX41 U8454 ( .I0(ram[15770]), .I1(ram[15762]), .I2(ram[15754]), .I3(
        ram[15746]), .S0(n27140), .S1(n26665), .ZN(n22638) );
  MUX41 U8455 ( .I0(ram[15514]), .I1(ram[15506]), .I2(ram[15498]), .I3(
        ram[15490]), .S0(n27139), .S1(n26664), .ZN(n22628) );
  MUX41 U8456 ( .I0(ram[15386]), .I1(ram[15378]), .I2(ram[15370]), .I3(
        ram[15362]), .S0(n27139), .S1(n26664), .ZN(n22623) );
  MUX41 U8457 ( .I0(ram[13722]), .I1(ram[13714]), .I2(ram[13706]), .I3(
        ram[13698]), .S0(n27135), .S1(n26660), .ZN(n22553) );
  MUX41 U8458 ( .I0(ram[13466]), .I1(ram[13458]), .I2(ram[13450]), .I3(
        ram[13442]), .S0(n27135), .S1(n26660), .ZN(n22543) );
  MUX41 U8459 ( .I0(ram[13338]), .I1(ram[13330]), .I2(ram[13322]), .I3(
        ram[13314]), .S0(n27134), .S1(n26659), .ZN(n22538) );
  MUX41 U8460 ( .I0(n22002), .I1(n22003), .I2(n22004), .I3(n22005), .S0(
        n26214), .S1(n26332), .ZN(n22001) );
  MUX41 U8461 ( .I0(ram[538]), .I1(ram[530]), .I2(ram[522]), .I3(ram[514]), .S0(n27103), .S1(n26628), .ZN(n22005) );
  MUX41 U8462 ( .I0(ram[570]), .I1(ram[562]), .I2(ram[554]), .I3(ram[546]), .S0(n27104), .S1(n26629), .ZN(n22003) );
  MUX41 U8463 ( .I0(ram[634]), .I1(ram[626]), .I2(ram[618]), .I3(ram[610]), .S0(n27104), .S1(n26629), .ZN(n22002) );
  MUX41 U8464 ( .I0(ram[7578]), .I1(ram[7570]), .I2(ram[7562]), .I3(
        ram[7554]), .S0(n27120), .S1(n26645), .ZN(n22296) );
  MUX41 U8465 ( .I0(ram[7322]), .I1(ram[7314]), .I2(ram[7306]), .I3(
        ram[7298]), .S0(n27120), .S1(n26645), .ZN(n22286) );
  MUX41 U8466 ( .I0(ram[7194]), .I1(ram[7186]), .I2(ram[7178]), .I3(
        ram[7170]), .S0(n27119), .S1(n26644), .ZN(n22281) );
  MUX41 U8467 ( .I0(ram[5530]), .I1(ram[5522]), .I2(ram[5514]), .I3(
        ram[5506]), .S0(n27115), .S1(n26640), .ZN(n22211) );
  MUX41 U8468 ( .I0(ram[11674]), .I1(ram[11666]), .I2(ram[11658]), .I3(
        ram[11650]), .S0(n27130), .S1(n26655), .ZN(n22467) );
  MUX41 U8469 ( .I0(ram[11418]), .I1(ram[11410]), .I2(ram[11402]), .I3(
        ram[11394]), .S0(n27130), .S1(n26655), .ZN(n22457) );
  MUX41 U8470 ( .I0(ram[11290]), .I1(ram[11282]), .I2(ram[11274]), .I3(
        ram[11266]), .S0(n27129), .S1(n26654), .ZN(n22452) );
  MUX41 U8471 ( .I0(ram[9626]), .I1(ram[9618]), .I2(ram[9610]), .I3(
        ram[9602]), .S0(n27125), .S1(n26650), .ZN(n22382) );
  MUX41 U8472 ( .I0(ram[9370]), .I1(ram[9362]), .I2(ram[9354]), .I3(
        ram[9346]), .S0(n27125), .S1(n26650), .ZN(n22372) );
  MUX41 U8473 ( .I0(ram[9242]), .I1(ram[9234]), .I2(ram[9226]), .I3(
        ram[9218]), .S0(n27124), .S1(n26649), .ZN(n22367) );
  MUX41 U8474 ( .I0(ram[15771]), .I1(ram[15763]), .I2(ram[15755]), .I3(
        ram[15747]), .S0(n27179), .S1(n26704), .ZN(n23322) );
  MUX41 U8475 ( .I0(ram[15515]), .I1(ram[15507]), .I2(ram[15499]), .I3(
        ram[15491]), .S0(n27179), .S1(n26704), .ZN(n23312) );
  MUX41 U8476 ( .I0(ram[15387]), .I1(ram[15379]), .I2(ram[15371]), .I3(
        ram[15363]), .S0(n27179), .S1(n26704), .ZN(n23307) );
  MUX41 U8477 ( .I0(ram[13723]), .I1(ram[13715]), .I2(ram[13707]), .I3(
        ram[13699]), .S0(n27175), .S1(n26700), .ZN(n23237) );
  MUX41 U8478 ( .I0(ram[13467]), .I1(ram[13459]), .I2(ram[13451]), .I3(
        ram[13443]), .S0(n27174), .S1(n26699), .ZN(n23227) );
  MUX41 U8479 ( .I0(ram[13339]), .I1(ram[13331]), .I2(ram[13323]), .I3(
        ram[13315]), .S0(n27174), .S1(n26699), .ZN(n23222) );
  MUX41 U8480 ( .I0(n22686), .I1(n22687), .I2(n22688), .I3(n22689), .S0(
        n26224), .S1(n26342), .ZN(n22685) );
  MUX41 U8481 ( .I0(ram[539]), .I1(ram[531]), .I2(ram[523]), .I3(ram[515]), .S0(n27143), .S1(n26668), .ZN(n22689) );
  MUX41 U8482 ( .I0(ram[571]), .I1(ram[563]), .I2(ram[555]), .I3(ram[547]), .S0(n27143), .S1(n26668), .ZN(n22687) );
  MUX41 U8483 ( .I0(ram[635]), .I1(ram[627]), .I2(ram[619]), .I3(ram[611]), .S0(n27143), .S1(n26668), .ZN(n22686) );
  MUX41 U8484 ( .I0(ram[7579]), .I1(ram[7571]), .I2(ram[7563]), .I3(
        ram[7555]), .S0(n27160), .S1(n26685), .ZN(n22980) );
  MUX41 U8485 ( .I0(ram[7323]), .I1(ram[7315]), .I2(ram[7307]), .I3(
        ram[7299]), .S0(n27159), .S1(n26684), .ZN(n22970) );
  MUX41 U8486 ( .I0(ram[7195]), .I1(ram[7187]), .I2(ram[7179]), .I3(
        ram[7171]), .S0(n27159), .S1(n26684), .ZN(n22965) );
  MUX41 U8487 ( .I0(ram[5531]), .I1(ram[5523]), .I2(ram[5515]), .I3(
        ram[5507]), .S0(n27155), .S1(n26680), .ZN(n22895) );
  MUX41 U8488 ( .I0(ram[11675]), .I1(ram[11667]), .I2(ram[11659]), .I3(
        ram[11651]), .S0(n27170), .S1(n26695), .ZN(n23151) );
  MUX41 U8489 ( .I0(ram[11419]), .I1(ram[11411]), .I2(ram[11403]), .I3(
        ram[11395]), .S0(n27169), .S1(n26694), .ZN(n23141) );
  MUX41 U8490 ( .I0(ram[11291]), .I1(ram[11283]), .I2(ram[11275]), .I3(
        ram[11267]), .S0(n27169), .S1(n26694), .ZN(n23136) );
  MUX41 U8491 ( .I0(ram[9627]), .I1(ram[9619]), .I2(ram[9611]), .I3(
        ram[9603]), .S0(n27165), .S1(n26690), .ZN(n23066) );
  MUX41 U8492 ( .I0(ram[9371]), .I1(ram[9363]), .I2(ram[9355]), .I3(
        ram[9347]), .S0(n27164), .S1(n26689), .ZN(n23056) );
  MUX41 U8493 ( .I0(ram[9243]), .I1(ram[9235]), .I2(ram[9227]), .I3(
        ram[9219]), .S0(n27164), .S1(n26689), .ZN(n23051) );
  MUX41 U8494 ( .I0(ram[15772]), .I1(ram[15764]), .I2(ram[15756]), .I3(
        ram[15748]), .S0(n27219), .S1(n26744), .ZN(n24006) );
  MUX41 U8495 ( .I0(ram[15516]), .I1(ram[15508]), .I2(ram[15500]), .I3(
        ram[15492]), .S0(n27218), .S1(n26743), .ZN(n23996) );
  MUX41 U8496 ( .I0(ram[15388]), .I1(ram[15380]), .I2(ram[15372]), .I3(
        ram[15364]), .S0(n27218), .S1(n26743), .ZN(n23991) );
  MUX41 U8497 ( .I0(ram[13724]), .I1(ram[13716]), .I2(ram[13708]), .I3(
        ram[13700]), .S0(n27214), .S1(n26739), .ZN(n23921) );
  MUX41 U8498 ( .I0(ram[13468]), .I1(ram[13460]), .I2(ram[13452]), .I3(
        ram[13444]), .S0(n27213), .S1(n26738), .ZN(n23911) );
  MUX41 U8499 ( .I0(ram[13340]), .I1(ram[13332]), .I2(ram[13324]), .I3(
        ram[13316]), .S0(n27213), .S1(n26738), .ZN(n23906) );
  MUX41 U8500 ( .I0(n23370), .I1(n23371), .I2(n23372), .I3(n23373), .S0(
        n26233), .S1(n26351), .ZN(n23369) );
  MUX41 U8501 ( .I0(ram[540]), .I1(ram[532]), .I2(ram[524]), .I3(ram[516]), .S0(n27182), .S1(n26707), .ZN(n23373) );
  MUX41 U8502 ( .I0(ram[572]), .I1(ram[564]), .I2(ram[556]), .I3(ram[548]), .S0(n27182), .S1(n26707), .ZN(n23371) );
  MUX41 U8503 ( .I0(ram[636]), .I1(ram[628]), .I2(ram[620]), .I3(ram[612]), .S0(n27182), .S1(n26707), .ZN(n23370) );
  MUX41 U8504 ( .I0(ram[7580]), .I1(ram[7572]), .I2(ram[7564]), .I3(
        ram[7556]), .S0(n27199), .S1(n26724), .ZN(n23664) );
  MUX41 U8505 ( .I0(ram[7324]), .I1(ram[7316]), .I2(ram[7308]), .I3(
        ram[7300]), .S0(n27199), .S1(n26724), .ZN(n23654) );
  MUX41 U8506 ( .I0(ram[7196]), .I1(ram[7188]), .I2(ram[7180]), .I3(
        ram[7172]), .S0(n27198), .S1(n26723), .ZN(n23649) );
  MUX41 U8507 ( .I0(ram[5532]), .I1(ram[5524]), .I2(ram[5516]), .I3(
        ram[5508]), .S0(n27194), .S1(n26719), .ZN(n23579) );
  MUX41 U8508 ( .I0(ram[11676]), .I1(ram[11668]), .I2(ram[11660]), .I3(
        ram[11652]), .S0(n27209), .S1(n26734), .ZN(n23835) );
  MUX41 U8509 ( .I0(ram[11420]), .I1(ram[11412]), .I2(ram[11404]), .I3(
        ram[11396]), .S0(n27208), .S1(n26733), .ZN(n23825) );
  MUX41 U8510 ( .I0(ram[11292]), .I1(ram[11284]), .I2(ram[11276]), .I3(
        ram[11268]), .S0(n27208), .S1(n26733), .ZN(n23820) );
  MUX41 U8511 ( .I0(ram[9628]), .I1(ram[9620]), .I2(ram[9612]), .I3(
        ram[9604]), .S0(n27204), .S1(n26729), .ZN(n23750) );
  MUX41 U8512 ( .I0(ram[9372]), .I1(ram[9364]), .I2(ram[9356]), .I3(
        ram[9348]), .S0(n27203), .S1(n26728), .ZN(n23740) );
  MUX41 U8513 ( .I0(ram[9244]), .I1(ram[9236]), .I2(ram[9228]), .I3(
        ram[9220]), .S0(n27203), .S1(n26728), .ZN(n23735) );
  MUX41 U8514 ( .I0(ram[15773]), .I1(ram[15765]), .I2(ram[15757]), .I3(
        ram[15749]), .S0(n27258), .S1(n26783), .ZN(n24690) );
  MUX41 U8515 ( .I0(ram[15517]), .I1(ram[15509]), .I2(ram[15501]), .I3(
        ram[15493]), .S0(n27258), .S1(n26783), .ZN(n24680) );
  MUX41 U8516 ( .I0(ram[15389]), .I1(ram[15381]), .I2(ram[15373]), .I3(
        ram[15365]), .S0(n27257), .S1(n26782), .ZN(n24675) );
  MUX41 U8517 ( .I0(ram[13725]), .I1(ram[13717]), .I2(ram[13709]), .I3(
        ram[13701]), .S0(n27253), .S1(n26778), .ZN(n24605) );
  MUX41 U8518 ( .I0(ram[13469]), .I1(ram[13461]), .I2(ram[13453]), .I3(
        ram[13445]), .S0(n27253), .S1(n26778), .ZN(n24595) );
  MUX41 U8519 ( .I0(ram[13341]), .I1(ram[13333]), .I2(ram[13325]), .I3(
        ram[13317]), .S0(n27252), .S1(n26777), .ZN(n24590) );
  MUX41 U8520 ( .I0(n24054), .I1(n24055), .I2(n24056), .I3(n24057), .S0(
        n26243), .S1(n26361), .ZN(n24053) );
  MUX41 U8521 ( .I0(ram[541]), .I1(ram[533]), .I2(ram[525]), .I3(ram[517]), .S0(n27222), .S1(n26747), .ZN(n24057) );
  MUX41 U8522 ( .I0(ram[573]), .I1(ram[565]), .I2(ram[557]), .I3(ram[549]), .S0(n27222), .S1(n26747), .ZN(n24055) );
  MUX41 U8523 ( .I0(ram[637]), .I1(ram[629]), .I2(ram[621]), .I3(ram[613]), .S0(n27222), .S1(n26747), .ZN(n24054) );
  MUX41 U8524 ( .I0(ram[7581]), .I1(ram[7573]), .I2(ram[7565]), .I3(
        ram[7557]), .S0(n27239), .S1(n26764), .ZN(n24348) );
  MUX41 U8525 ( .I0(ram[7325]), .I1(ram[7317]), .I2(ram[7309]), .I3(
        ram[7301]), .S0(n27238), .S1(n26763), .ZN(n24338) );
  MUX41 U8526 ( .I0(ram[7197]), .I1(ram[7189]), .I2(ram[7181]), .I3(
        ram[7173]), .S0(n27238), .S1(n26763), .ZN(n24333) );
  MUX41 U8527 ( .I0(ram[5533]), .I1(ram[5525]), .I2(ram[5517]), .I3(
        ram[5509]), .S0(n27234), .S1(n26759), .ZN(n24263) );
  MUX41 U8528 ( .I0(ram[11677]), .I1(ram[11669]), .I2(ram[11661]), .I3(
        ram[11653]), .S0(n27248), .S1(n26773), .ZN(n24519) );
  MUX41 U8529 ( .I0(ram[11421]), .I1(ram[11413]), .I2(ram[11405]), .I3(
        ram[11397]), .S0(n27248), .S1(n26773), .ZN(n24509) );
  MUX41 U8530 ( .I0(ram[11293]), .I1(ram[11285]), .I2(ram[11277]), .I3(
        ram[11269]), .S0(n27247), .S1(n26772), .ZN(n24504) );
  MUX41 U8531 ( .I0(ram[9629]), .I1(ram[9621]), .I2(ram[9613]), .I3(
        ram[9605]), .S0(n27243), .S1(n26768), .ZN(n24434) );
  MUX41 U8532 ( .I0(ram[9373]), .I1(ram[9365]), .I2(ram[9357]), .I3(
        ram[9349]), .S0(n27243), .S1(n26768), .ZN(n24424) );
  MUX41 U8533 ( .I0(ram[9245]), .I1(ram[9237]), .I2(ram[9229]), .I3(
        ram[9221]), .S0(n27243), .S1(n26768), .ZN(n24419) );
  MUX41 U8534 ( .I0(ram[15774]), .I1(ram[15766]), .I2(ram[15758]), .I3(
        ram[15750]), .S0(n27298), .S1(n26823), .ZN(n25374) );
  MUX41 U8535 ( .I0(ram[15518]), .I1(ram[15510]), .I2(ram[15502]), .I3(
        ram[15494]), .S0(n27297), .S1(n26822), .ZN(n25364) );
  MUX41 U8536 ( .I0(ram[15390]), .I1(ram[15382]), .I2(ram[15374]), .I3(
        ram[15366]), .S0(n27297), .S1(n26822), .ZN(n25359) );
  MUX41 U8537 ( .I0(ram[13726]), .I1(ram[13718]), .I2(ram[13710]), .I3(
        ram[13702]), .S0(n27293), .S1(n26818), .ZN(n25289) );
  MUX41 U8538 ( .I0(ram[13470]), .I1(ram[13462]), .I2(ram[13454]), .I3(
        ram[13446]), .S0(n27292), .S1(n26817), .ZN(n25279) );
  MUX41 U8539 ( .I0(ram[13342]), .I1(ram[13334]), .I2(ram[13326]), .I3(
        ram[13318]), .S0(n27292), .S1(n26817), .ZN(n25274) );
  MUX41 U8540 ( .I0(n24738), .I1(n24739), .I2(n24740), .I3(n24741), .S0(
        n26253), .S1(n26371), .ZN(n24737) );
  MUX41 U8541 ( .I0(ram[542]), .I1(ram[534]), .I2(ram[526]), .I3(ram[518]), .S0(n27261), .S1(n26786), .ZN(n24741) );
  MUX41 U8542 ( .I0(ram[574]), .I1(ram[566]), .I2(ram[558]), .I3(ram[550]), .S0(n27261), .S1(n26786), .ZN(n24739) );
  MUX41 U8543 ( .I0(ram[638]), .I1(ram[630]), .I2(ram[622]), .I3(ram[614]), .S0(n27261), .S1(n26786), .ZN(n24738) );
  MUX41 U8544 ( .I0(ram[7582]), .I1(ram[7574]), .I2(ram[7566]), .I3(
        ram[7558]), .S0(n27278), .S1(n26803), .ZN(n25032) );
  MUX41 U8545 ( .I0(ram[7326]), .I1(ram[7318]), .I2(ram[7310]), .I3(
        ram[7302]), .S0(n27277), .S1(n26802), .ZN(n25022) );
  MUX41 U8546 ( .I0(ram[7198]), .I1(ram[7190]), .I2(ram[7182]), .I3(
        ram[7174]), .S0(n27277), .S1(n26802), .ZN(n25017) );
  MUX41 U8547 ( .I0(ram[5534]), .I1(ram[5526]), .I2(ram[5518]), .I3(
        ram[5510]), .S0(n27273), .S1(n26798), .ZN(n24947) );
  MUX41 U8548 ( .I0(ram[11678]), .I1(ram[11670]), .I2(ram[11662]), .I3(
        ram[11654]), .S0(n27288), .S1(n26813), .ZN(n25203) );
  MUX41 U8549 ( .I0(ram[11422]), .I1(ram[11414]), .I2(ram[11406]), .I3(
        ram[11398]), .S0(n27287), .S1(n26812), .ZN(n25193) );
  MUX41 U8550 ( .I0(ram[11294]), .I1(ram[11286]), .I2(ram[11278]), .I3(
        ram[11270]), .S0(n27287), .S1(n26812), .ZN(n25188) );
  MUX41 U8551 ( .I0(ram[9630]), .I1(ram[9622]), .I2(ram[9614]), .I3(
        ram[9606]), .S0(n27283), .S1(n26808), .ZN(n25118) );
  MUX41 U8552 ( .I0(ram[9374]), .I1(ram[9366]), .I2(ram[9358]), .I3(
        ram[9350]), .S0(n27282), .S1(n26807), .ZN(n25108) );
  MUX41 U8553 ( .I0(ram[9246]), .I1(ram[9238]), .I2(ram[9230]), .I3(
        ram[9222]), .S0(n27282), .S1(n26807), .ZN(n25103) );
  MUX41 U8554 ( .I0(ram[15775]), .I1(ram[15767]), .I2(ram[15759]), .I3(
        ram[15751]), .S0(n27337), .S1(n26862), .ZN(n26058) );
  MUX41 U8555 ( .I0(ram[15519]), .I1(ram[15511]), .I2(ram[15503]), .I3(
        ram[15495]), .S0(n27336), .S1(n26861), .ZN(n26048) );
  MUX41 U8556 ( .I0(ram[15391]), .I1(ram[15383]), .I2(ram[15375]), .I3(
        ram[15367]), .S0(n27336), .S1(n26861), .ZN(n26043) );
  MUX41 U8557 ( .I0(ram[13727]), .I1(ram[13719]), .I2(ram[13711]), .I3(
        ram[13703]), .S0(n27332), .S1(n26857), .ZN(n25973) );
  MUX41 U8558 ( .I0(ram[13471]), .I1(ram[13463]), .I2(ram[13455]), .I3(
        ram[13447]), .S0(n27331), .S1(n26856), .ZN(n25963) );
  MUX41 U8559 ( .I0(ram[13343]), .I1(ram[13335]), .I2(ram[13327]), .I3(
        ram[13319]), .S0(n27331), .S1(n26856), .ZN(n25958) );
  MUX41 U8560 ( .I0(n25422), .I1(n25423), .I2(n25424), .I3(n25425), .S0(
        n26263), .S1(n26381), .ZN(n25421) );
  MUX41 U8561 ( .I0(ram[543]), .I1(ram[535]), .I2(ram[527]), .I3(ram[519]), .S0(n27300), .S1(n26825), .ZN(n25425) );
  MUX41 U8562 ( .I0(ram[575]), .I1(ram[567]), .I2(ram[559]), .I3(ram[551]), .S0(n27300), .S1(n26825), .ZN(n25423) );
  MUX41 U8563 ( .I0(ram[639]), .I1(ram[631]), .I2(ram[623]), .I3(ram[615]), .S0(n27301), .S1(n26826), .ZN(n25422) );
  MUX41 U8564 ( .I0(ram[7583]), .I1(ram[7575]), .I2(ram[7567]), .I3(
        ram[7559]), .S0(n27317), .S1(n26842), .ZN(n25716) );
  MUX41 U8565 ( .I0(ram[7327]), .I1(ram[7319]), .I2(ram[7311]), .I3(
        ram[7303]), .S0(n27317), .S1(n26842), .ZN(n25706) );
  MUX41 U8566 ( .I0(ram[7199]), .I1(ram[7191]), .I2(ram[7183]), .I3(
        ram[7175]), .S0(n27316), .S1(n26841), .ZN(n25701) );
  MUX41 U8567 ( .I0(ram[5535]), .I1(ram[5527]), .I2(ram[5519]), .I3(
        ram[5511]), .S0(n27312), .S1(n26837), .ZN(n25631) );
  MUX41 U8568 ( .I0(ram[11679]), .I1(ram[11671]), .I2(ram[11663]), .I3(
        ram[11655]), .S0(n27327), .S1(n26852), .ZN(n25887) );
  MUX41 U8569 ( .I0(ram[11423]), .I1(ram[11415]), .I2(ram[11407]), .I3(
        ram[11399]), .S0(n27327), .S1(n26852), .ZN(n25877) );
  MUX41 U8570 ( .I0(ram[11295]), .I1(ram[11287]), .I2(ram[11279]), .I3(
        ram[11271]), .S0(n27326), .S1(n26851), .ZN(n25872) );
  MUX41 U8571 ( .I0(ram[9631]), .I1(ram[9623]), .I2(ram[9615]), .I3(
        ram[9607]), .S0(n27322), .S1(n26847), .ZN(n25802) );
  MUX41 U8572 ( .I0(ram[9375]), .I1(ram[9367]), .I2(ram[9359]), .I3(
        ram[9351]), .S0(n27322), .S1(n26847), .ZN(n25792) );
  MUX41 U8573 ( .I0(ram[9247]), .I1(ram[9239]), .I2(ram[9231]), .I3(
        ram[9223]), .S0(n27321), .S1(n26846), .ZN(n25787) );
  MUX41 U8574 ( .I0(n21272), .I1(n21273), .I2(n21274), .I3(n21275), .S0(
        n26203), .S1(n26321), .ZN(n21271) );
  MUX41 U8575 ( .I0(ram[15896]), .I1(ram[15888]), .I2(ram[15880]), .I3(
        ram[15872]), .S0(n27062), .S1(n26587), .ZN(n21275) );
  MUX41 U8576 ( .I0(ram[15928]), .I1(ram[15920]), .I2(ram[15912]), .I3(
        ram[15904]), .S0(n27062), .S1(n26587), .ZN(n21273) );
  MUX41 U8577 ( .I0(ram[15992]), .I1(ram[15984]), .I2(ram[15976]), .I3(
        ram[15968]), .S0(n27062), .S1(n26587), .ZN(n21272) );
  MUX41 U8578 ( .I0(n21232), .I1(n21233), .I2(n21234), .I3(n21235), .S0(
        n26203), .S1(n26321), .ZN(n21231) );
  MUX41 U8579 ( .I0(ram[14872]), .I1(ram[14864]), .I2(ram[14856]), .I3(
        ram[14848]), .S0(n27059), .S1(n26584), .ZN(n21235) );
  MUX41 U8580 ( .I0(ram[14904]), .I1(ram[14896]), .I2(ram[14888]), .I3(
        ram[14880]), .S0(n27059), .S1(n26584), .ZN(n21233) );
  MUX41 U8581 ( .I0(ram[14968]), .I1(ram[14960]), .I2(ram[14952]), .I3(
        ram[14944]), .S0(n27059), .S1(n26584), .ZN(n21232) );
  MUX41 U8582 ( .I0(n21212), .I1(n21213), .I2(n21214), .I3(n21215), .S0(
        n26202), .S1(n26320), .ZN(n21211) );
  MUX41 U8583 ( .I0(ram[14360]), .I1(ram[14352]), .I2(ram[14344]), .I3(
        ram[14336]), .S0(n27058), .S1(n26583), .ZN(n21215) );
  MUX41 U8584 ( .I0(ram[14392]), .I1(ram[14384]), .I2(ram[14376]), .I3(
        ram[14368]), .S0(n27058), .S1(n26583), .ZN(n21213) );
  MUX41 U8585 ( .I0(ram[14456]), .I1(ram[14448]), .I2(ram[14440]), .I3(
        ram[14432]), .S0(n27058), .S1(n26583), .ZN(n21212) );
  MUX41 U8586 ( .I0(n21187), .I1(n21188), .I2(n21189), .I3(n21190), .S0(
        n26202), .S1(n26320), .ZN(n21186) );
  MUX41 U8587 ( .I0(ram[13848]), .I1(ram[13840]), .I2(ram[13832]), .I3(
        ram[13824]), .S0(n27057), .S1(n26582), .ZN(n21190) );
  MUX41 U8588 ( .I0(ram[13880]), .I1(ram[13872]), .I2(ram[13864]), .I3(
        ram[13856]), .S0(n27057), .S1(n26582), .ZN(n21188) );
  MUX41 U8589 ( .I0(ram[13944]), .I1(ram[13936]), .I2(ram[13928]), .I3(
        ram[13920]), .S0(n27057), .S1(n26582), .ZN(n21187) );
  MUX41 U8590 ( .I0(n21147), .I1(n21148), .I2(n21149), .I3(n21150), .S0(
        n26201), .S1(n26319), .ZN(n21146) );
  MUX41 U8591 ( .I0(ram[12824]), .I1(ram[12816]), .I2(ram[12808]), .I3(
        ram[12800]), .S0(n27054), .S1(n26579), .ZN(n21150) );
  MUX41 U8592 ( .I0(ram[12856]), .I1(ram[12848]), .I2(ram[12840]), .I3(
        ram[12832]), .S0(n27054), .S1(n26579), .ZN(n21148) );
  MUX41 U8593 ( .I0(ram[12920]), .I1(ram[12912]), .I2(ram[12904]), .I3(
        ram[12896]), .S0(n27054), .S1(n26579), .ZN(n21147) );
  MUX41 U8594 ( .I0(n21127), .I1(n21128), .I2(n21129), .I3(n21130), .S0(
        n26201), .S1(n26319), .ZN(n21126) );
  MUX41 U8595 ( .I0(ram[12312]), .I1(ram[12304]), .I2(ram[12296]), .I3(
        ram[12288]), .S0(n27053), .S1(n26578), .ZN(n21130) );
  MUX41 U8596 ( .I0(ram[12344]), .I1(ram[12336]), .I2(ram[12328]), .I3(
        ram[12320]), .S0(n27053), .S1(n26578), .ZN(n21128) );
  MUX41 U8597 ( .I0(ram[12408]), .I1(ram[12400]), .I2(ram[12392]), .I3(
        ram[12384]), .S0(n27053), .S1(n26578), .ZN(n21127) );
  MUX41 U8598 ( .I0(n20930), .I1(n20931), .I2(n20932), .I3(n20933), .S0(
        n26198), .S1(n26316), .ZN(n20929) );
  MUX41 U8599 ( .I0(ram[7736]), .I1(ram[7728]), .I2(ram[7720]), .I3(
        ram[7712]), .S0(n27042), .S1(n26567), .ZN(n20931) );
  MUX41 U8600 ( .I0(ram[7704]), .I1(ram[7696]), .I2(ram[7688]), .I3(
        ram[7680]), .S0(n27042), .S1(n26567), .ZN(n20933) );
  MUX41 U8601 ( .I0(ram[7800]), .I1(ram[7792]), .I2(ram[7784]), .I3(
        ram[7776]), .S0(n27042), .S1(n26567), .ZN(n20930) );
  MUX41 U8602 ( .I0(n20870), .I1(n20871), .I2(n20872), .I3(n20873), .S0(
        n26197), .S1(n26315), .ZN(n20869) );
  MUX41 U8603 ( .I0(ram[6200]), .I1(ram[6192]), .I2(ram[6184]), .I3(
        ram[6176]), .S0(n27038), .S1(n26563), .ZN(n20871) );
  MUX41 U8604 ( .I0(ram[6168]), .I1(ram[6160]), .I2(ram[6152]), .I3(
        ram[6144]), .S0(n27038), .S1(n26563), .ZN(n20873) );
  MUX41 U8605 ( .I0(ram[6264]), .I1(ram[6256]), .I2(ram[6248]), .I3(
        ram[6240]), .S0(n27038), .S1(n26563), .ZN(n20870) );
  MUX41 U8606 ( .I0(n20845), .I1(n20846), .I2(n20847), .I3(n20848), .S0(
        n26197), .S1(n26315), .ZN(n20844) );
  MUX41 U8607 ( .I0(ram[5688]), .I1(ram[5680]), .I2(ram[5672]), .I3(
        ram[5664]), .S0(n27037), .S1(n26562), .ZN(n20846) );
  MUX41 U8608 ( .I0(ram[5656]), .I1(ram[5648]), .I2(ram[5640]), .I3(
        ram[5632]), .S0(n27037), .S1(n26562), .ZN(n20848) );
  MUX41 U8609 ( .I0(ram[5752]), .I1(ram[5744]), .I2(ram[5736]), .I3(
        ram[5728]), .S0(n27037), .S1(n26562), .ZN(n20845) );
  MUX41 U8610 ( .I0(n21101), .I1(n21102), .I2(n21103), .I3(n21104), .S0(
        n26201), .S1(n26319), .ZN(n21100) );
  MUX41 U8611 ( .I0(ram[11832]), .I1(ram[11824]), .I2(ram[11816]), .I3(
        ram[11808]), .S0(n27052), .S1(n26577), .ZN(n21102) );
  MUX41 U8612 ( .I0(ram[11800]), .I1(ram[11792]), .I2(ram[11784]), .I3(
        ram[11776]), .S0(n27052), .S1(n26577), .ZN(n21104) );
  MUX41 U8613 ( .I0(ram[11896]), .I1(ram[11888]), .I2(ram[11880]), .I3(
        ram[11872]), .S0(n27052), .S1(n26577), .ZN(n21101) );
  MUX41 U8614 ( .I0(n21041), .I1(n21042), .I2(n21043), .I3(n21044), .S0(
        n26200), .S1(n26318), .ZN(n21040) );
  MUX41 U8615 ( .I0(ram[10296]), .I1(ram[10288]), .I2(ram[10280]), .I3(
        ram[10272]), .S0(n27048), .S1(n26573), .ZN(n21042) );
  MUX41 U8616 ( .I0(ram[10264]), .I1(ram[10256]), .I2(ram[10248]), .I3(
        ram[10240]), .S0(n27048), .S1(n26573), .ZN(n21044) );
  MUX41 U8617 ( .I0(ram[10360]), .I1(ram[10352]), .I2(ram[10344]), .I3(
        ram[10336]), .S0(n27048), .S1(n26573), .ZN(n21041) );
  MUX41 U8618 ( .I0(n21016), .I1(n21017), .I2(n21018), .I3(n21019), .S0(
        n26200), .S1(n26318), .ZN(n21015) );
  MUX41 U8619 ( .I0(ram[9784]), .I1(ram[9776]), .I2(ram[9768]), .I3(
        ram[9760]), .S0(n27047), .S1(n26572), .ZN(n21017) );
  MUX41 U8620 ( .I0(ram[9752]), .I1(ram[9744]), .I2(ram[9736]), .I3(
        ram[9728]), .S0(n27047), .S1(n26572), .ZN(n21019) );
  MUX41 U8621 ( .I0(ram[9848]), .I1(ram[9840]), .I2(ram[9832]), .I3(
        ram[9824]), .S0(n27047), .S1(n26572), .ZN(n21016) );
  MUX41 U8622 ( .I0(n21956), .I1(n21957), .I2(n21958), .I3(n21959), .S0(
        n26213), .S1(n26331), .ZN(n21955) );
  MUX41 U8623 ( .I0(ram[15929]), .I1(ram[15921]), .I2(ram[15913]), .I3(
        ram[15905]), .S0(n27101), .S1(n26626), .ZN(n21957) );
  MUX41 U8624 ( .I0(ram[15897]), .I1(ram[15889]), .I2(ram[15881]), .I3(
        ram[15873]), .S0(n27101), .S1(n26626), .ZN(n21959) );
  MUX41 U8625 ( .I0(ram[15993]), .I1(ram[15985]), .I2(ram[15977]), .I3(
        ram[15969]), .S0(n27101), .S1(n26626), .ZN(n21956) );
  MUX41 U8626 ( .I0(n21916), .I1(n21917), .I2(n21918), .I3(n21919), .S0(
        n26213), .S1(n26331), .ZN(n21915) );
  MUX41 U8627 ( .I0(ram[14873]), .I1(ram[14865]), .I2(ram[14857]), .I3(
        ram[14849]), .S0(n27099), .S1(n26624), .ZN(n21919) );
  MUX41 U8628 ( .I0(ram[14905]), .I1(ram[14897]), .I2(ram[14889]), .I3(
        ram[14881]), .S0(n27099), .S1(n26624), .ZN(n21917) );
  MUX41 U8629 ( .I0(ram[14969]), .I1(ram[14961]), .I2(ram[14953]), .I3(
        ram[14945]), .S0(n27099), .S1(n26624), .ZN(n21916) );
  MUX41 U8630 ( .I0(n21896), .I1(n21897), .I2(n21898), .I3(n21899), .S0(
        n26212), .S1(n26330), .ZN(n21895) );
  MUX41 U8631 ( .I0(ram[14361]), .I1(ram[14353]), .I2(ram[14345]), .I3(
        ram[14337]), .S0(n27097), .S1(n26622), .ZN(n21899) );
  MUX41 U8632 ( .I0(ram[14393]), .I1(ram[14385]), .I2(ram[14377]), .I3(
        ram[14369]), .S0(n27097), .S1(n26622), .ZN(n21897) );
  MUX41 U8633 ( .I0(ram[14457]), .I1(ram[14449]), .I2(ram[14441]), .I3(
        ram[14433]), .S0(n27098), .S1(n26623), .ZN(n21896) );
  MUX41 U8634 ( .I0(n21871), .I1(n21872), .I2(n21873), .I3(n21874), .S0(
        n26212), .S1(n26330), .ZN(n21870) );
  MUX41 U8635 ( .I0(ram[13849]), .I1(ram[13841]), .I2(ram[13833]), .I3(
        ram[13825]), .S0(n27096), .S1(n26621), .ZN(n21874) );
  MUX41 U8636 ( .I0(ram[13881]), .I1(ram[13873]), .I2(ram[13865]), .I3(
        ram[13857]), .S0(n27096), .S1(n26621), .ZN(n21872) );
  MUX41 U8637 ( .I0(ram[13945]), .I1(ram[13937]), .I2(ram[13929]), .I3(
        ram[13921]), .S0(n27096), .S1(n26621), .ZN(n21871) );
  MUX41 U8638 ( .I0(n21831), .I1(n21832), .I2(n21833), .I3(n21834), .S0(
        n26211), .S1(n26329), .ZN(n21830) );
  MUX41 U8639 ( .I0(ram[12825]), .I1(ram[12817]), .I2(ram[12809]), .I3(
        ram[12801]), .S0(n27094), .S1(n26619), .ZN(n21834) );
  MUX41 U8640 ( .I0(ram[12857]), .I1(ram[12849]), .I2(ram[12841]), .I3(
        ram[12833]), .S0(n27094), .S1(n26619), .ZN(n21832) );
  MUX41 U8641 ( .I0(ram[12921]), .I1(ram[12913]), .I2(ram[12905]), .I3(
        ram[12897]), .S0(n27094), .S1(n26619), .ZN(n21831) );
  MUX41 U8642 ( .I0(n21811), .I1(n21812), .I2(n21813), .I3(n21814), .S0(
        n26211), .S1(n26329), .ZN(n21810) );
  MUX41 U8643 ( .I0(ram[12313]), .I1(ram[12305]), .I2(ram[12297]), .I3(
        ram[12289]), .S0(n27092), .S1(n26617), .ZN(n21814) );
  MUX41 U8644 ( .I0(ram[12345]), .I1(ram[12337]), .I2(ram[12329]), .I3(
        ram[12321]), .S0(n27092), .S1(n26617), .ZN(n21812) );
  MUX41 U8645 ( .I0(ram[12409]), .I1(ram[12401]), .I2(ram[12393]), .I3(
        ram[12385]), .S0(n27093), .S1(n26618), .ZN(n21811) );
  MUX41 U8646 ( .I0(n21614), .I1(n21615), .I2(n21616), .I3(n21617), .S0(
        n26208), .S1(n26326), .ZN(n21613) );
  MUX41 U8647 ( .I0(ram[7737]), .I1(ram[7729]), .I2(ram[7721]), .I3(
        ram[7713]), .S0(n27081), .S1(n26606), .ZN(n21615) );
  MUX41 U8648 ( .I0(ram[7705]), .I1(ram[7697]), .I2(ram[7689]), .I3(
        ram[7681]), .S0(n27081), .S1(n26606), .ZN(n21617) );
  MUX41 U8649 ( .I0(ram[7801]), .I1(ram[7793]), .I2(ram[7785]), .I3(
        ram[7777]), .S0(n27082), .S1(n26607), .ZN(n21614) );
  MUX41 U8650 ( .I0(n21554), .I1(n21555), .I2(n21556), .I3(n21557), .S0(
        n26207), .S1(n26325), .ZN(n21553) );
  MUX41 U8651 ( .I0(ram[6201]), .I1(ram[6193]), .I2(ram[6185]), .I3(
        ram[6177]), .S0(n27078), .S1(n26603), .ZN(n21555) );
  MUX41 U8652 ( .I0(ram[6169]), .I1(ram[6161]), .I2(ram[6153]), .I3(
        ram[6145]), .S0(n27078), .S1(n26603), .ZN(n21557) );
  MUX41 U8653 ( .I0(ram[6265]), .I1(ram[6257]), .I2(ram[6249]), .I3(
        ram[6241]), .S0(n27078), .S1(n26603), .ZN(n21554) );
  MUX41 U8654 ( .I0(n21529), .I1(n21530), .I2(n21531), .I3(n21532), .S0(
        n26207), .S1(n26325), .ZN(n21528) );
  MUX41 U8655 ( .I0(ram[5689]), .I1(ram[5681]), .I2(ram[5673]), .I3(
        ram[5665]), .S0(n27076), .S1(n26601), .ZN(n21530) );
  MUX41 U8656 ( .I0(ram[5657]), .I1(ram[5649]), .I2(ram[5641]), .I3(
        ram[5633]), .S0(n27076), .S1(n26601), .ZN(n21532) );
  MUX41 U8657 ( .I0(ram[5753]), .I1(ram[5745]), .I2(ram[5737]), .I3(
        ram[5729]), .S0(n27077), .S1(n26602), .ZN(n21529) );
  MUX41 U8658 ( .I0(n21785), .I1(n21786), .I2(n21787), .I3(n21788), .S0(
        n26211), .S1(n26329), .ZN(n21784) );
  MUX41 U8659 ( .I0(ram[11833]), .I1(ram[11825]), .I2(ram[11817]), .I3(
        ram[11809]), .S0(n27091), .S1(n26616), .ZN(n21786) );
  MUX41 U8660 ( .I0(ram[11801]), .I1(ram[11793]), .I2(ram[11785]), .I3(
        ram[11777]), .S0(n27091), .S1(n26616), .ZN(n21788) );
  MUX41 U8661 ( .I0(ram[11897]), .I1(ram[11889]), .I2(ram[11881]), .I3(
        ram[11873]), .S0(n27091), .S1(n26616), .ZN(n21785) );
  MUX41 U8662 ( .I0(n21725), .I1(n21726), .I2(n21727), .I3(n21728), .S0(
        n26210), .S1(n26328), .ZN(n21724) );
  MUX41 U8663 ( .I0(ram[10297]), .I1(ram[10289]), .I2(ram[10281]), .I3(
        ram[10273]), .S0(n27088), .S1(n26613), .ZN(n21726) );
  MUX41 U8664 ( .I0(ram[10265]), .I1(ram[10257]), .I2(ram[10249]), .I3(
        ram[10241]), .S0(n27087), .S1(n26612), .ZN(n21728) );
  MUX41 U8665 ( .I0(ram[10361]), .I1(ram[10353]), .I2(ram[10345]), .I3(
        ram[10337]), .S0(n27088), .S1(n26613), .ZN(n21725) );
  MUX41 U8666 ( .I0(n21700), .I1(n21701), .I2(n21702), .I3(n21703), .S0(
        n26209), .S1(n26327), .ZN(n21699) );
  MUX41 U8667 ( .I0(ram[9785]), .I1(ram[9777]), .I2(ram[9769]), .I3(
        ram[9761]), .S0(n27086), .S1(n26611), .ZN(n21701) );
  MUX41 U8668 ( .I0(ram[9753]), .I1(ram[9745]), .I2(ram[9737]), .I3(
        ram[9729]), .S0(n27086), .S1(n26611), .ZN(n21703) );
  MUX41 U8669 ( .I0(ram[9849]), .I1(ram[9841]), .I2(ram[9833]), .I3(
        ram[9825]), .S0(n27086), .S1(n26611), .ZN(n21700) );
  MUX41 U8670 ( .I0(n22640), .I1(n22641), .I2(n22642), .I3(n22643), .S0(
        n26223), .S1(n26341), .ZN(n22639) );
  MUX41 U8671 ( .I0(ram[15930]), .I1(ram[15922]), .I2(ram[15914]), .I3(
        ram[15906]), .S0(n27140), .S1(n26665), .ZN(n22641) );
  MUX41 U8672 ( .I0(ram[15898]), .I1(ram[15890]), .I2(ram[15882]), .I3(
        ram[15874]), .S0(n27140), .S1(n26665), .ZN(n22643) );
  MUX41 U8673 ( .I0(ram[15994]), .I1(ram[15986]), .I2(ram[15978]), .I3(
        ram[15970]), .S0(n27141), .S1(n26666), .ZN(n22640) );
  MUX41 U8674 ( .I0(n22600), .I1(n22601), .I2(n22602), .I3(n22603), .S0(
        n26222), .S1(n26340), .ZN(n22599) );
  MUX41 U8675 ( .I0(ram[14874]), .I1(ram[14866]), .I2(ram[14858]), .I3(
        ram[14850]), .S0(n27138), .S1(n26663), .ZN(n22603) );
  MUX41 U8676 ( .I0(ram[14906]), .I1(ram[14898]), .I2(ram[14890]), .I3(
        ram[14882]), .S0(n27138), .S1(n26663), .ZN(n22601) );
  MUX41 U8677 ( .I0(ram[14970]), .I1(ram[14962]), .I2(ram[14954]), .I3(
        ram[14946]), .S0(n27138), .S1(n26663), .ZN(n22600) );
  MUX41 U8678 ( .I0(n22580), .I1(n22581), .I2(n22582), .I3(n22583), .S0(
        n26222), .S1(n26340), .ZN(n22579) );
  MUX41 U8679 ( .I0(ram[14362]), .I1(ram[14354]), .I2(ram[14346]), .I3(
        ram[14338]), .S0(n27137), .S1(n26662), .ZN(n22583) );
  MUX41 U8680 ( .I0(ram[14394]), .I1(ram[14386]), .I2(ram[14378]), .I3(
        ram[14370]), .S0(n27137), .S1(n26662), .ZN(n22581) );
  MUX41 U8681 ( .I0(ram[14458]), .I1(ram[14450]), .I2(ram[14442]), .I3(
        ram[14434]), .S0(n27137), .S1(n26662), .ZN(n22580) );
  MUX41 U8682 ( .I0(n22555), .I1(n22556), .I2(n22557), .I3(n22558), .S0(
        n26222), .S1(n26340), .ZN(n22554) );
  MUX41 U8683 ( .I0(ram[13850]), .I1(ram[13842]), .I2(ram[13834]), .I3(
        ram[13826]), .S0(n27135), .S1(n26660), .ZN(n22558) );
  MUX41 U8684 ( .I0(ram[13882]), .I1(ram[13874]), .I2(ram[13866]), .I3(
        ram[13858]), .S0(n27136), .S1(n26661), .ZN(n22556) );
  MUX41 U8685 ( .I0(ram[13946]), .I1(ram[13938]), .I2(ram[13930]), .I3(
        ram[13922]), .S0(n27136), .S1(n26661), .ZN(n22555) );
  MUX41 U8686 ( .I0(n22515), .I1(n22516), .I2(n22517), .I3(n22518), .S0(
        n26221), .S1(n26339), .ZN(n22514) );
  MUX41 U8687 ( .I0(ram[12826]), .I1(ram[12818]), .I2(ram[12810]), .I3(
        ram[12802]), .S0(n27133), .S1(n26658), .ZN(n22518) );
  MUX41 U8688 ( .I0(ram[12858]), .I1(ram[12850]), .I2(ram[12842]), .I3(
        ram[12834]), .S0(n27133), .S1(n26658), .ZN(n22516) );
  MUX41 U8689 ( .I0(ram[12922]), .I1(ram[12914]), .I2(ram[12906]), .I3(
        ram[12898]), .S0(n27133), .S1(n26658), .ZN(n22515) );
  MUX41 U8690 ( .I0(n22495), .I1(n22496), .I2(n22497), .I3(n22498), .S0(
        n26221), .S1(n26339), .ZN(n22494) );
  MUX41 U8691 ( .I0(ram[12314]), .I1(ram[12306]), .I2(ram[12298]), .I3(
        ram[12290]), .S0(n27132), .S1(n26657), .ZN(n22498) );
  MUX41 U8692 ( .I0(ram[12346]), .I1(ram[12338]), .I2(ram[12330]), .I3(
        ram[12322]), .S0(n27132), .S1(n26657), .ZN(n22496) );
  MUX41 U8693 ( .I0(ram[12410]), .I1(ram[12402]), .I2(ram[12394]), .I3(
        ram[12386]), .S0(n27132), .S1(n26657), .ZN(n22495) );
  MUX41 U8694 ( .I0(n22298), .I1(n22299), .I2(n22300), .I3(n22301), .S0(
        n26218), .S1(n26336), .ZN(n22297) );
  MUX41 U8695 ( .I0(ram[7738]), .I1(ram[7730]), .I2(ram[7722]), .I3(
        ram[7714]), .S0(n27121), .S1(n26646), .ZN(n22299) );
  MUX41 U8696 ( .I0(ram[7706]), .I1(ram[7698]), .I2(ram[7690]), .I3(
        ram[7682]), .S0(n27121), .S1(n26646), .ZN(n22301) );
  MUX41 U8697 ( .I0(ram[7802]), .I1(ram[7794]), .I2(ram[7786]), .I3(
        ram[7778]), .S0(n27121), .S1(n26646), .ZN(n22298) );
  MUX41 U8698 ( .I0(n22238), .I1(n22239), .I2(n22240), .I3(n22241), .S0(
        n26217), .S1(n26335), .ZN(n22237) );
  MUX41 U8699 ( .I0(ram[6202]), .I1(ram[6194]), .I2(ram[6186]), .I3(
        ram[6178]), .S0(n27117), .S1(n26642), .ZN(n22239) );
  MUX41 U8700 ( .I0(ram[6170]), .I1(ram[6162]), .I2(ram[6154]), .I3(
        ram[6146]), .S0(n27117), .S1(n26642), .ZN(n22241) );
  MUX41 U8701 ( .I0(ram[6266]), .I1(ram[6258]), .I2(ram[6250]), .I3(
        ram[6242]), .S0(n27117), .S1(n26642), .ZN(n22238) );
  MUX41 U8702 ( .I0(n22258), .I1(n22259), .I2(n22260), .I3(n22261), .S0(
        n26217), .S1(n26335), .ZN(n22257) );
  MUX41 U8703 ( .I0(ram[6682]), .I1(ram[6674]), .I2(ram[6666]), .I3(
        ram[6658]), .S0(n27118), .S1(n26643), .ZN(n22261) );
  MUX41 U8704 ( .I0(ram[6714]), .I1(ram[6706]), .I2(ram[6698]), .I3(
        ram[6690]), .S0(n27118), .S1(n26643), .ZN(n22259) );
  MUX41 U8705 ( .I0(ram[6778]), .I1(ram[6770]), .I2(ram[6762]), .I3(
        ram[6754]), .S0(n27118), .S1(n26643), .ZN(n22258) );
  MUX41 U8706 ( .I0(n22213), .I1(n22214), .I2(n22215), .I3(n22216), .S0(
        n26217), .S1(n26335), .ZN(n22212) );
  MUX41 U8707 ( .I0(ram[5690]), .I1(ram[5682]), .I2(ram[5674]), .I3(
        ram[5666]), .S0(n27116), .S1(n26641), .ZN(n22214) );
  MUX41 U8708 ( .I0(ram[5658]), .I1(ram[5650]), .I2(ram[5642]), .I3(
        ram[5634]), .S0(n27116), .S1(n26641), .ZN(n22216) );
  MUX41 U8709 ( .I0(ram[5754]), .I1(ram[5746]), .I2(ram[5738]), .I3(
        ram[5730]), .S0(n27116), .S1(n26641), .ZN(n22213) );
  MUX41 U8710 ( .I0(n22469), .I1(n22470), .I2(n22471), .I3(n22472), .S0(
        n26221), .S1(n26339), .ZN(n22468) );
  MUX41 U8711 ( .I0(ram[11834]), .I1(ram[11826]), .I2(ram[11818]), .I3(
        ram[11810]), .S0(n27131), .S1(n26656), .ZN(n22470) );
  MUX41 U8712 ( .I0(ram[11802]), .I1(ram[11794]), .I2(ram[11786]), .I3(
        ram[11778]), .S0(n27131), .S1(n26656), .ZN(n22472) );
  MUX41 U8713 ( .I0(ram[11898]), .I1(ram[11890]), .I2(ram[11882]), .I3(
        ram[11874]), .S0(n27131), .S1(n26656), .ZN(n22469) );
  MUX41 U8714 ( .I0(n22409), .I1(n22410), .I2(n22411), .I3(n22412), .S0(
        n26220), .S1(n26338), .ZN(n22408) );
  MUX41 U8715 ( .I0(ram[10298]), .I1(ram[10290]), .I2(ram[10282]), .I3(
        ram[10274]), .S0(n27127), .S1(n26652), .ZN(n22410) );
  MUX41 U8716 ( .I0(ram[10266]), .I1(ram[10258]), .I2(ram[10250]), .I3(
        ram[10242]), .S0(n27127), .S1(n26652), .ZN(n22412) );
  MUX41 U8717 ( .I0(ram[10362]), .I1(ram[10354]), .I2(ram[10346]), .I3(
        ram[10338]), .S0(n27127), .S1(n26652), .ZN(n22409) );
  MUX41 U8718 ( .I0(n22384), .I1(n22385), .I2(n22386), .I3(n22387), .S0(
        n26219), .S1(n26337), .ZN(n22383) );
  MUX41 U8719 ( .I0(ram[9786]), .I1(ram[9778]), .I2(ram[9770]), .I3(
        ram[9762]), .S0(n27126), .S1(n26651), .ZN(n22385) );
  MUX41 U8720 ( .I0(ram[9754]), .I1(ram[9746]), .I2(ram[9738]), .I3(
        ram[9730]), .S0(n27126), .S1(n26651), .ZN(n22387) );
  MUX41 U8721 ( .I0(ram[9850]), .I1(ram[9842]), .I2(ram[9834]), .I3(
        ram[9826]), .S0(n27126), .S1(n26651), .ZN(n22384) );
  MUX41 U8722 ( .I0(n22324), .I1(n22325), .I2(n22326), .I3(n22327), .S0(
        n26218), .S1(n26336), .ZN(n22323) );
  MUX41 U8723 ( .I0(ram[8250]), .I1(ram[8242]), .I2(ram[8234]), .I3(
        ram[8226]), .S0(n27122), .S1(n26647), .ZN(n22325) );
  MUX41 U8724 ( .I0(ram[8218]), .I1(ram[8210]), .I2(ram[8202]), .I3(
        ram[8194]), .S0(n27122), .S1(n26647), .ZN(n22327) );
  MUX41 U8725 ( .I0(ram[8314]), .I1(ram[8306]), .I2(ram[8298]), .I3(
        ram[8290]), .S0(n27122), .S1(n26647), .ZN(n22324) );
  MUX41 U8726 ( .I0(n23324), .I1(n23325), .I2(n23326), .I3(n23327), .S0(
        n26233), .S1(n26351), .ZN(n23323) );
  MUX41 U8727 ( .I0(ram[15931]), .I1(ram[15923]), .I2(ram[15915]), .I3(
        ram[15907]), .S0(n27180), .S1(n26705), .ZN(n23325) );
  MUX41 U8728 ( .I0(ram[15899]), .I1(ram[15891]), .I2(ram[15883]), .I3(
        ram[15875]), .S0(n27180), .S1(n26705), .ZN(n23327) );
  MUX41 U8729 ( .I0(ram[15995]), .I1(ram[15987]), .I2(ram[15979]), .I3(
        ram[15971]), .S0(n27180), .S1(n26705), .ZN(n23324) );
  MUX41 U8730 ( .I0(n23284), .I1(n23285), .I2(n23286), .I3(n23287), .S0(
        n26232), .S1(n26350), .ZN(n23283) );
  MUX41 U8731 ( .I0(ram[14875]), .I1(ram[14867]), .I2(ram[14859]), .I3(
        ram[14851]), .S0(n27177), .S1(n26702), .ZN(n23287) );
  MUX41 U8732 ( .I0(ram[14907]), .I1(ram[14899]), .I2(ram[14891]), .I3(
        ram[14883]), .S0(n27177), .S1(n26702), .ZN(n23285) );
  MUX41 U8733 ( .I0(ram[14971]), .I1(ram[14963]), .I2(ram[14955]), .I3(
        ram[14947]), .S0(n27178), .S1(n26703), .ZN(n23284) );
  MUX41 U8734 ( .I0(n23264), .I1(n23265), .I2(n23266), .I3(n23267), .S0(
        n26232), .S1(n26350), .ZN(n23263) );
  MUX41 U8735 ( .I0(ram[14363]), .I1(ram[14355]), .I2(ram[14347]), .I3(
        ram[14339]), .S0(n27176), .S1(n26701), .ZN(n23267) );
  MUX41 U8736 ( .I0(ram[14395]), .I1(ram[14387]), .I2(ram[14379]), .I3(
        ram[14371]), .S0(n27176), .S1(n26701), .ZN(n23265) );
  MUX41 U8737 ( .I0(ram[14459]), .I1(ram[14451]), .I2(ram[14443]), .I3(
        ram[14435]), .S0(n27176), .S1(n26701), .ZN(n23264) );
  MUX41 U8738 ( .I0(n23239), .I1(n23240), .I2(n23241), .I3(n23242), .S0(
        n26232), .S1(n26350), .ZN(n23238) );
  MUX41 U8739 ( .I0(ram[13851]), .I1(ram[13843]), .I2(ram[13835]), .I3(
        ram[13827]), .S0(n27175), .S1(n26700), .ZN(n23242) );
  MUX41 U8740 ( .I0(ram[13883]), .I1(ram[13875]), .I2(ram[13867]), .I3(
        ram[13859]), .S0(n27175), .S1(n26700), .ZN(n23240) );
  MUX41 U8741 ( .I0(ram[13947]), .I1(ram[13939]), .I2(ram[13931]), .I3(
        ram[13923]), .S0(n27175), .S1(n26700), .ZN(n23239) );
  MUX41 U8742 ( .I0(n23199), .I1(n23200), .I2(n23201), .I3(n23202), .S0(
        n26231), .S1(n26349), .ZN(n23198) );
  MUX41 U8743 ( .I0(ram[12827]), .I1(ram[12819]), .I2(ram[12811]), .I3(
        ram[12803]), .S0(n27172), .S1(n26697), .ZN(n23202) );
  MUX41 U8744 ( .I0(ram[12859]), .I1(ram[12851]), .I2(ram[12843]), .I3(
        ram[12835]), .S0(n27172), .S1(n26697), .ZN(n23200) );
  MUX41 U8745 ( .I0(ram[12923]), .I1(ram[12915]), .I2(ram[12907]), .I3(
        ram[12899]), .S0(n27173), .S1(n26698), .ZN(n23199) );
  MUX41 U8746 ( .I0(n23179), .I1(n23180), .I2(n23181), .I3(n23182), .S0(
        n26231), .S1(n26349), .ZN(n23178) );
  MUX41 U8747 ( .I0(ram[12315]), .I1(ram[12307]), .I2(ram[12299]), .I3(
        ram[12291]), .S0(n27171), .S1(n26696), .ZN(n23182) );
  MUX41 U8748 ( .I0(ram[12347]), .I1(ram[12339]), .I2(ram[12331]), .I3(
        ram[12323]), .S0(n27171), .S1(n26696), .ZN(n23180) );
  MUX41 U8749 ( .I0(ram[12411]), .I1(ram[12403]), .I2(ram[12395]), .I3(
        ram[12387]), .S0(n27171), .S1(n26696), .ZN(n23179) );
  MUX41 U8750 ( .I0(n22982), .I1(n22983), .I2(n22984), .I3(n22985), .S0(
        n26228), .S1(n26346), .ZN(n22981) );
  MUX41 U8751 ( .I0(ram[7739]), .I1(ram[7731]), .I2(ram[7723]), .I3(
        ram[7715]), .S0(n27160), .S1(n26685), .ZN(n22983) );
  MUX41 U8752 ( .I0(ram[7707]), .I1(ram[7699]), .I2(ram[7691]), .I3(
        ram[7683]), .S0(n27160), .S1(n26685), .ZN(n22985) );
  MUX41 U8753 ( .I0(ram[7803]), .I1(ram[7795]), .I2(ram[7787]), .I3(
        ram[7779]), .S0(n27160), .S1(n26685), .ZN(n22982) );
  MUX41 U8754 ( .I0(n22922), .I1(n22923), .I2(n22924), .I3(n22925), .S0(
        n26227), .S1(n26345), .ZN(n22921) );
  MUX41 U8755 ( .I0(ram[6203]), .I1(ram[6195]), .I2(ram[6187]), .I3(
        ram[6179]), .S0(n27156), .S1(n26681), .ZN(n22923) );
  MUX41 U8756 ( .I0(ram[6171]), .I1(ram[6163]), .I2(ram[6155]), .I3(
        ram[6147]), .S0(n27156), .S1(n26681), .ZN(n22925) );
  MUX41 U8757 ( .I0(ram[6267]), .I1(ram[6259]), .I2(ram[6251]), .I3(
        ram[6243]), .S0(n27157), .S1(n26682), .ZN(n22922) );
  MUX41 U8758 ( .I0(n22942), .I1(n22943), .I2(n22944), .I3(n22945), .S0(
        n26227), .S1(n26345), .ZN(n22941) );
  MUX41 U8759 ( .I0(ram[6683]), .I1(ram[6675]), .I2(ram[6667]), .I3(
        ram[6659]), .S0(n27158), .S1(n26683), .ZN(n22945) );
  MUX41 U8760 ( .I0(ram[6715]), .I1(ram[6707]), .I2(ram[6699]), .I3(
        ram[6691]), .S0(n27158), .S1(n26683), .ZN(n22943) );
  MUX41 U8761 ( .I0(ram[6779]), .I1(ram[6771]), .I2(ram[6763]), .I3(
        ram[6755]), .S0(n27158), .S1(n26683), .ZN(n22942) );
  MUX41 U8762 ( .I0(n22897), .I1(n22898), .I2(n22899), .I3(n22900), .S0(
        n26227), .S1(n26345), .ZN(n22896) );
  MUX41 U8763 ( .I0(ram[5691]), .I1(ram[5683]), .I2(ram[5675]), .I3(
        ram[5667]), .S0(n27155), .S1(n26680), .ZN(n22898) );
  MUX41 U8764 ( .I0(ram[5659]), .I1(ram[5651]), .I2(ram[5643]), .I3(
        ram[5635]), .S0(n27155), .S1(n26680), .ZN(n22900) );
  MUX41 U8765 ( .I0(ram[5755]), .I1(ram[5747]), .I2(ram[5739]), .I3(
        ram[5731]), .S0(n27155), .S1(n26680), .ZN(n22897) );
  MUX41 U8766 ( .I0(n23153), .I1(n23154), .I2(n23155), .I3(n23156), .S0(
        n26230), .S1(n26348), .ZN(n23152) );
  MUX41 U8767 ( .I0(ram[11835]), .I1(ram[11827]), .I2(ram[11819]), .I3(
        ram[11811]), .S0(n27170), .S1(n26695), .ZN(n23154) );
  MUX41 U8768 ( .I0(ram[11803]), .I1(ram[11795]), .I2(ram[11787]), .I3(
        ram[11779]), .S0(n27170), .S1(n26695), .ZN(n23156) );
  MUX41 U8769 ( .I0(ram[11899]), .I1(ram[11891]), .I2(ram[11883]), .I3(
        ram[11875]), .S0(n27170), .S1(n26695), .ZN(n23153) );
  MUX41 U8770 ( .I0(n23093), .I1(n23094), .I2(n23095), .I3(n23096), .S0(
        n26229), .S1(n26347), .ZN(n23092) );
  MUX41 U8771 ( .I0(ram[10299]), .I1(ram[10291]), .I2(ram[10283]), .I3(
        ram[10275]), .S0(n27166), .S1(n26691), .ZN(n23094) );
  MUX41 U8772 ( .I0(ram[10267]), .I1(ram[10259]), .I2(ram[10251]), .I3(
        ram[10243]), .S0(n27166), .S1(n26691), .ZN(n23096) );
  MUX41 U8773 ( .I0(ram[10363]), .I1(ram[10355]), .I2(ram[10347]), .I3(
        ram[10339]), .S0(n27166), .S1(n26691), .ZN(n23093) );
  MUX41 U8774 ( .I0(n23068), .I1(n23069), .I2(n23070), .I3(n23071), .S0(
        n26229), .S1(n26347), .ZN(n23067) );
  MUX41 U8775 ( .I0(ram[9787]), .I1(ram[9779]), .I2(ram[9771]), .I3(
        ram[9763]), .S0(n27165), .S1(n26690), .ZN(n23069) );
  MUX41 U8776 ( .I0(ram[9755]), .I1(ram[9747]), .I2(ram[9739]), .I3(
        ram[9731]), .S0(n27165), .S1(n26690), .ZN(n23071) );
  MUX41 U8777 ( .I0(ram[9851]), .I1(ram[9843]), .I2(ram[9835]), .I3(
        ram[9827]), .S0(n27165), .S1(n26690), .ZN(n23068) );
  MUX41 U8778 ( .I0(n23008), .I1(n23009), .I2(n23010), .I3(n23011), .S0(
        n26228), .S1(n26346), .ZN(n23007) );
  MUX41 U8779 ( .I0(ram[8251]), .I1(ram[8243]), .I2(ram[8235]), .I3(
        ram[8227]), .S0(n27161), .S1(n26686), .ZN(n23009) );
  MUX41 U8780 ( .I0(ram[8219]), .I1(ram[8211]), .I2(ram[8203]), .I3(
        ram[8195]), .S0(n27161), .S1(n26686), .ZN(n23011) );
  MUX41 U8781 ( .I0(ram[8315]), .I1(ram[8307]), .I2(ram[8299]), .I3(
        ram[8291]), .S0(n27162), .S1(n26687), .ZN(n23008) );
  MUX41 U8782 ( .I0(n24008), .I1(n24009), .I2(n24010), .I3(n24011), .S0(
        n26243), .S1(n26361), .ZN(n24007) );
  MUX41 U8783 ( .I0(ram[15932]), .I1(ram[15924]), .I2(ram[15916]), .I3(
        ram[15908]), .S0(n27219), .S1(n26744), .ZN(n24009) );
  MUX41 U8784 ( .I0(ram[15900]), .I1(ram[15892]), .I2(ram[15884]), .I3(
        ram[15876]), .S0(n27219), .S1(n26744), .ZN(n24011) );
  MUX41 U8785 ( .I0(ram[15996]), .I1(ram[15988]), .I2(ram[15980]), .I3(
        ram[15972]), .S0(n27219), .S1(n26744), .ZN(n24008) );
  MUX41 U8786 ( .I0(n23968), .I1(n23969), .I2(n23970), .I3(n23971), .S0(
        n26242), .S1(n26360), .ZN(n23967) );
  MUX41 U8787 ( .I0(ram[14876]), .I1(ram[14868]), .I2(ram[14860]), .I3(
        ram[14852]), .S0(n27217), .S1(n26742), .ZN(n23971) );
  MUX41 U8788 ( .I0(ram[14908]), .I1(ram[14900]), .I2(ram[14892]), .I3(
        ram[14884]), .S0(n27217), .S1(n26742), .ZN(n23969) );
  MUX41 U8789 ( .I0(ram[14972]), .I1(ram[14964]), .I2(ram[14956]), .I3(
        ram[14948]), .S0(n27217), .S1(n26742), .ZN(n23968) );
  MUX41 U8790 ( .I0(n23948), .I1(n23949), .I2(n23950), .I3(n23951), .S0(
        n26242), .S1(n26360), .ZN(n23947) );
  MUX41 U8791 ( .I0(ram[14364]), .I1(ram[14356]), .I2(ram[14348]), .I3(
        ram[14340]), .S0(n27215), .S1(n26740), .ZN(n23951) );
  MUX41 U8792 ( .I0(ram[14396]), .I1(ram[14388]), .I2(ram[14380]), .I3(
        ram[14372]), .S0(n27216), .S1(n26741), .ZN(n23949) );
  MUX41 U8793 ( .I0(ram[14460]), .I1(ram[14452]), .I2(ram[14444]), .I3(
        ram[14436]), .S0(n27216), .S1(n26741), .ZN(n23948) );
  MUX41 U8794 ( .I0(n23923), .I1(n23924), .I2(n23925), .I3(n23926), .S0(
        n26241), .S1(n26359), .ZN(n23922) );
  MUX41 U8795 ( .I0(ram[13852]), .I1(ram[13844]), .I2(ram[13836]), .I3(
        ram[13828]), .S0(n27214), .S1(n26739), .ZN(n23926) );
  MUX41 U8796 ( .I0(ram[13884]), .I1(ram[13876]), .I2(ram[13868]), .I3(
        ram[13860]), .S0(n27214), .S1(n26739), .ZN(n23924) );
  MUX41 U8797 ( .I0(ram[13948]), .I1(ram[13940]), .I2(ram[13932]), .I3(
        ram[13924]), .S0(n27214), .S1(n26739), .ZN(n23923) );
  MUX41 U8798 ( .I0(n23883), .I1(n23884), .I2(n23885), .I3(n23886), .S0(
        n26241), .S1(n26359), .ZN(n23882) );
  MUX41 U8799 ( .I0(ram[12828]), .I1(ram[12820]), .I2(ram[12812]), .I3(
        ram[12804]), .S0(n27212), .S1(n26737), .ZN(n23886) );
  MUX41 U8800 ( .I0(ram[12860]), .I1(ram[12852]), .I2(ram[12844]), .I3(
        ram[12836]), .S0(n27212), .S1(n26737), .ZN(n23884) );
  MUX41 U8801 ( .I0(ram[12924]), .I1(ram[12916]), .I2(ram[12908]), .I3(
        ram[12900]), .S0(n27212), .S1(n26737), .ZN(n23883) );
  MUX41 U8802 ( .I0(n23863), .I1(n23864), .I2(n23865), .I3(n23866), .S0(
        n26241), .S1(n26359), .ZN(n23862) );
  MUX41 U8803 ( .I0(ram[12316]), .I1(ram[12308]), .I2(ram[12300]), .I3(
        ram[12292]), .S0(n27211), .S1(n26736), .ZN(n23866) );
  MUX41 U8804 ( .I0(ram[12348]), .I1(ram[12340]), .I2(ram[12332]), .I3(
        ram[12324]), .S0(n27211), .S1(n26736), .ZN(n23864) );
  MUX41 U8805 ( .I0(ram[12412]), .I1(ram[12404]), .I2(ram[12396]), .I3(
        ram[12388]), .S0(n27211), .S1(n26736), .ZN(n23863) );
  MUX41 U8806 ( .I0(n23666), .I1(n23667), .I2(n23668), .I3(n23669), .S0(
        n26238), .S1(n26356), .ZN(n23665) );
  MUX41 U8807 ( .I0(ram[7740]), .I1(ram[7732]), .I2(ram[7724]), .I3(
        ram[7716]), .S0(n27200), .S1(n26725), .ZN(n23667) );
  MUX41 U8808 ( .I0(ram[7708]), .I1(ram[7700]), .I2(ram[7692]), .I3(
        ram[7684]), .S0(n27199), .S1(n26724), .ZN(n23669) );
  MUX41 U8809 ( .I0(ram[7804]), .I1(ram[7796]), .I2(ram[7788]), .I3(
        ram[7780]), .S0(n27200), .S1(n26725), .ZN(n23666) );
  MUX41 U8810 ( .I0(n23606), .I1(n23607), .I2(n23608), .I3(n23609), .S0(
        n26237), .S1(n26355), .ZN(n23605) );
  MUX41 U8811 ( .I0(ram[6204]), .I1(ram[6196]), .I2(ram[6188]), .I3(
        ram[6180]), .S0(n27196), .S1(n26721), .ZN(n23607) );
  MUX41 U8812 ( .I0(ram[6172]), .I1(ram[6164]), .I2(ram[6156]), .I3(
        ram[6148]), .S0(n27196), .S1(n26721), .ZN(n23609) );
  MUX41 U8813 ( .I0(ram[6268]), .I1(ram[6260]), .I2(ram[6252]), .I3(
        ram[6244]), .S0(n27196), .S1(n26721), .ZN(n23606) );
  MUX41 U8814 ( .I0(n23626), .I1(n23627), .I2(n23628), .I3(n23629), .S0(
        n26237), .S1(n26355), .ZN(n23625) );
  MUX41 U8815 ( .I0(ram[6684]), .I1(ram[6676]), .I2(ram[6668]), .I3(
        ram[6660]), .S0(n27197), .S1(n26722), .ZN(n23629) );
  MUX41 U8816 ( .I0(ram[6716]), .I1(ram[6708]), .I2(ram[6700]), .I3(
        ram[6692]), .S0(n27197), .S1(n26722), .ZN(n23627) );
  MUX41 U8817 ( .I0(ram[6780]), .I1(ram[6772]), .I2(ram[6764]), .I3(
        ram[6756]), .S0(n27197), .S1(n26722), .ZN(n23626) );
  MUX41 U8818 ( .I0(n23581), .I1(n23582), .I2(n23583), .I3(n23584), .S0(
        n26237), .S1(n26355), .ZN(n23580) );
  MUX41 U8819 ( .I0(ram[5692]), .I1(ram[5684]), .I2(ram[5676]), .I3(
        ram[5668]), .S0(n27195), .S1(n26720), .ZN(n23582) );
  MUX41 U8820 ( .I0(ram[5660]), .I1(ram[5652]), .I2(ram[5644]), .I3(
        ram[5636]), .S0(n27195), .S1(n26720), .ZN(n23584) );
  MUX41 U8821 ( .I0(ram[5756]), .I1(ram[5748]), .I2(ram[5740]), .I3(
        ram[5732]), .S0(n27195), .S1(n26720), .ZN(n23581) );
  MUX41 U8822 ( .I0(n23837), .I1(n23838), .I2(n23839), .I3(n23840), .S0(
        n26240), .S1(n26358), .ZN(n23836) );
  MUX41 U8823 ( .I0(ram[11836]), .I1(ram[11828]), .I2(ram[11820]), .I3(
        ram[11812]), .S0(n27209), .S1(n26734), .ZN(n23838) );
  MUX41 U8824 ( .I0(ram[11804]), .I1(ram[11796]), .I2(ram[11788]), .I3(
        ram[11780]), .S0(n27209), .S1(n26734), .ZN(n23840) );
  MUX41 U8825 ( .I0(ram[11900]), .I1(ram[11892]), .I2(ram[11884]), .I3(
        ram[11876]), .S0(n27210), .S1(n26735), .ZN(n23837) );
  MUX41 U8826 ( .I0(n23777), .I1(n23778), .I2(n23779), .I3(n23780), .S0(
        n26239), .S1(n26357), .ZN(n23776) );
  MUX41 U8827 ( .I0(ram[10300]), .I1(ram[10292]), .I2(ram[10284]), .I3(
        ram[10276]), .S0(n27206), .S1(n26731), .ZN(n23778) );
  MUX41 U8828 ( .I0(ram[10268]), .I1(ram[10260]), .I2(ram[10252]), .I3(
        ram[10244]), .S0(n27206), .S1(n26731), .ZN(n23780) );
  MUX41 U8829 ( .I0(ram[10364]), .I1(ram[10356]), .I2(ram[10348]), .I3(
        ram[10340]), .S0(n27206), .S1(n26731), .ZN(n23777) );
  MUX41 U8830 ( .I0(n23752), .I1(n23753), .I2(n23754), .I3(n23755), .S0(
        n26239), .S1(n26357), .ZN(n23751) );
  MUX41 U8831 ( .I0(ram[9788]), .I1(ram[9780]), .I2(ram[9772]), .I3(
        ram[9764]), .S0(n27204), .S1(n26729), .ZN(n23753) );
  MUX41 U8832 ( .I0(ram[9756]), .I1(ram[9748]), .I2(ram[9740]), .I3(
        ram[9732]), .S0(n27204), .S1(n26729), .ZN(n23755) );
  MUX41 U8833 ( .I0(ram[9852]), .I1(ram[9844]), .I2(ram[9836]), .I3(
        ram[9828]), .S0(n27205), .S1(n26730), .ZN(n23752) );
  MUX41 U8834 ( .I0(n23692), .I1(n23693), .I2(n23694), .I3(n23695), .S0(
        n26238), .S1(n26356), .ZN(n23691) );
  MUX41 U8835 ( .I0(ram[8252]), .I1(ram[8244]), .I2(ram[8236]), .I3(
        ram[8228]), .S0(n27201), .S1(n26726), .ZN(n23693) );
  MUX41 U8836 ( .I0(ram[8220]), .I1(ram[8212]), .I2(ram[8204]), .I3(
        ram[8196]), .S0(n27201), .S1(n26726), .ZN(n23695) );
  MUX41 U8837 ( .I0(ram[8316]), .I1(ram[8308]), .I2(ram[8300]), .I3(
        ram[8292]), .S0(n27201), .S1(n26726), .ZN(n23692) );
  MUX41 U8838 ( .I0(n24692), .I1(n24693), .I2(n24694), .I3(n24695), .S0(
        n26253), .S1(n26371), .ZN(n24691) );
  MUX41 U8839 ( .I0(ram[15933]), .I1(ram[15925]), .I2(ram[15917]), .I3(
        ram[15909]), .S0(n27259), .S1(n26784), .ZN(n24693) );
  MUX41 U8840 ( .I0(ram[15901]), .I1(ram[15893]), .I2(ram[15885]), .I3(
        ram[15877]), .S0(n27259), .S1(n26784), .ZN(n24695) );
  MUX41 U8841 ( .I0(ram[15997]), .I1(ram[15989]), .I2(ram[15981]), .I3(
        ram[15973]), .S0(n27259), .S1(n26784), .ZN(n24692) );
  MUX41 U8842 ( .I0(n24652), .I1(n24653), .I2(n24654), .I3(n24655), .S0(
        n26252), .S1(n26370), .ZN(n24651) );
  MUX41 U8843 ( .I0(ram[14877]), .I1(ram[14869]), .I2(ram[14861]), .I3(
        ram[14853]), .S0(n27256), .S1(n26781), .ZN(n24655) );
  MUX41 U8844 ( .I0(ram[14909]), .I1(ram[14901]), .I2(ram[14893]), .I3(
        ram[14885]), .S0(n27256), .S1(n26781), .ZN(n24653) );
  MUX41 U8845 ( .I0(ram[14973]), .I1(ram[14965]), .I2(ram[14957]), .I3(
        ram[14949]), .S0(n27256), .S1(n26781), .ZN(n24652) );
  MUX41 U8846 ( .I0(n24632), .I1(n24633), .I2(n24634), .I3(n24635), .S0(
        n26252), .S1(n26370), .ZN(n24631) );
  MUX41 U8847 ( .I0(ram[14365]), .I1(ram[14357]), .I2(ram[14349]), .I3(
        ram[14341]), .S0(n27255), .S1(n26780), .ZN(n24635) );
  MUX41 U8848 ( .I0(ram[14397]), .I1(ram[14389]), .I2(ram[14381]), .I3(
        ram[14373]), .S0(n27255), .S1(n26780), .ZN(n24633) );
  MUX41 U8849 ( .I0(ram[14461]), .I1(ram[14453]), .I2(ram[14445]), .I3(
        ram[14437]), .S0(n27255), .S1(n26780), .ZN(n24632) );
  MUX41 U8850 ( .I0(n24607), .I1(n24608), .I2(n24609), .I3(n24610), .S0(
        n26251), .S1(n26369), .ZN(n24606) );
  MUX41 U8851 ( .I0(ram[13853]), .I1(ram[13845]), .I2(ram[13837]), .I3(
        ram[13829]), .S0(n27254), .S1(n26779), .ZN(n24610) );
  MUX41 U8852 ( .I0(ram[13885]), .I1(ram[13877]), .I2(ram[13869]), .I3(
        ram[13861]), .S0(n27254), .S1(n26779), .ZN(n24608) );
  MUX41 U8853 ( .I0(ram[13949]), .I1(ram[13941]), .I2(ram[13933]), .I3(
        ram[13925]), .S0(n27254), .S1(n26779), .ZN(n24607) );
  MUX41 U8854 ( .I0(n24567), .I1(n24568), .I2(n24569), .I3(n24570), .S0(
        n26251), .S1(n26369), .ZN(n24566) );
  MUX41 U8855 ( .I0(ram[12829]), .I1(ram[12821]), .I2(ram[12813]), .I3(
        ram[12805]), .S0(n27251), .S1(n26776), .ZN(n24570) );
  MUX41 U8856 ( .I0(ram[12861]), .I1(ram[12853]), .I2(ram[12845]), .I3(
        ram[12837]), .S0(n27251), .S1(n26776), .ZN(n24568) );
  MUX41 U8857 ( .I0(ram[12925]), .I1(ram[12917]), .I2(ram[12909]), .I3(
        ram[12901]), .S0(n27251), .S1(n26776), .ZN(n24567) );
  MUX41 U8858 ( .I0(n24547), .I1(n24548), .I2(n24549), .I3(n24550), .S0(
        n26250), .S1(n26368), .ZN(n24546) );
  MUX41 U8859 ( .I0(ram[12317]), .I1(ram[12309]), .I2(ram[12301]), .I3(
        ram[12293]), .S0(n27250), .S1(n26775), .ZN(n24550) );
  MUX41 U8860 ( .I0(ram[12349]), .I1(ram[12341]), .I2(ram[12333]), .I3(
        ram[12325]), .S0(n27250), .S1(n26775), .ZN(n24548) );
  MUX41 U8861 ( .I0(ram[12413]), .I1(ram[12405]), .I2(ram[12397]), .I3(
        ram[12389]), .S0(n27250), .S1(n26775), .ZN(n24547) );
  MUX41 U8862 ( .I0(n24350), .I1(n24351), .I2(n24352), .I3(n24353), .S0(
        n26248), .S1(n26366), .ZN(n24349) );
  MUX41 U8863 ( .I0(ram[7741]), .I1(ram[7733]), .I2(ram[7725]), .I3(
        ram[7717]), .S0(n27239), .S1(n26764), .ZN(n24351) );
  MUX41 U8864 ( .I0(ram[7709]), .I1(ram[7701]), .I2(ram[7693]), .I3(
        ram[7685]), .S0(n27239), .S1(n26764), .ZN(n24353) );
  MUX41 U8865 ( .I0(ram[7805]), .I1(ram[7797]), .I2(ram[7789]), .I3(
        ram[7781]), .S0(n27239), .S1(n26764), .ZN(n24350) );
  MUX41 U8866 ( .I0(n24290), .I1(n24291), .I2(n24292), .I3(n24293), .S0(
        n26247), .S1(n26365), .ZN(n24289) );
  MUX41 U8867 ( .I0(ram[6205]), .I1(ram[6197]), .I2(ram[6189]), .I3(
        ram[6181]), .S0(n27235), .S1(n26760), .ZN(n24291) );
  MUX41 U8868 ( .I0(ram[6173]), .I1(ram[6165]), .I2(ram[6157]), .I3(
        ram[6149]), .S0(n27235), .S1(n26760), .ZN(n24293) );
  MUX41 U8869 ( .I0(ram[6269]), .I1(ram[6261]), .I2(ram[6253]), .I3(
        ram[6245]), .S0(n27235), .S1(n26760), .ZN(n24290) );
  MUX41 U8870 ( .I0(n24310), .I1(n24311), .I2(n24312), .I3(n24313), .S0(
        n26247), .S1(n26365), .ZN(n24309) );
  MUX41 U8871 ( .I0(ram[6685]), .I1(ram[6677]), .I2(ram[6669]), .I3(
        ram[6661]), .S0(n27236), .S1(n26761), .ZN(n24313) );
  MUX41 U8872 ( .I0(ram[6717]), .I1(ram[6709]), .I2(ram[6701]), .I3(
        ram[6693]), .S0(n27236), .S1(n26761), .ZN(n24311) );
  MUX41 U8873 ( .I0(ram[6781]), .I1(ram[6773]), .I2(ram[6765]), .I3(
        ram[6757]), .S0(n27237), .S1(n26762), .ZN(n24310) );
  MUX41 U8874 ( .I0(n24265), .I1(n24266), .I2(n24267), .I3(n24268), .S0(
        n26246), .S1(n26364), .ZN(n24264) );
  MUX41 U8875 ( .I0(ram[5693]), .I1(ram[5685]), .I2(ram[5677]), .I3(
        ram[5669]), .S0(n27234), .S1(n26759), .ZN(n24266) );
  MUX41 U8876 ( .I0(ram[5661]), .I1(ram[5653]), .I2(ram[5645]), .I3(
        ram[5637]), .S0(n27234), .S1(n26759), .ZN(n24268) );
  MUX41 U8877 ( .I0(ram[5757]), .I1(ram[5749]), .I2(ram[5741]), .I3(
        ram[5733]), .S0(n27234), .S1(n26759), .ZN(n24265) );
  MUX41 U8878 ( .I0(n24521), .I1(n24522), .I2(n24523), .I3(n24524), .S0(
        n26250), .S1(n26368), .ZN(n24520) );
  MUX41 U8879 ( .I0(ram[11837]), .I1(ram[11829]), .I2(ram[11821]), .I3(
        ram[11813]), .S0(n27249), .S1(n26774), .ZN(n24522) );
  MUX41 U8880 ( .I0(ram[11805]), .I1(ram[11797]), .I2(ram[11789]), .I3(
        ram[11781]), .S0(n27249), .S1(n26774), .ZN(n24524) );
  MUX41 U8881 ( .I0(ram[11901]), .I1(ram[11893]), .I2(ram[11885]), .I3(
        ram[11877]), .S0(n27249), .S1(n26774), .ZN(n24521) );
  MUX41 U8882 ( .I0(n24461), .I1(n24462), .I2(n24463), .I3(n24464), .S0(
        n26249), .S1(n26367), .ZN(n24460) );
  MUX41 U8883 ( .I0(ram[10301]), .I1(ram[10293]), .I2(ram[10285]), .I3(
        ram[10277]), .S0(n27245), .S1(n26770), .ZN(n24462) );
  MUX41 U8884 ( .I0(ram[10269]), .I1(ram[10261]), .I2(ram[10253]), .I3(
        ram[10245]), .S0(n27245), .S1(n26770), .ZN(n24464) );
  MUX41 U8885 ( .I0(ram[10365]), .I1(ram[10357]), .I2(ram[10349]), .I3(
        ram[10341]), .S0(n27245), .S1(n26770), .ZN(n24461) );
  MUX41 U8886 ( .I0(n24436), .I1(n24437), .I2(n24438), .I3(n24439), .S0(
        n26249), .S1(n26367), .ZN(n24435) );
  MUX41 U8887 ( .I0(ram[9789]), .I1(ram[9781]), .I2(ram[9773]), .I3(
        ram[9765]), .S0(n27244), .S1(n26769), .ZN(n24437) );
  MUX41 U8888 ( .I0(ram[9757]), .I1(ram[9749]), .I2(ram[9741]), .I3(
        ram[9733]), .S0(n27244), .S1(n26769), .ZN(n24439) );
  MUX41 U8889 ( .I0(ram[9853]), .I1(ram[9845]), .I2(ram[9837]), .I3(
        ram[9829]), .S0(n27244), .S1(n26769), .ZN(n24436) );
  MUX41 U8890 ( .I0(n24376), .I1(n24377), .I2(n24378), .I3(n24379), .S0(
        n26248), .S1(n26366), .ZN(n24375) );
  MUX41 U8891 ( .I0(ram[8253]), .I1(ram[8245]), .I2(ram[8237]), .I3(
        ram[8229]), .S0(n27240), .S1(n26765), .ZN(n24377) );
  MUX41 U8892 ( .I0(ram[8221]), .I1(ram[8213]), .I2(ram[8205]), .I3(
        ram[8197]), .S0(n27240), .S1(n26765), .ZN(n24379) );
  MUX41 U8893 ( .I0(ram[8317]), .I1(ram[8309]), .I2(ram[8301]), .I3(
        ram[8293]), .S0(n27240), .S1(n26765), .ZN(n24376) );
  MUX41 U8894 ( .I0(n25376), .I1(n25377), .I2(n25378), .I3(n25379), .S0(
        n26262), .S1(n26380), .ZN(n25375) );
  MUX41 U8895 ( .I0(ram[15934]), .I1(ram[15926]), .I2(ram[15918]), .I3(
        ram[15910]), .S0(n27298), .S1(n26823), .ZN(n25377) );
  MUX41 U8896 ( .I0(ram[15902]), .I1(ram[15894]), .I2(ram[15886]), .I3(
        ram[15878]), .S0(n27298), .S1(n26823), .ZN(n25379) );
  MUX41 U8897 ( .I0(ram[15998]), .I1(ram[15990]), .I2(ram[15982]), .I3(
        ram[15974]), .S0(n27298), .S1(n26823), .ZN(n25376) );
  MUX41 U8898 ( .I0(n25336), .I1(n25337), .I2(n25338), .I3(n25339), .S0(
        n26262), .S1(n26380), .ZN(n25335) );
  MUX41 U8899 ( .I0(ram[14878]), .I1(ram[14870]), .I2(ram[14862]), .I3(
        ram[14854]), .S0(n27295), .S1(n26820), .ZN(n25339) );
  MUX41 U8900 ( .I0(ram[14910]), .I1(ram[14902]), .I2(ram[14894]), .I3(
        ram[14886]), .S0(n27296), .S1(n26821), .ZN(n25337) );
  MUX41 U8901 ( .I0(ram[14974]), .I1(ram[14966]), .I2(ram[14958]), .I3(
        ram[14950]), .S0(n27296), .S1(n26821), .ZN(n25336) );
  MUX41 U8902 ( .I0(n25316), .I1(n25317), .I2(n25318), .I3(n25319), .S0(
        n26261), .S1(n26379), .ZN(n25315) );
  MUX41 U8903 ( .I0(ram[14366]), .I1(ram[14358]), .I2(ram[14350]), .I3(
        ram[14342]), .S0(n27294), .S1(n26819), .ZN(n25319) );
  MUX41 U8904 ( .I0(ram[14398]), .I1(ram[14390]), .I2(ram[14382]), .I3(
        ram[14374]), .S0(n27294), .S1(n26819), .ZN(n25317) );
  MUX41 U8905 ( .I0(ram[14462]), .I1(ram[14454]), .I2(ram[14446]), .I3(
        ram[14438]), .S0(n27294), .S1(n26819), .ZN(n25316) );
  MUX41 U8906 ( .I0(n25291), .I1(n25292), .I2(n25293), .I3(n25294), .S0(
        n26261), .S1(n26379), .ZN(n25290) );
  MUX41 U8907 ( .I0(ram[13854]), .I1(ram[13846]), .I2(ram[13838]), .I3(
        ram[13830]), .S0(n27293), .S1(n26818), .ZN(n25294) );
  MUX41 U8908 ( .I0(ram[13886]), .I1(ram[13878]), .I2(ram[13870]), .I3(
        ram[13862]), .S0(n27293), .S1(n26818), .ZN(n25292) );
  MUX41 U8909 ( .I0(ram[13950]), .I1(ram[13942]), .I2(ram[13934]), .I3(
        ram[13926]), .S0(n27293), .S1(n26818), .ZN(n25291) );
  MUX41 U8910 ( .I0(n25251), .I1(n25252), .I2(n25253), .I3(n25254), .S0(
        n26261), .S1(n26379), .ZN(n25250) );
  MUX41 U8911 ( .I0(ram[12830]), .I1(ram[12822]), .I2(ram[12814]), .I3(
        ram[12806]), .S0(n27291), .S1(n26816), .ZN(n25254) );
  MUX41 U8912 ( .I0(ram[12862]), .I1(ram[12854]), .I2(ram[12846]), .I3(
        ram[12838]), .S0(n27291), .S1(n26816), .ZN(n25252) );
  MUX41 U8913 ( .I0(ram[12926]), .I1(ram[12918]), .I2(ram[12910]), .I3(
        ram[12902]), .S0(n27291), .S1(n26816), .ZN(n25251) );
  MUX41 U8914 ( .I0(n25231), .I1(n25232), .I2(n25233), .I3(n25234), .S0(
        n26260), .S1(n26378), .ZN(n25230) );
  MUX41 U8915 ( .I0(ram[12318]), .I1(ram[12310]), .I2(ram[12302]), .I3(
        ram[12294]), .S0(n27289), .S1(n26814), .ZN(n25234) );
  MUX41 U8916 ( .I0(ram[12350]), .I1(ram[12342]), .I2(ram[12334]), .I3(
        ram[12326]), .S0(n27289), .S1(n26814), .ZN(n25232) );
  MUX41 U8917 ( .I0(ram[12414]), .I1(ram[12406]), .I2(ram[12398]), .I3(
        ram[12390]), .S0(n27290), .S1(n26815), .ZN(n25231) );
  MUX41 U8918 ( .I0(n25034), .I1(n25035), .I2(n25036), .I3(n25037), .S0(
        n26257), .S1(n26375), .ZN(n25033) );
  MUX41 U8919 ( .I0(ram[7742]), .I1(ram[7734]), .I2(ram[7726]), .I3(
        ram[7718]), .S0(n27278), .S1(n26803), .ZN(n25035) );
  MUX41 U8920 ( .I0(ram[7710]), .I1(ram[7702]), .I2(ram[7694]), .I3(
        ram[7686]), .S0(n27278), .S1(n26803), .ZN(n25037) );
  MUX41 U8921 ( .I0(ram[7806]), .I1(ram[7798]), .I2(ram[7790]), .I3(
        ram[7782]), .S0(n27278), .S1(n26803), .ZN(n25034) );
  MUX41 U8922 ( .I0(n24974), .I1(n24975), .I2(n24976), .I3(n24977), .S0(
        n26257), .S1(n26375), .ZN(n24973) );
  MUX41 U8923 ( .I0(ram[6206]), .I1(ram[6198]), .I2(ram[6190]), .I3(
        ram[6182]), .S0(n27275), .S1(n26800), .ZN(n24975) );
  MUX41 U8924 ( .I0(ram[6174]), .I1(ram[6166]), .I2(ram[6158]), .I3(
        ram[6150]), .S0(n27275), .S1(n26800), .ZN(n24977) );
  MUX41 U8925 ( .I0(ram[6270]), .I1(ram[6262]), .I2(ram[6254]), .I3(
        ram[6246]), .S0(n27275), .S1(n26800), .ZN(n24974) );
  MUX41 U8926 ( .I0(n24994), .I1(n24995), .I2(n24996), .I3(n24997), .S0(
        n26257), .S1(n26375), .ZN(n24993) );
  MUX41 U8927 ( .I0(ram[6686]), .I1(ram[6678]), .I2(ram[6670]), .I3(
        ram[6662]), .S0(n27276), .S1(n26801), .ZN(n24997) );
  MUX41 U8928 ( .I0(ram[6718]), .I1(ram[6710]), .I2(ram[6702]), .I3(
        ram[6694]), .S0(n27276), .S1(n26801), .ZN(n24995) );
  MUX41 U8929 ( .I0(ram[6782]), .I1(ram[6774]), .I2(ram[6766]), .I3(
        ram[6758]), .S0(n27276), .S1(n26801), .ZN(n24994) );
  MUX41 U8930 ( .I0(n24949), .I1(n24950), .I2(n24951), .I3(n24952), .S0(
        n26256), .S1(n26374), .ZN(n24948) );
  MUX41 U8931 ( .I0(ram[5694]), .I1(ram[5686]), .I2(ram[5678]), .I3(
        ram[5670]), .S0(n27273), .S1(n26798), .ZN(n24950) );
  MUX41 U8932 ( .I0(ram[5662]), .I1(ram[5654]), .I2(ram[5646]), .I3(
        ram[5638]), .S0(n27273), .S1(n26798), .ZN(n24952) );
  MUX41 U8933 ( .I0(ram[5758]), .I1(ram[5750]), .I2(ram[5742]), .I3(
        ram[5734]), .S0(n27274), .S1(n26799), .ZN(n24949) );
  MUX41 U8934 ( .I0(n25205), .I1(n25206), .I2(n25207), .I3(n25208), .S0(
        n26260), .S1(n26378), .ZN(n25204) );
  MUX41 U8935 ( .I0(ram[11838]), .I1(ram[11830]), .I2(ram[11822]), .I3(
        ram[11814]), .S0(n27288), .S1(n26813), .ZN(n25206) );
  MUX41 U8936 ( .I0(ram[11806]), .I1(ram[11798]), .I2(ram[11790]), .I3(
        ram[11782]), .S0(n27288), .S1(n26813), .ZN(n25208) );
  MUX41 U8937 ( .I0(ram[11902]), .I1(ram[11894]), .I2(ram[11886]), .I3(
        ram[11878]), .S0(n27288), .S1(n26813), .ZN(n25205) );
  MUX41 U8938 ( .I0(n25145), .I1(n25146), .I2(n25147), .I3(n25148), .S0(
        n26259), .S1(n26377), .ZN(n25144) );
  MUX41 U8939 ( .I0(ram[10302]), .I1(ram[10294]), .I2(ram[10286]), .I3(
        ram[10278]), .S0(n27284), .S1(n26809), .ZN(n25146) );
  MUX41 U8940 ( .I0(ram[10270]), .I1(ram[10262]), .I2(ram[10254]), .I3(
        ram[10246]), .S0(n27284), .S1(n26809), .ZN(n25148) );
  MUX41 U8941 ( .I0(ram[10366]), .I1(ram[10358]), .I2(ram[10350]), .I3(
        ram[10342]), .S0(n27285), .S1(n26810), .ZN(n25145) );
  MUX41 U8942 ( .I0(n25120), .I1(n25121), .I2(n25122), .I3(n25123), .S0(
        n26259), .S1(n26377), .ZN(n25119) );
  MUX41 U8943 ( .I0(ram[9790]), .I1(ram[9782]), .I2(ram[9774]), .I3(
        ram[9766]), .S0(n27283), .S1(n26808), .ZN(n25121) );
  MUX41 U8944 ( .I0(ram[9758]), .I1(ram[9750]), .I2(ram[9742]), .I3(
        ram[9734]), .S0(n27283), .S1(n26808), .ZN(n25123) );
  MUX41 U8945 ( .I0(ram[9854]), .I1(ram[9846]), .I2(ram[9838]), .I3(
        ram[9830]), .S0(n27283), .S1(n26808), .ZN(n25120) );
  MUX41 U8946 ( .I0(n25060), .I1(n25061), .I2(n25062), .I3(n25063), .S0(
        n26258), .S1(n26376), .ZN(n25059) );
  MUX41 U8947 ( .I0(ram[8254]), .I1(ram[8246]), .I2(ram[8238]), .I3(
        ram[8230]), .S0(n27280), .S1(n26805), .ZN(n25061) );
  MUX41 U8948 ( .I0(ram[8222]), .I1(ram[8214]), .I2(ram[8206]), .I3(
        ram[8198]), .S0(n27279), .S1(n26804), .ZN(n25063) );
  MUX41 U8949 ( .I0(ram[8318]), .I1(ram[8310]), .I2(ram[8302]), .I3(
        ram[8294]), .S0(n27280), .S1(n26805), .ZN(n25060) );
  MUX41 U8950 ( .I0(n26060), .I1(n26061), .I2(n26062), .I3(n26063), .S0(
        n26272), .S1(n26390), .ZN(n26059) );
  MUX41 U8951 ( .I0(ram[15935]), .I1(ram[15927]), .I2(ram[15919]), .I3(
        ram[15911]), .S0(n27337), .S1(n26862), .ZN(n26061) );
  MUX41 U8952 ( .I0(ram[15903]), .I1(ram[15895]), .I2(ram[15887]), .I3(
        ram[15879]), .S0(n27337), .S1(n26862), .ZN(n26063) );
  MUX41 U8953 ( .I0(ram[15999]), .I1(ram[15991]), .I2(ram[15983]), .I3(
        ram[15975]), .S0(n27338), .S1(n26863), .ZN(n26060) );
  MUX41 U8954 ( .I0(n26020), .I1(n26021), .I2(n26022), .I3(n26023), .S0(
        n26272), .S1(n26390), .ZN(n26019) );
  MUX41 U8955 ( .I0(ram[14879]), .I1(ram[14871]), .I2(ram[14863]), .I3(
        ram[14855]), .S0(n27335), .S1(n26860), .ZN(n26023) );
  MUX41 U8956 ( .I0(ram[14911]), .I1(ram[14903]), .I2(ram[14895]), .I3(
        ram[14887]), .S0(n27335), .S1(n26860), .ZN(n26021) );
  MUX41 U8957 ( .I0(ram[14975]), .I1(ram[14967]), .I2(ram[14959]), .I3(
        ram[14951]), .S0(n27335), .S1(n26860), .ZN(n26020) );
  MUX41 U8958 ( .I0(n26000), .I1(n26001), .I2(n26002), .I3(n26003), .S0(
        n26271), .S1(n26389), .ZN(n25999) );
  MUX41 U8959 ( .I0(ram[14367]), .I1(ram[14359]), .I2(ram[14351]), .I3(
        ram[14343]), .S0(n27334), .S1(n26859), .ZN(n26003) );
  MUX41 U8960 ( .I0(ram[14399]), .I1(ram[14391]), .I2(ram[14383]), .I3(
        ram[14375]), .S0(n27334), .S1(n26859), .ZN(n26001) );
  MUX41 U8961 ( .I0(ram[14463]), .I1(ram[14455]), .I2(ram[14447]), .I3(
        ram[14439]), .S0(n27334), .S1(n26859), .ZN(n26000) );
  MUX41 U8962 ( .I0(n25975), .I1(n25976), .I2(n25977), .I3(n25978), .S0(
        n26271), .S1(n26389), .ZN(n25974) );
  MUX41 U8963 ( .I0(ram[13855]), .I1(ram[13847]), .I2(ram[13839]), .I3(
        ram[13831]), .S0(n27332), .S1(n26857), .ZN(n25978) );
  MUX41 U8964 ( .I0(ram[13887]), .I1(ram[13879]), .I2(ram[13871]), .I3(
        ram[13863]), .S0(n27332), .S1(n26857), .ZN(n25976) );
  MUX41 U8965 ( .I0(ram[13951]), .I1(ram[13943]), .I2(ram[13935]), .I3(
        ram[13927]), .S0(n27333), .S1(n26858), .ZN(n25975) );
  MUX41 U8966 ( .I0(n25935), .I1(n25936), .I2(n25937), .I3(n25938), .S0(
        n26270), .S1(n26388), .ZN(n25934) );
  MUX41 U8967 ( .I0(ram[12831]), .I1(ram[12823]), .I2(ram[12815]), .I3(
        ram[12807]), .S0(n27330), .S1(n26855), .ZN(n25938) );
  MUX41 U8968 ( .I0(ram[12863]), .I1(ram[12855]), .I2(ram[12847]), .I3(
        ram[12839]), .S0(n27330), .S1(n26855), .ZN(n25936) );
  MUX41 U8969 ( .I0(ram[12927]), .I1(ram[12919]), .I2(ram[12911]), .I3(
        ram[12903]), .S0(n27330), .S1(n26855), .ZN(n25935) );
  MUX41 U8970 ( .I0(n25915), .I1(n25916), .I2(n25917), .I3(n25918), .S0(
        n26270), .S1(n26388), .ZN(n25914) );
  MUX41 U8971 ( .I0(ram[12319]), .I1(ram[12311]), .I2(ram[12303]), .I3(
        ram[12295]), .S0(n27329), .S1(n26854), .ZN(n25918) );
  MUX41 U8972 ( .I0(ram[12351]), .I1(ram[12343]), .I2(ram[12335]), .I3(
        ram[12327]), .S0(n27329), .S1(n26854), .ZN(n25916) );
  MUX41 U8973 ( .I0(ram[12415]), .I1(ram[12407]), .I2(ram[12399]), .I3(
        ram[12391]), .S0(n27329), .S1(n26854), .ZN(n25915) );
  MUX41 U8974 ( .I0(n25718), .I1(n25719), .I2(n25720), .I3(n25721), .S0(
        n26267), .S1(n26385), .ZN(n25717) );
  MUX41 U8975 ( .I0(ram[7743]), .I1(ram[7735]), .I2(ram[7727]), .I3(
        ram[7719]), .S0(n27318), .S1(n26843), .ZN(n25719) );
  MUX41 U8976 ( .I0(ram[7711]), .I1(ram[7703]), .I2(ram[7695]), .I3(
        ram[7687]), .S0(n27318), .S1(n26843), .ZN(n25721) );
  MUX41 U8977 ( .I0(ram[7807]), .I1(ram[7799]), .I2(ram[7791]), .I3(
        ram[7783]), .S0(n27318), .S1(n26843), .ZN(n25718) );
  MUX41 U8978 ( .I0(n25658), .I1(n25659), .I2(n25660), .I3(n25661), .S0(
        n26266), .S1(n26384), .ZN(n25657) );
  MUX41 U8979 ( .I0(ram[6207]), .I1(ram[6199]), .I2(ram[6191]), .I3(
        ram[6183]), .S0(n27314), .S1(n26839), .ZN(n25659) );
  MUX41 U8980 ( .I0(ram[6175]), .I1(ram[6167]), .I2(ram[6159]), .I3(
        ram[6151]), .S0(n27314), .S1(n26839), .ZN(n25661) );
  MUX41 U8981 ( .I0(ram[6271]), .I1(ram[6263]), .I2(ram[6255]), .I3(
        ram[6247]), .S0(n27314), .S1(n26839), .ZN(n25658) );
  MUX41 U8982 ( .I0(n25678), .I1(n25679), .I2(n25680), .I3(n25681), .S0(
        n26267), .S1(n26385), .ZN(n25677) );
  MUX41 U8983 ( .I0(ram[6687]), .I1(ram[6679]), .I2(ram[6671]), .I3(
        ram[6663]), .S0(n27315), .S1(n26840), .ZN(n25681) );
  MUX41 U8984 ( .I0(ram[6719]), .I1(ram[6711]), .I2(ram[6703]), .I3(
        ram[6695]), .S0(n27315), .S1(n26840), .ZN(n25679) );
  MUX41 U8985 ( .I0(ram[6783]), .I1(ram[6775]), .I2(ram[6767]), .I3(
        ram[6759]), .S0(n27315), .S1(n26840), .ZN(n25678) );
  MUX41 U8986 ( .I0(n25633), .I1(n25634), .I2(n25635), .I3(n25636), .S0(
        n26266), .S1(n26384), .ZN(n25632) );
  MUX41 U8987 ( .I0(ram[5695]), .I1(ram[5687]), .I2(ram[5679]), .I3(
        ram[5671]), .S0(n27313), .S1(n26838), .ZN(n25634) );
  MUX41 U8988 ( .I0(ram[5663]), .I1(ram[5655]), .I2(ram[5647]), .I3(
        ram[5639]), .S0(n27313), .S1(n26838), .ZN(n25636) );
  MUX41 U8989 ( .I0(ram[5759]), .I1(ram[5751]), .I2(ram[5743]), .I3(
        ram[5735]), .S0(n27313), .S1(n26838), .ZN(n25633) );
  MUX41 U8990 ( .I0(n25889), .I1(n25890), .I2(n25891), .I3(n25892), .S0(
        n26270), .S1(n26388), .ZN(n25888) );
  MUX41 U8991 ( .I0(ram[11839]), .I1(ram[11831]), .I2(ram[11823]), .I3(
        ram[11815]), .S0(n27328), .S1(n26853), .ZN(n25890) );
  MUX41 U8992 ( .I0(ram[11807]), .I1(ram[11799]), .I2(ram[11791]), .I3(
        ram[11783]), .S0(n27327), .S1(n26852), .ZN(n25892) );
  MUX41 U8993 ( .I0(ram[11903]), .I1(ram[11895]), .I2(ram[11887]), .I3(
        ram[11879]), .S0(n27328), .S1(n26853), .ZN(n25889) );
  MUX41 U8994 ( .I0(n25829), .I1(n25830), .I2(n25831), .I3(n25832), .S0(
        n26269), .S1(n26387), .ZN(n25828) );
  MUX41 U8995 ( .I0(ram[10303]), .I1(ram[10295]), .I2(ram[10287]), .I3(
        ram[10279]), .S0(n27324), .S1(n26849), .ZN(n25830) );
  MUX41 U8996 ( .I0(ram[10271]), .I1(ram[10263]), .I2(ram[10255]), .I3(
        ram[10247]), .S0(n27324), .S1(n26849), .ZN(n25832) );
  MUX41 U8997 ( .I0(ram[10367]), .I1(ram[10359]), .I2(ram[10351]), .I3(
        ram[10343]), .S0(n27324), .S1(n26849), .ZN(n25829) );
  MUX41 U8998 ( .I0(n25804), .I1(n25805), .I2(n25806), .I3(n25807), .S0(
        n26269), .S1(n26387), .ZN(n25803) );
  MUX41 U8999 ( .I0(ram[9791]), .I1(ram[9783]), .I2(ram[9775]), .I3(
        ram[9767]), .S0(n27323), .S1(n26848), .ZN(n25805) );
  MUX41 U9000 ( .I0(ram[9759]), .I1(ram[9751]), .I2(ram[9743]), .I3(
        ram[9735]), .S0(n27323), .S1(n26848), .ZN(n25807) );
  MUX41 U9001 ( .I0(ram[9855]), .I1(ram[9847]), .I2(ram[9839]), .I3(
        ram[9831]), .S0(n27323), .S1(n26848), .ZN(n25804) );
  MUX41 U9002 ( .I0(n25744), .I1(n25745), .I2(n25746), .I3(n25747), .S0(
        n26268), .S1(n26386), .ZN(n25743) );
  MUX41 U9003 ( .I0(ram[8255]), .I1(ram[8247]), .I2(ram[8239]), .I3(
        ram[8231]), .S0(n27319), .S1(n26844), .ZN(n25745) );
  MUX41 U9004 ( .I0(ram[8223]), .I1(ram[8215]), .I2(ram[8207]), .I3(
        ram[8199]), .S0(n27319), .S1(n26844), .ZN(n25747) );
  MUX41 U9005 ( .I0(ram[8319]), .I1(ram[8311]), .I2(ram[8303]), .I3(
        ram[8295]), .S0(n27319), .S1(n26844), .ZN(n25744) );
  MUX41 U9006 ( .I0(ram[3512]), .I1(ram[3504]), .I2(ram[3496]), .I3(
        ram[3488]), .S0(n27032), .S1(n26557), .ZN(n20755) );
  MUX41 U9007 ( .I0(ram[3256]), .I1(ram[3248]), .I2(ram[3240]), .I3(
        ram[3232]), .S0(n27031), .S1(n26556), .ZN(n20745) );
  MUX41 U9008 ( .I0(ram[3128]), .I1(ram[3120]), .I2(ram[3112]), .I3(
        ram[3104]), .S0(n27031), .S1(n26556), .ZN(n20740) );
  MUX41 U9009 ( .I0(ram[1464]), .I1(ram[1456]), .I2(ram[1448]), .I3(
        ram[1440]), .S0(n27027), .S1(n26552), .ZN(n20670) );
  MUX41 U9010 ( .I0(ram[1208]), .I1(ram[1200]), .I2(ram[1192]), .I3(
        ram[1184]), .S0(n27026), .S1(n26551), .ZN(n20660) );
  MUX41 U9011 ( .I0(ram[3513]), .I1(ram[3505]), .I2(ram[3497]), .I3(
        ram[3489]), .S0(n27071), .S1(n26596), .ZN(n21439) );
  MUX41 U9012 ( .I0(ram[3257]), .I1(ram[3249]), .I2(ram[3241]), .I3(
        ram[3233]), .S0(n27071), .S1(n26596), .ZN(n21429) );
  MUX41 U9013 ( .I0(ram[3129]), .I1(ram[3121]), .I2(ram[3113]), .I3(
        ram[3105]), .S0(n27070), .S1(n26595), .ZN(n21424) );
  MUX41 U9014 ( .I0(ram[1465]), .I1(ram[1457]), .I2(ram[1449]), .I3(
        ram[1441]), .S0(n27066), .S1(n26591), .ZN(n21354) );
  MUX41 U9015 ( .I0(ram[1209]), .I1(ram[1201]), .I2(ram[1193]), .I3(
        ram[1185]), .S0(n27066), .S1(n26591), .ZN(n21344) );
  MUX41 U9016 ( .I0(ram[3514]), .I1(ram[3506]), .I2(ram[3498]), .I3(
        ram[3490]), .S0(n27111), .S1(n26636), .ZN(n22123) );
  MUX41 U9017 ( .I0(ram[3258]), .I1(ram[3250]), .I2(ram[3242]), .I3(
        ram[3234]), .S0(n27110), .S1(n26635), .ZN(n22113) );
  MUX41 U9018 ( .I0(ram[3130]), .I1(ram[3122]), .I2(ram[3114]), .I3(
        ram[3106]), .S0(n27110), .S1(n26635), .ZN(n22108) );
  MUX41 U9019 ( .I0(ram[1466]), .I1(ram[1458]), .I2(ram[1450]), .I3(
        ram[1442]), .S0(n27106), .S1(n26631), .ZN(n22038) );
  MUX41 U9020 ( .I0(ram[1210]), .I1(ram[1202]), .I2(ram[1194]), .I3(
        ram[1186]), .S0(n27105), .S1(n26630), .ZN(n22028) );
  MUX41 U9021 ( .I0(ram[1082]), .I1(ram[1074]), .I2(ram[1066]), .I3(
        ram[1058]), .S0(n27105), .S1(n26630), .ZN(n22023) );
  MUX41 U9022 ( .I0(ram[3515]), .I1(ram[3507]), .I2(ram[3499]), .I3(
        ram[3491]), .S0(n27150), .S1(n26675), .ZN(n22807) );
  MUX41 U9023 ( .I0(ram[3259]), .I1(ram[3251]), .I2(ram[3243]), .I3(
        ram[3235]), .S0(n27149), .S1(n26674), .ZN(n22797) );
  MUX41 U9024 ( .I0(ram[3131]), .I1(ram[3123]), .I2(ram[3115]), .I3(
        ram[3107]), .S0(n27149), .S1(n26674), .ZN(n22792) );
  MUX41 U9025 ( .I0(ram[1467]), .I1(ram[1459]), .I2(ram[1451]), .I3(
        ram[1443]), .S0(n27145), .S1(n26670), .ZN(n22722) );
  MUX41 U9026 ( .I0(ram[1211]), .I1(ram[1203]), .I2(ram[1195]), .I3(
        ram[1187]), .S0(n27144), .S1(n26669), .ZN(n22712) );
  MUX41 U9027 ( .I0(ram[1083]), .I1(ram[1075]), .I2(ram[1067]), .I3(
        ram[1059]), .S0(n27144), .S1(n26669), .ZN(n22707) );
  MUX41 U9028 ( .I0(ram[3516]), .I1(ram[3508]), .I2(ram[3500]), .I3(
        ram[3492]), .S0(n27189), .S1(n26714), .ZN(n23491) );
  MUX41 U9029 ( .I0(ram[3260]), .I1(ram[3252]), .I2(ram[3244]), .I3(
        ram[3236]), .S0(n27189), .S1(n26714), .ZN(n23481) );
  MUX41 U9030 ( .I0(ram[3132]), .I1(ram[3124]), .I2(ram[3116]), .I3(
        ram[3108]), .S0(n27188), .S1(n26713), .ZN(n23476) );
  MUX41 U9031 ( .I0(ram[1468]), .I1(ram[1460]), .I2(ram[1452]), .I3(
        ram[1444]), .S0(n27184), .S1(n26709), .ZN(n23406) );
  MUX41 U9032 ( .I0(ram[1212]), .I1(ram[1204]), .I2(ram[1196]), .I3(
        ram[1188]), .S0(n27184), .S1(n26709), .ZN(n23396) );
  MUX41 U9033 ( .I0(ram[1084]), .I1(ram[1076]), .I2(ram[1068]), .I3(
        ram[1060]), .S0(n27184), .S1(n26709), .ZN(n23391) );
  MUX41 U9034 ( .I0(ram[3517]), .I1(ram[3509]), .I2(ram[3501]), .I3(
        ram[3493]), .S0(n27229), .S1(n26754), .ZN(n24175) );
  MUX41 U9035 ( .I0(ram[3261]), .I1(ram[3253]), .I2(ram[3245]), .I3(
        ram[3237]), .S0(n27228), .S1(n26753), .ZN(n24165) );
  MUX41 U9036 ( .I0(ram[3133]), .I1(ram[3125]), .I2(ram[3117]), .I3(
        ram[3109]), .S0(n27228), .S1(n26753), .ZN(n24160) );
  MUX41 U9037 ( .I0(ram[1469]), .I1(ram[1461]), .I2(ram[1453]), .I3(
        ram[1445]), .S0(n27224), .S1(n26749), .ZN(n24090) );
  MUX41 U9038 ( .I0(ram[1213]), .I1(ram[1205]), .I2(ram[1197]), .I3(
        ram[1189]), .S0(n27223), .S1(n26748), .ZN(n24080) );
  MUX41 U9039 ( .I0(ram[1085]), .I1(ram[1077]), .I2(ram[1069]), .I3(
        ram[1061]), .S0(n27223), .S1(n26748), .ZN(n24075) );
  MUX41 U9040 ( .I0(ram[3518]), .I1(ram[3510]), .I2(ram[3502]), .I3(
        ram[3494]), .S0(n27268), .S1(n26793), .ZN(n24859) );
  MUX41 U9041 ( .I0(ram[3262]), .I1(ram[3254]), .I2(ram[3246]), .I3(
        ram[3238]), .S0(n27268), .S1(n26793), .ZN(n24849) );
  MUX41 U9042 ( .I0(ram[3134]), .I1(ram[3126]), .I2(ram[3118]), .I3(
        ram[3110]), .S0(n27267), .S1(n26792), .ZN(n24844) );
  MUX41 U9043 ( .I0(ram[1470]), .I1(ram[1462]), .I2(ram[1454]), .I3(
        ram[1446]), .S0(n27263), .S1(n26788), .ZN(n24774) );
  MUX41 U9044 ( .I0(ram[1214]), .I1(ram[1206]), .I2(ram[1198]), .I3(
        ram[1190]), .S0(n27263), .S1(n26788), .ZN(n24764) );
  MUX41 U9045 ( .I0(ram[1086]), .I1(ram[1078]), .I2(ram[1070]), .I3(
        ram[1062]), .S0(n27262), .S1(n26787), .ZN(n24759) );
  MUX41 U9046 ( .I0(ram[3519]), .I1(ram[3511]), .I2(ram[3503]), .I3(
        ram[3495]), .S0(n27308), .S1(n26833), .ZN(n25543) );
  MUX41 U9047 ( .I0(ram[3263]), .I1(ram[3255]), .I2(ram[3247]), .I3(
        ram[3239]), .S0(n27307), .S1(n26832), .ZN(n25533) );
  MUX41 U9048 ( .I0(ram[3135]), .I1(ram[3127]), .I2(ram[3119]), .I3(
        ram[3111]), .S0(n27307), .S1(n26832), .ZN(n25528) );
  MUX41 U9049 ( .I0(ram[1471]), .I1(ram[1463]), .I2(ram[1455]), .I3(
        ram[1447]), .S0(n27303), .S1(n26828), .ZN(n25458) );
  MUX41 U9050 ( .I0(ram[1215]), .I1(ram[1207]), .I2(ram[1199]), .I3(
        ram[1191]), .S0(n27302), .S1(n26827), .ZN(n25448) );
  MUX41 U9051 ( .I0(ram[1087]), .I1(ram[1079]), .I2(ram[1071]), .I3(
        ram[1063]), .S0(n27302), .S1(n26827), .ZN(n25443) );
  MUX41 U9052 ( .I0(ram[15800]), .I1(ram[15792]), .I2(ram[15784]), .I3(
        ram[15776]), .S0(n27061), .S1(n26586), .ZN(n21268) );
  MUX41 U9053 ( .I0(ram[15544]), .I1(ram[15536]), .I2(ram[15528]), .I3(
        ram[15520]), .S0(n27061), .S1(n26586), .ZN(n21258) );
  MUX41 U9054 ( .I0(ram[15416]), .I1(ram[15408]), .I2(ram[15400]), .I3(
        ram[15392]), .S0(n27060), .S1(n26585), .ZN(n21253) );
  MUX41 U9055 ( .I0(ram[13752]), .I1(ram[13744]), .I2(ram[13736]), .I3(
        ram[13728]), .S0(n27056), .S1(n26581), .ZN(n21183) );
  MUX41 U9056 ( .I0(ram[13496]), .I1(ram[13488]), .I2(ram[13480]), .I3(
        ram[13472]), .S0(n27056), .S1(n26581), .ZN(n21173) );
  MUX41 U9057 ( .I0(ram[13368]), .I1(ram[13360]), .I2(ram[13352]), .I3(
        ram[13344]), .S0(n27056), .S1(n26581), .ZN(n21168) );
  MUX41 U9058 ( .I0(ram[7608]), .I1(ram[7600]), .I2(ram[7592]), .I3(
        ram[7584]), .S0(n27042), .S1(n26567), .ZN(n20926) );
  MUX41 U9059 ( .I0(ram[7352]), .I1(ram[7344]), .I2(ram[7336]), .I3(
        ram[7328]), .S0(n27041), .S1(n26566), .ZN(n20916) );
  MUX41 U9060 ( .I0(ram[11704]), .I1(ram[11696]), .I2(ram[11688]), .I3(
        ram[11680]), .S0(n27052), .S1(n26577), .ZN(n21097) );
  MUX41 U9061 ( .I0(ram[9656]), .I1(ram[9648]), .I2(ram[9640]), .I3(
        ram[9632]), .S0(n27047), .S1(n26572), .ZN(n21012) );
  MUX41 U9062 ( .I0(ram[15801]), .I1(ram[15793]), .I2(ram[15785]), .I3(
        ram[15777]), .S0(n27101), .S1(n26626), .ZN(n21952) );
  MUX41 U9063 ( .I0(ram[15545]), .I1(ram[15537]), .I2(ram[15529]), .I3(
        ram[15521]), .S0(n27100), .S1(n26625), .ZN(n21942) );
  MUX41 U9064 ( .I0(ram[15417]), .I1(ram[15409]), .I2(ram[15401]), .I3(
        ram[15393]), .S0(n27100), .S1(n26625), .ZN(n21937) );
  MUX41 U9065 ( .I0(ram[13753]), .I1(ram[13745]), .I2(ram[13737]), .I3(
        ram[13729]), .S0(n27096), .S1(n26621), .ZN(n21867) );
  MUX41 U9066 ( .I0(ram[13497]), .I1(ram[13489]), .I2(ram[13481]), .I3(
        ram[13473]), .S0(n27095), .S1(n26620), .ZN(n21857) );
  MUX41 U9067 ( .I0(ram[13369]), .I1(ram[13361]), .I2(ram[13353]), .I3(
        ram[13345]), .S0(n27095), .S1(n26620), .ZN(n21852) );
  MUX41 U9068 ( .I0(n21323), .I1(n21324), .I2(n21325), .I3(n21326), .S0(
        n26204), .S1(n26322), .ZN(n21322) );
  MUX41 U9069 ( .I0(ram[697]), .I1(ram[689]), .I2(ram[681]), .I3(ram[673]), .S0(n27064), .S1(n26589), .ZN(n21324) );
  MUX41 U9070 ( .I0(ram[665]), .I1(ram[657]), .I2(ram[649]), .I3(ram[641]), .S0(n27064), .S1(n26589), .ZN(n21326) );
  MUX41 U9071 ( .I0(ram[761]), .I1(ram[753]), .I2(ram[745]), .I3(ram[737]), .S0(n27065), .S1(n26590), .ZN(n21323) );
  MUX41 U9072 ( .I0(ram[7609]), .I1(ram[7601]), .I2(ram[7593]), .I3(
        ram[7585]), .S0(n27081), .S1(n26606), .ZN(n21610) );
  MUX41 U9073 ( .I0(ram[7353]), .I1(ram[7345]), .I2(ram[7337]), .I3(
        ram[7329]), .S0(n27080), .S1(n26605), .ZN(n21600) );
  MUX41 U9074 ( .I0(ram[11705]), .I1(ram[11697]), .I2(ram[11689]), .I3(
        ram[11681]), .S0(n27091), .S1(n26616), .ZN(n21781) );
  MUX41 U9075 ( .I0(ram[9657]), .I1(ram[9649]), .I2(ram[9641]), .I3(
        ram[9633]), .S0(n27086), .S1(n26611), .ZN(n21696) );
  MUX41 U9076 ( .I0(ram[15802]), .I1(ram[15794]), .I2(ram[15786]), .I3(
        ram[15778]), .S0(n27140), .S1(n26665), .ZN(n22636) );
  MUX41 U9077 ( .I0(ram[15546]), .I1(ram[15538]), .I2(ram[15530]), .I3(
        ram[15522]), .S0(n27140), .S1(n26665), .ZN(n22626) );
  MUX41 U9078 ( .I0(ram[15418]), .I1(ram[15410]), .I2(ram[15402]), .I3(
        ram[15394]), .S0(n27139), .S1(n26664), .ZN(n22621) );
  MUX41 U9079 ( .I0(ram[13754]), .I1(ram[13746]), .I2(ram[13738]), .I3(
        ram[13730]), .S0(n27135), .S1(n26660), .ZN(n22551) );
  MUX41 U9080 ( .I0(ram[13498]), .I1(ram[13490]), .I2(ram[13482]), .I3(
        ram[13474]), .S0(n27135), .S1(n26660), .ZN(n22541) );
  MUX41 U9081 ( .I0(ram[13370]), .I1(ram[13362]), .I2(ram[13354]), .I3(
        ram[13346]), .S0(n27134), .S1(n26659), .ZN(n22536) );
  MUX41 U9082 ( .I0(n22007), .I1(n22008), .I2(n22009), .I3(n22010), .S0(
        n26214), .S1(n26332), .ZN(n22006) );
  MUX41 U9083 ( .I0(ram[698]), .I1(ram[690]), .I2(ram[682]), .I3(ram[674]), .S0(n27104), .S1(n26629), .ZN(n22008) );
  MUX41 U9084 ( .I0(ram[666]), .I1(ram[658]), .I2(ram[650]), .I3(ram[642]), .S0(n27104), .S1(n26629), .ZN(n22010) );
  MUX41 U9085 ( .I0(ram[762]), .I1(ram[754]), .I2(ram[746]), .I3(ram[738]), .S0(n27104), .S1(n26629), .ZN(n22007) );
  MUX41 U9086 ( .I0(ram[7610]), .I1(ram[7602]), .I2(ram[7594]), .I3(
        ram[7586]), .S0(n27120), .S1(n26645), .ZN(n22294) );
  MUX41 U9087 ( .I0(ram[7354]), .I1(ram[7346]), .I2(ram[7338]), .I3(
        ram[7330]), .S0(n27120), .S1(n26645), .ZN(n22284) );
  MUX41 U9088 ( .I0(ram[7226]), .I1(ram[7218]), .I2(ram[7210]), .I3(
        ram[7202]), .S0(n27120), .S1(n26645), .ZN(n22279) );
  MUX41 U9089 ( .I0(ram[11706]), .I1(ram[11698]), .I2(ram[11690]), .I3(
        ram[11682]), .S0(n27130), .S1(n26655), .ZN(n22465) );
  MUX41 U9090 ( .I0(ram[11450]), .I1(ram[11442]), .I2(ram[11434]), .I3(
        ram[11426]), .S0(n27130), .S1(n26655), .ZN(n22455) );
  MUX41 U9091 ( .I0(ram[9658]), .I1(ram[9650]), .I2(ram[9642]), .I3(
        ram[9634]), .S0(n27125), .S1(n26650), .ZN(n22380) );
  MUX41 U9092 ( .I0(ram[15803]), .I1(ram[15795]), .I2(ram[15787]), .I3(
        ram[15779]), .S0(n27180), .S1(n26705), .ZN(n23320) );
  MUX41 U9093 ( .I0(ram[15547]), .I1(ram[15539]), .I2(ram[15531]), .I3(
        ram[15523]), .S0(n27179), .S1(n26704), .ZN(n23310) );
  MUX41 U9094 ( .I0(ram[15419]), .I1(ram[15411]), .I2(ram[15403]), .I3(
        ram[15395]), .S0(n27179), .S1(n26704), .ZN(n23305) );
  MUX41 U9095 ( .I0(ram[13755]), .I1(ram[13747]), .I2(ram[13739]), .I3(
        ram[13731]), .S0(n27175), .S1(n26700), .ZN(n23235) );
  MUX41 U9096 ( .I0(ram[13499]), .I1(ram[13491]), .I2(ram[13483]), .I3(
        ram[13475]), .S0(n27174), .S1(n26699), .ZN(n23225) );
  MUX41 U9097 ( .I0(ram[13371]), .I1(ram[13363]), .I2(ram[13355]), .I3(
        ram[13347]), .S0(n27174), .S1(n26699), .ZN(n23220) );
  MUX41 U9098 ( .I0(n22691), .I1(n22692), .I2(n22693), .I3(n22694), .S0(
        n26224), .S1(n26342), .ZN(n22690) );
  MUX41 U9099 ( .I0(ram[699]), .I1(ram[691]), .I2(ram[683]), .I3(ram[675]), .S0(n27143), .S1(n26668), .ZN(n22692) );
  MUX41 U9100 ( .I0(ram[667]), .I1(ram[659]), .I2(ram[651]), .I3(ram[643]), .S0(n27143), .S1(n26668), .ZN(n22694) );
  MUX41 U9101 ( .I0(ram[763]), .I1(ram[755]), .I2(ram[747]), .I3(ram[739]), .S0(n27143), .S1(n26668), .ZN(n22691) );
  MUX41 U9102 ( .I0(ram[7611]), .I1(ram[7603]), .I2(ram[7595]), .I3(
        ram[7587]), .S0(n27160), .S1(n26685), .ZN(n22978) );
  MUX41 U9103 ( .I0(ram[7355]), .I1(ram[7347]), .I2(ram[7339]), .I3(
        ram[7331]), .S0(n27159), .S1(n26684), .ZN(n22968) );
  MUX41 U9104 ( .I0(ram[7227]), .I1(ram[7219]), .I2(ram[7211]), .I3(
        ram[7203]), .S0(n27159), .S1(n26684), .ZN(n22963) );
  MUX41 U9105 ( .I0(ram[11707]), .I1(ram[11699]), .I2(ram[11691]), .I3(
        ram[11683]), .S0(n27170), .S1(n26695), .ZN(n23149) );
  MUX41 U9106 ( .I0(ram[11451]), .I1(ram[11443]), .I2(ram[11435]), .I3(
        ram[11427]), .S0(n27169), .S1(n26694), .ZN(n23139) );
  MUX41 U9107 ( .I0(ram[9659]), .I1(ram[9651]), .I2(ram[9643]), .I3(
        ram[9635]), .S0(n27165), .S1(n26690), .ZN(n23064) );
  MUX41 U9108 ( .I0(ram[15804]), .I1(ram[15796]), .I2(ram[15788]), .I3(
        ram[15780]), .S0(n27219), .S1(n26744), .ZN(n24004) );
  MUX41 U9109 ( .I0(ram[15548]), .I1(ram[15540]), .I2(ram[15532]), .I3(
        ram[15524]), .S0(n27218), .S1(n26743), .ZN(n23994) );
  MUX41 U9110 ( .I0(ram[15420]), .I1(ram[15412]), .I2(ram[15404]), .I3(
        ram[15396]), .S0(n27218), .S1(n26743), .ZN(n23989) );
  MUX41 U9111 ( .I0(ram[13756]), .I1(ram[13748]), .I2(ram[13740]), .I3(
        ram[13732]), .S0(n27214), .S1(n26739), .ZN(n23919) );
  MUX41 U9112 ( .I0(ram[13500]), .I1(ram[13492]), .I2(ram[13484]), .I3(
        ram[13476]), .S0(n27213), .S1(n26738), .ZN(n23909) );
  MUX41 U9113 ( .I0(ram[13372]), .I1(ram[13364]), .I2(ram[13356]), .I3(
        ram[13348]), .S0(n27213), .S1(n26738), .ZN(n23904) );
  MUX41 U9114 ( .I0(n23375), .I1(n23376), .I2(n23377), .I3(n23378), .S0(
        n26234), .S1(n26352), .ZN(n23374) );
  MUX41 U9115 ( .I0(ram[700]), .I1(ram[692]), .I2(ram[684]), .I3(ram[676]), .S0(n27183), .S1(n26708), .ZN(n23376) );
  MUX41 U9116 ( .I0(ram[668]), .I1(ram[660]), .I2(ram[652]), .I3(ram[644]), .S0(n27183), .S1(n26708), .ZN(n23378) );
  MUX41 U9117 ( .I0(ram[764]), .I1(ram[756]), .I2(ram[748]), .I3(ram[740]), .S0(n27183), .S1(n26708), .ZN(n23375) );
  MUX41 U9118 ( .I0(ram[7612]), .I1(ram[7604]), .I2(ram[7596]), .I3(
        ram[7588]), .S0(n27199), .S1(n26724), .ZN(n23662) );
  MUX41 U9119 ( .I0(ram[7356]), .I1(ram[7348]), .I2(ram[7340]), .I3(
        ram[7332]), .S0(n27199), .S1(n26724), .ZN(n23652) );
  MUX41 U9120 ( .I0(ram[7228]), .I1(ram[7220]), .I2(ram[7212]), .I3(
        ram[7204]), .S0(n27198), .S1(n26723), .ZN(n23647) );
  MUX41 U9121 ( .I0(ram[11708]), .I1(ram[11700]), .I2(ram[11692]), .I3(
        ram[11684]), .S0(n27209), .S1(n26734), .ZN(n23833) );
  MUX41 U9122 ( .I0(ram[11452]), .I1(ram[11444]), .I2(ram[11436]), .I3(
        ram[11428]), .S0(n27208), .S1(n26733), .ZN(n23823) );
  MUX41 U9123 ( .I0(ram[9660]), .I1(ram[9652]), .I2(ram[9644]), .I3(
        ram[9636]), .S0(n27204), .S1(n26729), .ZN(n23748) );
  MUX41 U9124 ( .I0(ram[15805]), .I1(ram[15797]), .I2(ram[15789]), .I3(
        ram[15781]), .S0(n27258), .S1(n26783), .ZN(n24688) );
  MUX41 U9125 ( .I0(ram[15549]), .I1(ram[15541]), .I2(ram[15533]), .I3(
        ram[15525]), .S0(n27258), .S1(n26783), .ZN(n24678) );
  MUX41 U9126 ( .I0(ram[15421]), .I1(ram[15413]), .I2(ram[15405]), .I3(
        ram[15397]), .S0(n27257), .S1(n26782), .ZN(n24673) );
  MUX41 U9127 ( .I0(ram[13757]), .I1(ram[13749]), .I2(ram[13741]), .I3(
        ram[13733]), .S0(n27253), .S1(n26778), .ZN(n24603) );
  MUX41 U9128 ( .I0(ram[13501]), .I1(ram[13493]), .I2(ram[13485]), .I3(
        ram[13477]), .S0(n27253), .S1(n26778), .ZN(n24593) );
  MUX41 U9129 ( .I0(ram[13373]), .I1(ram[13365]), .I2(ram[13357]), .I3(
        ram[13349]), .S0(n27252), .S1(n26777), .ZN(n24588) );
  MUX41 U9130 ( .I0(n24059), .I1(n24060), .I2(n24061), .I3(n24062), .S0(
        n26243), .S1(n26361), .ZN(n24058) );
  MUX41 U9131 ( .I0(ram[701]), .I1(ram[693]), .I2(ram[685]), .I3(ram[677]), .S0(n27222), .S1(n26747), .ZN(n24060) );
  MUX41 U9132 ( .I0(ram[669]), .I1(ram[661]), .I2(ram[653]), .I3(ram[645]), .S0(n27222), .S1(n26747), .ZN(n24062) );
  MUX41 U9133 ( .I0(ram[765]), .I1(ram[757]), .I2(ram[749]), .I3(ram[741]), .S0(n27222), .S1(n26747), .ZN(n24059) );
  MUX41 U9134 ( .I0(ram[7613]), .I1(ram[7605]), .I2(ram[7597]), .I3(
        ram[7589]), .S0(n27239), .S1(n26764), .ZN(n24346) );
  MUX41 U9135 ( .I0(ram[7357]), .I1(ram[7349]), .I2(ram[7341]), .I3(
        ram[7333]), .S0(n27238), .S1(n26763), .ZN(n24336) );
  MUX41 U9136 ( .I0(ram[7229]), .I1(ram[7221]), .I2(ram[7213]), .I3(
        ram[7205]), .S0(n27238), .S1(n26763), .ZN(n24331) );
  MUX41 U9137 ( .I0(ram[11709]), .I1(ram[11701]), .I2(ram[11693]), .I3(
        ram[11685]), .S0(n27248), .S1(n26773), .ZN(n24517) );
  MUX41 U9138 ( .I0(ram[11453]), .I1(ram[11445]), .I2(ram[11437]), .I3(
        ram[11429]), .S0(n27248), .S1(n26773), .ZN(n24507) );
  MUX41 U9139 ( .I0(ram[9661]), .I1(ram[9653]), .I2(ram[9645]), .I3(
        ram[9637]), .S0(n27244), .S1(n26769), .ZN(n24432) );
  MUX41 U9140 ( .I0(ram[15806]), .I1(ram[15798]), .I2(ram[15790]), .I3(
        ram[15782]), .S0(n27298), .S1(n26823), .ZN(n25372) );
  MUX41 U9141 ( .I0(ram[15550]), .I1(ram[15542]), .I2(ram[15534]), .I3(
        ram[15526]), .S0(n27297), .S1(n26822), .ZN(n25362) );
  MUX41 U9142 ( .I0(ram[15422]), .I1(ram[15414]), .I2(ram[15406]), .I3(
        ram[15398]), .S0(n27297), .S1(n26822), .ZN(n25357) );
  MUX41 U9143 ( .I0(ram[13758]), .I1(ram[13750]), .I2(ram[13742]), .I3(
        ram[13734]), .S0(n27293), .S1(n26818), .ZN(n25287) );
  MUX41 U9144 ( .I0(ram[13502]), .I1(ram[13494]), .I2(ram[13486]), .I3(
        ram[13478]), .S0(n27292), .S1(n26817), .ZN(n25277) );
  MUX41 U9145 ( .I0(ram[13374]), .I1(ram[13366]), .I2(ram[13358]), .I3(
        ram[13350]), .S0(n27292), .S1(n26817), .ZN(n25272) );
  MUX41 U9146 ( .I0(n24743), .I1(n24744), .I2(n24745), .I3(n24746), .S0(
        n26253), .S1(n26371), .ZN(n24742) );
  MUX41 U9147 ( .I0(ram[702]), .I1(ram[694]), .I2(ram[686]), .I3(ram[678]), .S0(n27261), .S1(n26786), .ZN(n24744) );
  MUX41 U9148 ( .I0(ram[670]), .I1(ram[662]), .I2(ram[654]), .I3(ram[646]), .S0(n27261), .S1(n26786), .ZN(n24746) );
  MUX41 U9149 ( .I0(ram[766]), .I1(ram[758]), .I2(ram[750]), .I3(ram[742]), .S0(n27262), .S1(n26787), .ZN(n24743) );
  MUX41 U9150 ( .I0(ram[7614]), .I1(ram[7606]), .I2(ram[7598]), .I3(
        ram[7590]), .S0(n27278), .S1(n26803), .ZN(n25030) );
  MUX41 U9151 ( .I0(ram[7358]), .I1(ram[7350]), .I2(ram[7342]), .I3(
        ram[7334]), .S0(n27277), .S1(n26802), .ZN(n25020) );
  MUX41 U9152 ( .I0(ram[7230]), .I1(ram[7222]), .I2(ram[7214]), .I3(
        ram[7206]), .S0(n27277), .S1(n26802), .ZN(n25015) );
  MUX41 U9153 ( .I0(ram[11710]), .I1(ram[11702]), .I2(ram[11694]), .I3(
        ram[11686]), .S0(n27288), .S1(n26813), .ZN(n25201) );
  MUX41 U9154 ( .I0(ram[11454]), .I1(ram[11446]), .I2(ram[11438]), .I3(
        ram[11430]), .S0(n27287), .S1(n26812), .ZN(n25191) );
  MUX41 U9155 ( .I0(ram[9662]), .I1(ram[9654]), .I2(ram[9646]), .I3(
        ram[9638]), .S0(n27283), .S1(n26808), .ZN(n25116) );
  MUX41 U9156 ( .I0(ram[15807]), .I1(ram[15799]), .I2(ram[15791]), .I3(
        ram[15783]), .S0(n27337), .S1(n26862), .ZN(n26056) );
  MUX41 U9157 ( .I0(ram[15551]), .I1(ram[15543]), .I2(ram[15535]), .I3(
        ram[15527]), .S0(n27336), .S1(n26861), .ZN(n26046) );
  MUX41 U9158 ( .I0(ram[15423]), .I1(ram[15415]), .I2(ram[15407]), .I3(
        ram[15399]), .S0(n27336), .S1(n26861), .ZN(n26041) );
  MUX41 U9159 ( .I0(ram[13759]), .I1(ram[13751]), .I2(ram[13743]), .I3(
        ram[13735]), .S0(n27332), .S1(n26857), .ZN(n25971) );
  MUX41 U9160 ( .I0(ram[13503]), .I1(ram[13495]), .I2(ram[13487]), .I3(
        ram[13479]), .S0(n27332), .S1(n26857), .ZN(n25961) );
  MUX41 U9161 ( .I0(ram[13375]), .I1(ram[13367]), .I2(ram[13359]), .I3(
        ram[13351]), .S0(n27331), .S1(n26856), .ZN(n25956) );
  MUX41 U9162 ( .I0(n25427), .I1(n25428), .I2(n25429), .I3(n25430), .S0(
        n26263), .S1(n26381), .ZN(n25426) );
  MUX41 U9163 ( .I0(ram[703]), .I1(ram[695]), .I2(ram[687]), .I3(ram[679]), .S0(n27301), .S1(n26826), .ZN(n25428) );
  MUX41 U9164 ( .I0(ram[671]), .I1(ram[663]), .I2(ram[655]), .I3(ram[647]), .S0(n27301), .S1(n26826), .ZN(n25430) );
  MUX41 U9165 ( .I0(ram[767]), .I1(ram[759]), .I2(ram[751]), .I3(ram[743]), .S0(n27301), .S1(n26826), .ZN(n25427) );
  MUX41 U9166 ( .I0(ram[7615]), .I1(ram[7607]), .I2(ram[7599]), .I3(
        ram[7591]), .S0(n27317), .S1(n26842), .ZN(n25714) );
  MUX41 U9167 ( .I0(ram[7359]), .I1(ram[7351]), .I2(ram[7343]), .I3(
        ram[7335]), .S0(n27317), .S1(n26842), .ZN(n25704) );
  MUX41 U9168 ( .I0(ram[7231]), .I1(ram[7223]), .I2(ram[7215]), .I3(
        ram[7207]), .S0(n27316), .S1(n26841), .ZN(n25699) );
  MUX41 U9169 ( .I0(ram[11711]), .I1(ram[11703]), .I2(ram[11695]), .I3(
        ram[11687]), .S0(n27327), .S1(n26852), .ZN(n25885) );
  MUX41 U9170 ( .I0(ram[11455]), .I1(ram[11447]), .I2(ram[11439]), .I3(
        ram[11431]), .S0(n27327), .S1(n26852), .ZN(n25875) );
  MUX41 U9171 ( .I0(ram[9663]), .I1(ram[9655]), .I2(ram[9647]), .I3(
        ram[9639]), .S0(n27322), .S1(n26847), .ZN(n25800) );
  MUX41 U9172 ( .I0(n21277), .I1(n21278), .I2(n21279), .I3(n21280), .S0(
        n26203), .S1(n26321), .ZN(n21276) );
  MUX41 U9173 ( .I0(ram[16056]), .I1(ram[16048]), .I2(ram[16040]), .I3(
        ram[16032]), .S0(n27062), .S1(n26587), .ZN(n21278) );
  MUX41 U9174 ( .I0(ram[16024]), .I1(ram[16016]), .I2(ram[16008]), .I3(
        ram[16000]), .S0(n27062), .S1(n26587), .ZN(n21280) );
  MUX41 U9175 ( .I0(ram[16120]), .I1(ram[16112]), .I2(ram[16104]), .I3(
        ram[16096]), .S0(n27062), .S1(n26587), .ZN(n21277) );
  MUX41 U9176 ( .I0(n21237), .I1(n21238), .I2(n21239), .I3(n21240), .S0(
        n26203), .S1(n26321), .ZN(n21236) );
  MUX41 U9177 ( .I0(ram[15000]), .I1(ram[14992]), .I2(ram[14984]), .I3(
        ram[14976]), .S0(n27059), .S1(n26584), .ZN(n21240) );
  MUX41 U9178 ( .I0(ram[15032]), .I1(ram[15024]), .I2(ram[15016]), .I3(
        ram[15008]), .S0(n27060), .S1(n26585), .ZN(n21238) );
  MUX41 U9179 ( .I0(ram[15096]), .I1(ram[15088]), .I2(ram[15080]), .I3(
        ram[15072]), .S0(n27060), .S1(n26585), .ZN(n21237) );
  MUX41 U9180 ( .I0(n21217), .I1(n21218), .I2(n21219), .I3(n21220), .S0(
        n26202), .S1(n26320), .ZN(n21216) );
  MUX41 U9181 ( .I0(ram[14520]), .I1(ram[14512]), .I2(ram[14504]), .I3(
        ram[14496]), .S0(n27058), .S1(n26583), .ZN(n21218) );
  MUX41 U9182 ( .I0(ram[14488]), .I1(ram[14480]), .I2(ram[14472]), .I3(
        ram[14464]), .S0(n27058), .S1(n26583), .ZN(n21220) );
  MUX41 U9183 ( .I0(ram[14584]), .I1(ram[14576]), .I2(ram[14568]), .I3(
        ram[14560]), .S0(n27058), .S1(n26583), .ZN(n21217) );
  MUX41 U9184 ( .I0(n21192), .I1(n21193), .I2(n21194), .I3(n21195), .S0(
        n26202), .S1(n26320), .ZN(n21191) );
  MUX41 U9185 ( .I0(ram[14008]), .I1(ram[14000]), .I2(ram[13992]), .I3(
        ram[13984]), .S0(n27057), .S1(n26582), .ZN(n21193) );
  MUX41 U9186 ( .I0(ram[13976]), .I1(ram[13968]), .I2(ram[13960]), .I3(
        ram[13952]), .S0(n27057), .S1(n26582), .ZN(n21195) );
  MUX41 U9187 ( .I0(ram[14072]), .I1(ram[14064]), .I2(ram[14056]), .I3(
        ram[14048]), .S0(n27057), .S1(n26582), .ZN(n21192) );
  MUX41 U9188 ( .I0(n21152), .I1(n21153), .I2(n21154), .I3(n21155), .S0(
        n26202), .S1(n26320), .ZN(n21151) );
  MUX41 U9189 ( .I0(ram[12952]), .I1(ram[12944]), .I2(ram[12936]), .I3(
        ram[12928]), .S0(n27055), .S1(n26580), .ZN(n21155) );
  MUX41 U9190 ( .I0(ram[12984]), .I1(ram[12976]), .I2(ram[12968]), .I3(
        ram[12960]), .S0(n27055), .S1(n26580), .ZN(n21153) );
  MUX41 U9191 ( .I0(ram[13048]), .I1(ram[13040]), .I2(ram[13032]), .I3(
        ram[13024]), .S0(n27055), .S1(n26580), .ZN(n21152) );
  MUX41 U9192 ( .I0(n21132), .I1(n21133), .I2(n21134), .I3(n21135), .S0(
        n26201), .S1(n26319), .ZN(n21131) );
  MUX41 U9193 ( .I0(ram[12472]), .I1(ram[12464]), .I2(ram[12456]), .I3(
        ram[12448]), .S0(n27053), .S1(n26578), .ZN(n21133) );
  MUX41 U9194 ( .I0(ram[12440]), .I1(ram[12432]), .I2(ram[12424]), .I3(
        ram[12416]), .S0(n27053), .S1(n26578), .ZN(n21135) );
  MUX41 U9195 ( .I0(ram[12536]), .I1(ram[12528]), .I2(ram[12520]), .I3(
        ram[12512]), .S0(n27054), .S1(n26579), .ZN(n21132) );
  MUX41 U9196 ( .I0(n20935), .I1(n20936), .I2(n20937), .I3(n20938), .S0(
        n26198), .S1(n26316), .ZN(n20934) );
  MUX41 U9197 ( .I0(ram[7864]), .I1(ram[7856]), .I2(ram[7848]), .I3(
        ram[7840]), .S0(n27042), .S1(n26567), .ZN(n20936) );
  MUX41 U9198 ( .I0(ram[7832]), .I1(ram[7824]), .I2(ram[7816]), .I3(
        ram[7808]), .S0(n27042), .S1(n26567), .ZN(n20938) );
  MUX41 U9199 ( .I0(ram[7928]), .I1(ram[7920]), .I2(ram[7912]), .I3(
        ram[7904]), .S0(n27042), .S1(n26567), .ZN(n20935) );
  MUX41 U9200 ( .I0(n20875), .I1(n20876), .I2(n20877), .I3(n20878), .S0(
        n26198), .S1(n26316), .ZN(n20874) );
  MUX41 U9201 ( .I0(ram[6328]), .I1(ram[6320]), .I2(ram[6312]), .I3(
        ram[6304]), .S0(n27039), .S1(n26564), .ZN(n20876) );
  MUX41 U9202 ( .I0(ram[6296]), .I1(ram[6288]), .I2(ram[6280]), .I3(
        ram[6272]), .S0(n27039), .S1(n26564), .ZN(n20878) );
  MUX41 U9203 ( .I0(ram[6392]), .I1(ram[6384]), .I2(ram[6376]), .I3(
        ram[6368]), .S0(n27039), .S1(n26564), .ZN(n20875) );
  MUX41 U9204 ( .I0(n20895), .I1(n20896), .I2(n20897), .I3(n20898), .S0(
        n26198), .S1(n26316), .ZN(n20894) );
  MUX41 U9205 ( .I0(ram[6840]), .I1(ram[6832]), .I2(ram[6824]), .I3(
        ram[6816]), .S0(n27040), .S1(n26565), .ZN(n20896) );
  MUX41 U9206 ( .I0(ram[6808]), .I1(ram[6800]), .I2(ram[6792]), .I3(
        ram[6784]), .S0(n27040), .S1(n26565), .ZN(n20898) );
  MUX41 U9207 ( .I0(ram[6904]), .I1(ram[6896]), .I2(ram[6888]), .I3(
        ram[6880]), .S0(n27040), .S1(n26565), .ZN(n20895) );
  MUX41 U9208 ( .I0(n20850), .I1(n20851), .I2(n20852), .I3(n20853), .S0(
        n26197), .S1(n26315), .ZN(n20849) );
  MUX41 U9209 ( .I0(ram[5816]), .I1(ram[5808]), .I2(ram[5800]), .I3(
        ram[5792]), .S0(n27037), .S1(n26562), .ZN(n20851) );
  MUX41 U9210 ( .I0(ram[5784]), .I1(ram[5776]), .I2(ram[5768]), .I3(
        ram[5760]), .S0(n27037), .S1(n26562), .ZN(n20853) );
  MUX41 U9211 ( .I0(ram[5880]), .I1(ram[5872]), .I2(ram[5864]), .I3(
        ram[5856]), .S0(n27038), .S1(n26563), .ZN(n20850) );
  MUX41 U9212 ( .I0(n21106), .I1(n21107), .I2(n21108), .I3(n21109), .S0(
        n26201), .S1(n26319), .ZN(n21105) );
  MUX41 U9213 ( .I0(ram[11960]), .I1(ram[11952]), .I2(ram[11944]), .I3(
        ram[11936]), .S0(n27052), .S1(n26577), .ZN(n21107) );
  MUX41 U9214 ( .I0(ram[11928]), .I1(ram[11920]), .I2(ram[11912]), .I3(
        ram[11904]), .S0(n27052), .S1(n26577), .ZN(n21109) );
  MUX41 U9215 ( .I0(ram[12024]), .I1(ram[12016]), .I2(ram[12008]), .I3(
        ram[12000]), .S0(n27052), .S1(n26577), .ZN(n21106) );
  MUX41 U9216 ( .I0(n21046), .I1(n21047), .I2(n21048), .I3(n21049), .S0(
        n26200), .S1(n26318), .ZN(n21045) );
  MUX41 U9217 ( .I0(ram[10424]), .I1(ram[10416]), .I2(ram[10408]), .I3(
        ram[10400]), .S0(n27048), .S1(n26573), .ZN(n21047) );
  MUX41 U9218 ( .I0(ram[10392]), .I1(ram[10384]), .I2(ram[10376]), .I3(
        ram[10368]), .S0(n27048), .S1(n26573), .ZN(n21049) );
  MUX41 U9219 ( .I0(ram[10488]), .I1(ram[10480]), .I2(ram[10472]), .I3(
        ram[10464]), .S0(n27049), .S1(n26574), .ZN(n21046) );
  MUX41 U9220 ( .I0(n21021), .I1(n21022), .I2(n21023), .I3(n21024), .S0(
        n26200), .S1(n26318), .ZN(n21020) );
  MUX41 U9221 ( .I0(ram[9912]), .I1(ram[9904]), .I2(ram[9896]), .I3(
        ram[9888]), .S0(n27047), .S1(n26572), .ZN(n21022) );
  MUX41 U9222 ( .I0(ram[9880]), .I1(ram[9872]), .I2(ram[9864]), .I3(
        ram[9856]), .S0(n27047), .S1(n26572), .ZN(n21024) );
  MUX41 U9223 ( .I0(ram[9976]), .I1(ram[9968]), .I2(ram[9960]), .I3(
        ram[9952]), .S0(n27047), .S1(n26572), .ZN(n21021) );
  MUX41 U9224 ( .I0(n20961), .I1(n20962), .I2(n20963), .I3(n20964), .S0(
        n26199), .S1(n26317), .ZN(n20960) );
  MUX41 U9225 ( .I0(ram[8376]), .I1(ram[8368]), .I2(ram[8360]), .I3(
        ram[8352]), .S0(n27044), .S1(n26569), .ZN(n20962) );
  MUX41 U9226 ( .I0(ram[8344]), .I1(ram[8336]), .I2(ram[8328]), .I3(
        ram[8320]), .S0(n27043), .S1(n26568), .ZN(n20964) );
  MUX41 U9227 ( .I0(ram[8440]), .I1(ram[8432]), .I2(ram[8424]), .I3(
        ram[8416]), .S0(n27044), .S1(n26569), .ZN(n20961) );
  MUX41 U9228 ( .I0(n21961), .I1(n21962), .I2(n21963), .I3(n21964), .S0(
        n26213), .S1(n26331), .ZN(n21960) );
  MUX41 U9229 ( .I0(ram[16057]), .I1(ram[16049]), .I2(ram[16041]), .I3(
        ram[16033]), .S0(n27101), .S1(n26626), .ZN(n21962) );
  MUX41 U9230 ( .I0(ram[16025]), .I1(ram[16017]), .I2(ram[16009]), .I3(
        ram[16001]), .S0(n27101), .S1(n26626), .ZN(n21964) );
  MUX41 U9231 ( .I0(ram[16121]), .I1(ram[16113]), .I2(ram[16105]), .I3(
        ram[16097]), .S0(n27102), .S1(n26627), .ZN(n21961) );
  MUX41 U9232 ( .I0(n21921), .I1(n21922), .I2(n21923), .I3(n21924), .S0(
        n26213), .S1(n26331), .ZN(n21920) );
  MUX41 U9233 ( .I0(ram[15001]), .I1(ram[14993]), .I2(ram[14985]), .I3(
        ram[14977]), .S0(n27099), .S1(n26624), .ZN(n21924) );
  MUX41 U9234 ( .I0(ram[15033]), .I1(ram[15025]), .I2(ram[15017]), .I3(
        ram[15009]), .S0(n27099), .S1(n26624), .ZN(n21922) );
  MUX41 U9235 ( .I0(ram[15097]), .I1(ram[15089]), .I2(ram[15081]), .I3(
        ram[15073]), .S0(n27099), .S1(n26624), .ZN(n21921) );
  MUX41 U9236 ( .I0(n21901), .I1(n21902), .I2(n21903), .I3(n21904), .S0(
        n26212), .S1(n26330), .ZN(n21900) );
  MUX41 U9237 ( .I0(ram[14521]), .I1(ram[14513]), .I2(ram[14505]), .I3(
        ram[14497]), .S0(n27098), .S1(n26623), .ZN(n21902) );
  MUX41 U9238 ( .I0(ram[14489]), .I1(ram[14481]), .I2(ram[14473]), .I3(
        ram[14465]), .S0(n27098), .S1(n26623), .ZN(n21904) );
  MUX41 U9239 ( .I0(ram[14585]), .I1(ram[14577]), .I2(ram[14569]), .I3(
        ram[14561]), .S0(n27098), .S1(n26623), .ZN(n21901) );
  MUX41 U9240 ( .I0(n21876), .I1(n21877), .I2(n21878), .I3(n21879), .S0(
        n26212), .S1(n26330), .ZN(n21875) );
  MUX41 U9241 ( .I0(ram[14009]), .I1(ram[14001]), .I2(ram[13993]), .I3(
        ram[13985]), .S0(n27096), .S1(n26621), .ZN(n21877) );
  MUX41 U9242 ( .I0(ram[13977]), .I1(ram[13969]), .I2(ram[13961]), .I3(
        ram[13953]), .S0(n27096), .S1(n26621), .ZN(n21879) );
  MUX41 U9243 ( .I0(ram[14073]), .I1(ram[14065]), .I2(ram[14057]), .I3(
        ram[14049]), .S0(n27097), .S1(n26622), .ZN(n21876) );
  MUX41 U9244 ( .I0(n21836), .I1(n21837), .I2(n21838), .I3(n21839), .S0(
        n26211), .S1(n26329), .ZN(n21835) );
  MUX41 U9245 ( .I0(ram[12953]), .I1(ram[12945]), .I2(ram[12937]), .I3(
        ram[12929]), .S0(n27094), .S1(n26619), .ZN(n21839) );
  MUX41 U9246 ( .I0(ram[12985]), .I1(ram[12977]), .I2(ram[12969]), .I3(
        ram[12961]), .S0(n27094), .S1(n26619), .ZN(n21837) );
  MUX41 U9247 ( .I0(ram[13049]), .I1(ram[13041]), .I2(ram[13033]), .I3(
        ram[13025]), .S0(n27094), .S1(n26619), .ZN(n21836) );
  MUX41 U9248 ( .I0(n21816), .I1(n21817), .I2(n21818), .I3(n21819), .S0(
        n26211), .S1(n26329), .ZN(n21815) );
  MUX41 U9249 ( .I0(ram[12473]), .I1(ram[12465]), .I2(ram[12457]), .I3(
        ram[12449]), .S0(n27093), .S1(n26618), .ZN(n21817) );
  MUX41 U9250 ( .I0(ram[12441]), .I1(ram[12433]), .I2(ram[12425]), .I3(
        ram[12417]), .S0(n27093), .S1(n26618), .ZN(n21819) );
  MUX41 U9251 ( .I0(ram[12537]), .I1(ram[12529]), .I2(ram[12521]), .I3(
        ram[12513]), .S0(n27093), .S1(n26618), .ZN(n21816) );
  MUX41 U9252 ( .I0(n21619), .I1(n21620), .I2(n21621), .I3(n21622), .S0(
        n26208), .S1(n26326), .ZN(n21618) );
  MUX41 U9253 ( .I0(ram[7865]), .I1(ram[7857]), .I2(ram[7849]), .I3(
        ram[7841]), .S0(n27082), .S1(n26607), .ZN(n21620) );
  MUX41 U9254 ( .I0(ram[7833]), .I1(ram[7825]), .I2(ram[7817]), .I3(
        ram[7809]), .S0(n27082), .S1(n26607), .ZN(n21622) );
  MUX41 U9255 ( .I0(ram[7929]), .I1(ram[7921]), .I2(ram[7913]), .I3(
        ram[7905]), .S0(n27082), .S1(n26607), .ZN(n21619) );
  MUX41 U9256 ( .I0(n21559), .I1(n21560), .I2(n21561), .I3(n21562), .S0(
        n26207), .S1(n26325), .ZN(n21558) );
  MUX41 U9257 ( .I0(ram[6329]), .I1(ram[6321]), .I2(ram[6313]), .I3(
        ram[6305]), .S0(n27078), .S1(n26603), .ZN(n21560) );
  MUX41 U9258 ( .I0(ram[6297]), .I1(ram[6289]), .I2(ram[6281]), .I3(
        ram[6273]), .S0(n27078), .S1(n26603), .ZN(n21562) );
  MUX41 U9259 ( .I0(ram[6393]), .I1(ram[6385]), .I2(ram[6377]), .I3(
        ram[6369]), .S0(n27078), .S1(n26603), .ZN(n21559) );
  MUX41 U9260 ( .I0(n21579), .I1(n21580), .I2(n21581), .I3(n21582), .S0(
        n26208), .S1(n26326), .ZN(n21578) );
  MUX41 U9261 ( .I0(ram[6841]), .I1(ram[6833]), .I2(ram[6825]), .I3(
        ram[6817]), .S0(n27079), .S1(n26604), .ZN(n21580) );
  MUX41 U9262 ( .I0(ram[6809]), .I1(ram[6801]), .I2(ram[6793]), .I3(
        ram[6785]), .S0(n27079), .S1(n26604), .ZN(n21582) );
  MUX41 U9263 ( .I0(ram[6905]), .I1(ram[6897]), .I2(ram[6889]), .I3(
        ram[6881]), .S0(n27079), .S1(n26604), .ZN(n21579) );
  MUX41 U9264 ( .I0(n21534), .I1(n21535), .I2(n21536), .I3(n21537), .S0(
        n26207), .S1(n26325), .ZN(n21533) );
  MUX41 U9265 ( .I0(ram[5817]), .I1(ram[5809]), .I2(ram[5801]), .I3(
        ram[5793]), .S0(n27077), .S1(n26602), .ZN(n21535) );
  MUX41 U9266 ( .I0(ram[5785]), .I1(ram[5777]), .I2(ram[5769]), .I3(
        ram[5761]), .S0(n27077), .S1(n26602), .ZN(n21537) );
  MUX41 U9267 ( .I0(ram[5881]), .I1(ram[5873]), .I2(ram[5865]), .I3(
        ram[5857]), .S0(n27077), .S1(n26602), .ZN(n21534) );
  MUX41 U9268 ( .I0(n21790), .I1(n21791), .I2(n21792), .I3(n21793), .S0(
        n26211), .S1(n26329), .ZN(n21789) );
  MUX41 U9269 ( .I0(ram[11961]), .I1(ram[11953]), .I2(ram[11945]), .I3(
        ram[11937]), .S0(n27092), .S1(n26617), .ZN(n21791) );
  MUX41 U9270 ( .I0(ram[11929]), .I1(ram[11921]), .I2(ram[11913]), .I3(
        ram[11905]), .S0(n27091), .S1(n26616), .ZN(n21793) );
  MUX41 U9271 ( .I0(ram[12025]), .I1(ram[12017]), .I2(ram[12009]), .I3(
        ram[12001]), .S0(n27092), .S1(n26617), .ZN(n21790) );
  MUX41 U9272 ( .I0(n21730), .I1(n21731), .I2(n21732), .I3(n21733), .S0(
        n26210), .S1(n26328), .ZN(n21729) );
  MUX41 U9273 ( .I0(ram[10425]), .I1(ram[10417]), .I2(ram[10409]), .I3(
        ram[10401]), .S0(n27088), .S1(n26613), .ZN(n21731) );
  MUX41 U9274 ( .I0(ram[10393]), .I1(ram[10385]), .I2(ram[10377]), .I3(
        ram[10369]), .S0(n27088), .S1(n26613), .ZN(n21733) );
  MUX41 U9275 ( .I0(ram[10489]), .I1(ram[10481]), .I2(ram[10473]), .I3(
        ram[10465]), .S0(n27088), .S1(n26613), .ZN(n21730) );
  MUX41 U9276 ( .I0(n21705), .I1(n21706), .I2(n21707), .I3(n21708), .S0(
        n26210), .S1(n26328), .ZN(n21704) );
  MUX41 U9277 ( .I0(ram[9913]), .I1(ram[9905]), .I2(ram[9897]), .I3(
        ram[9889]), .S0(n27087), .S1(n26612), .ZN(n21706) );
  MUX41 U9278 ( .I0(ram[9881]), .I1(ram[9873]), .I2(ram[9865]), .I3(
        ram[9857]), .S0(n27087), .S1(n26612), .ZN(n21708) );
  MUX41 U9279 ( .I0(ram[9977]), .I1(ram[9969]), .I2(ram[9961]), .I3(
        ram[9953]), .S0(n27087), .S1(n26612), .ZN(n21705) );
  MUX41 U9280 ( .I0(n21645), .I1(n21646), .I2(n21647), .I3(n21648), .S0(
        n26209), .S1(n26327), .ZN(n21644) );
  MUX41 U9281 ( .I0(ram[8377]), .I1(ram[8369]), .I2(ram[8361]), .I3(
        ram[8353]), .S0(n27083), .S1(n26608), .ZN(n21646) );
  MUX41 U9282 ( .I0(ram[8345]), .I1(ram[8337]), .I2(ram[8329]), .I3(
        ram[8321]), .S0(n27083), .S1(n26608), .ZN(n21648) );
  MUX41 U9283 ( .I0(ram[8441]), .I1(ram[8433]), .I2(ram[8425]), .I3(
        ram[8417]), .S0(n27083), .S1(n26608), .ZN(n21645) );
  MUX41 U9284 ( .I0(n22645), .I1(n22646), .I2(n22647), .I3(n22648), .S0(
        n26223), .S1(n26341), .ZN(n22644) );
  MUX41 U9285 ( .I0(ram[16058]), .I1(ram[16050]), .I2(ram[16042]), .I3(
        ram[16034]), .S0(n27141), .S1(n26666), .ZN(n22646) );
  MUX41 U9286 ( .I0(ram[16026]), .I1(ram[16018]), .I2(ram[16010]), .I3(
        ram[16002]), .S0(n27141), .S1(n26666), .ZN(n22648) );
  MUX41 U9287 ( .I0(ram[16122]), .I1(ram[16114]), .I2(ram[16106]), .I3(
        ram[16098]), .S0(n27141), .S1(n26666), .ZN(n22645) );
  MUX41 U9288 ( .I0(n22605), .I1(n22606), .I2(n22607), .I3(n22608), .S0(
        n26222), .S1(n26340), .ZN(n22604) );
  MUX41 U9289 ( .I0(ram[15002]), .I1(ram[14994]), .I2(ram[14986]), .I3(
        ram[14978]), .S0(n27138), .S1(n26663), .ZN(n22608) );
  MUX41 U9290 ( .I0(ram[15034]), .I1(ram[15026]), .I2(ram[15018]), .I3(
        ram[15010]), .S0(n27138), .S1(n26663), .ZN(n22606) );
  MUX41 U9291 ( .I0(ram[15098]), .I1(ram[15090]), .I2(ram[15082]), .I3(
        ram[15074]), .S0(n27138), .S1(n26663), .ZN(n22605) );
  MUX41 U9292 ( .I0(n22585), .I1(n22586), .I2(n22587), .I3(n22588), .S0(
        n26222), .S1(n26340), .ZN(n22584) );
  MUX41 U9293 ( .I0(ram[14522]), .I1(ram[14514]), .I2(ram[14506]), .I3(
        ram[14498]), .S0(n27137), .S1(n26662), .ZN(n22586) );
  MUX41 U9294 ( .I0(ram[14490]), .I1(ram[14482]), .I2(ram[14474]), .I3(
        ram[14466]), .S0(n27137), .S1(n26662), .ZN(n22588) );
  MUX41 U9295 ( .I0(ram[14586]), .I1(ram[14578]), .I2(ram[14570]), .I3(
        ram[14562]), .S0(n27137), .S1(n26662), .ZN(n22585) );
  MUX41 U9296 ( .I0(n22560), .I1(n22561), .I2(n22562), .I3(n22563), .S0(
        n26222), .S1(n26340), .ZN(n22559) );
  MUX41 U9297 ( .I0(ram[14010]), .I1(ram[14002]), .I2(ram[13994]), .I3(
        ram[13986]), .S0(n27136), .S1(n26661), .ZN(n22561) );
  MUX41 U9298 ( .I0(ram[13978]), .I1(ram[13970]), .I2(ram[13962]), .I3(
        ram[13954]), .S0(n27136), .S1(n26661), .ZN(n22563) );
  MUX41 U9299 ( .I0(ram[14074]), .I1(ram[14066]), .I2(ram[14058]), .I3(
        ram[14050]), .S0(n27136), .S1(n26661), .ZN(n22560) );
  MUX41 U9300 ( .I0(n22520), .I1(n22521), .I2(n22522), .I3(n22523), .S0(
        n26221), .S1(n26339), .ZN(n22519) );
  MUX41 U9301 ( .I0(ram[12954]), .I1(ram[12946]), .I2(ram[12938]), .I3(
        ram[12930]), .S0(n27133), .S1(n26658), .ZN(n22523) );
  MUX41 U9302 ( .I0(ram[12986]), .I1(ram[12978]), .I2(ram[12970]), .I3(
        ram[12962]), .S0(n27133), .S1(n26658), .ZN(n22521) );
  MUX41 U9303 ( .I0(ram[13050]), .I1(ram[13042]), .I2(ram[13034]), .I3(
        ram[13026]), .S0(n27134), .S1(n26659), .ZN(n22520) );
  MUX41 U9304 ( .I0(n22500), .I1(n22501), .I2(n22502), .I3(n22503), .S0(
        n26221), .S1(n26339), .ZN(n22499) );
  MUX41 U9305 ( .I0(ram[12474]), .I1(ram[12466]), .I2(ram[12458]), .I3(
        ram[12450]), .S0(n27132), .S1(n26657), .ZN(n22501) );
  MUX41 U9306 ( .I0(ram[12442]), .I1(ram[12434]), .I2(ram[12426]), .I3(
        ram[12418]), .S0(n27132), .S1(n26657), .ZN(n22503) );
  MUX41 U9307 ( .I0(ram[12538]), .I1(ram[12530]), .I2(ram[12522]), .I3(
        ram[12514]), .S0(n27132), .S1(n26657), .ZN(n22500) );
  MUX41 U9308 ( .I0(n22303), .I1(n22304), .I2(n22305), .I3(n22306), .S0(
        n26218), .S1(n26336), .ZN(n22302) );
  MUX41 U9309 ( .I0(ram[7866]), .I1(ram[7858]), .I2(ram[7850]), .I3(
        ram[7842]), .S0(n27121), .S1(n26646), .ZN(n22304) );
  MUX41 U9310 ( .I0(ram[7834]), .I1(ram[7826]), .I2(ram[7818]), .I3(
        ram[7810]), .S0(n27121), .S1(n26646), .ZN(n22306) );
  MUX41 U9311 ( .I0(ram[7930]), .I1(ram[7922]), .I2(ram[7914]), .I3(
        ram[7906]), .S0(n27121), .S1(n26646), .ZN(n22303) );
  MUX41 U9312 ( .I0(n22243), .I1(n22244), .I2(n22245), .I3(n22246), .S0(
        n26217), .S1(n26335), .ZN(n22242) );
  MUX41 U9313 ( .I0(ram[6330]), .I1(ram[6322]), .I2(ram[6314]), .I3(
        ram[6306]), .S0(n27117), .S1(n26642), .ZN(n22244) );
  MUX41 U9314 ( .I0(ram[6298]), .I1(ram[6290]), .I2(ram[6282]), .I3(
        ram[6274]), .S0(n27117), .S1(n26642), .ZN(n22246) );
  MUX41 U9315 ( .I0(ram[6394]), .I1(ram[6386]), .I2(ram[6378]), .I3(
        ram[6370]), .S0(n27118), .S1(n26643), .ZN(n22243) );
  MUX41 U9316 ( .I0(n22263), .I1(n22264), .I2(n22265), .I3(n22266), .S0(
        n26218), .S1(n26336), .ZN(n22262) );
  MUX41 U9317 ( .I0(ram[6842]), .I1(ram[6834]), .I2(ram[6826]), .I3(
        ram[6818]), .S0(n27119), .S1(n26644), .ZN(n22264) );
  MUX41 U9318 ( .I0(ram[6810]), .I1(ram[6802]), .I2(ram[6794]), .I3(
        ram[6786]), .S0(n27119), .S1(n26644), .ZN(n22266) );
  MUX41 U9319 ( .I0(ram[6906]), .I1(ram[6898]), .I2(ram[6890]), .I3(
        ram[6882]), .S0(n27119), .S1(n26644), .ZN(n22263) );
  MUX41 U9320 ( .I0(n22218), .I1(n22219), .I2(n22220), .I3(n22221), .S0(
        n26217), .S1(n26335), .ZN(n22217) );
  MUX41 U9321 ( .I0(ram[5818]), .I1(ram[5810]), .I2(ram[5802]), .I3(
        ram[5794]), .S0(n27116), .S1(n26641), .ZN(n22219) );
  MUX41 U9322 ( .I0(ram[5786]), .I1(ram[5778]), .I2(ram[5770]), .I3(
        ram[5762]), .S0(n27116), .S1(n26641), .ZN(n22221) );
  MUX41 U9323 ( .I0(ram[5882]), .I1(ram[5874]), .I2(ram[5866]), .I3(
        ram[5858]), .S0(n27116), .S1(n26641), .ZN(n22218) );
  MUX41 U9324 ( .I0(n22474), .I1(n22475), .I2(n22476), .I3(n22477), .S0(
        n26221), .S1(n26339), .ZN(n22473) );
  MUX41 U9325 ( .I0(ram[11962]), .I1(ram[11954]), .I2(ram[11946]), .I3(
        ram[11938]), .S0(n27131), .S1(n26656), .ZN(n22475) );
  MUX41 U9326 ( .I0(ram[11930]), .I1(ram[11922]), .I2(ram[11914]), .I3(
        ram[11906]), .S0(n27131), .S1(n26656), .ZN(n22477) );
  MUX41 U9327 ( .I0(ram[12026]), .I1(ram[12018]), .I2(ram[12010]), .I3(
        ram[12002]), .S0(n27131), .S1(n26656), .ZN(n22474) );
  MUX41 U9328 ( .I0(n22414), .I1(n22415), .I2(n22416), .I3(n22417), .S0(
        n26220), .S1(n26338), .ZN(n22413) );
  MUX41 U9329 ( .I0(ram[10426]), .I1(ram[10418]), .I2(ram[10410]), .I3(
        ram[10402]), .S0(n27127), .S1(n26652), .ZN(n22415) );
  MUX41 U9330 ( .I0(ram[10394]), .I1(ram[10386]), .I2(ram[10378]), .I3(
        ram[10370]), .S0(n27127), .S1(n26652), .ZN(n22417) );
  MUX41 U9331 ( .I0(ram[10490]), .I1(ram[10482]), .I2(ram[10474]), .I3(
        ram[10466]), .S0(n27127), .S1(n26652), .ZN(n22414) );
  MUX41 U9332 ( .I0(n22434), .I1(n22435), .I2(n22436), .I3(n22437), .S0(
        n26220), .S1(n26338), .ZN(n22433) );
  MUX41 U9333 ( .I0(ram[10938]), .I1(ram[10930]), .I2(ram[10922]), .I3(
        ram[10914]), .S0(n27128), .S1(n26653), .ZN(n22435) );
  MUX41 U9334 ( .I0(ram[10906]), .I1(ram[10898]), .I2(ram[10890]), .I3(
        ram[10882]), .S0(n27128), .S1(n26653), .ZN(n22437) );
  MUX41 U9335 ( .I0(ram[11002]), .I1(ram[10994]), .I2(ram[10986]), .I3(
        ram[10978]), .S0(n27129), .S1(n26654), .ZN(n22434) );
  MUX41 U9336 ( .I0(n22389), .I1(n22390), .I2(n22391), .I3(n22392), .S0(
        n26219), .S1(n26337), .ZN(n22388) );
  MUX41 U9337 ( .I0(ram[9914]), .I1(ram[9906]), .I2(ram[9898]), .I3(
        ram[9890]), .S0(n27126), .S1(n26651), .ZN(n22390) );
  MUX41 U9338 ( .I0(ram[9882]), .I1(ram[9874]), .I2(ram[9866]), .I3(
        ram[9858]), .S0(n27126), .S1(n26651), .ZN(n22392) );
  MUX41 U9339 ( .I0(ram[9978]), .I1(ram[9970]), .I2(ram[9962]), .I3(
        ram[9954]), .S0(n27126), .S1(n26651), .ZN(n22389) );
  MUX41 U9340 ( .I0(n22329), .I1(n22330), .I2(n22331), .I3(n22332), .S0(
        n26218), .S1(n26336), .ZN(n22328) );
  MUX41 U9341 ( .I0(ram[8378]), .I1(ram[8370]), .I2(ram[8362]), .I3(
        ram[8354]), .S0(n27122), .S1(n26647), .ZN(n22330) );
  MUX41 U9342 ( .I0(ram[8346]), .I1(ram[8338]), .I2(ram[8330]), .I3(
        ram[8322]), .S0(n27122), .S1(n26647), .ZN(n22332) );
  MUX41 U9343 ( .I0(ram[8442]), .I1(ram[8434]), .I2(ram[8426]), .I3(
        ram[8418]), .S0(n27122), .S1(n26647), .ZN(n22329) );
  MUX41 U9344 ( .I0(n23329), .I1(n23330), .I2(n23331), .I3(n23332), .S0(
        n26233), .S1(n26351), .ZN(n23328) );
  MUX41 U9345 ( .I0(ram[16059]), .I1(ram[16051]), .I2(ram[16043]), .I3(
        ram[16035]), .S0(n27180), .S1(n26705), .ZN(n23330) );
  MUX41 U9346 ( .I0(ram[16027]), .I1(ram[16019]), .I2(ram[16011]), .I3(
        ram[16003]), .S0(n27180), .S1(n26705), .ZN(n23332) );
  MUX41 U9347 ( .I0(ram[16123]), .I1(ram[16115]), .I2(ram[16107]), .I3(
        ram[16099]), .S0(n27180), .S1(n26705), .ZN(n23329) );
  MUX41 U9348 ( .I0(n23289), .I1(n23290), .I2(n23291), .I3(n23292), .S0(
        n26232), .S1(n26350), .ZN(n23288) );
  MUX41 U9349 ( .I0(ram[15003]), .I1(ram[14995]), .I2(ram[14987]), .I3(
        ram[14979]), .S0(n27178), .S1(n26703), .ZN(n23292) );
  MUX41 U9350 ( .I0(ram[15035]), .I1(ram[15027]), .I2(ram[15019]), .I3(
        ram[15011]), .S0(n27178), .S1(n26703), .ZN(n23290) );
  MUX41 U9351 ( .I0(ram[15099]), .I1(ram[15091]), .I2(ram[15083]), .I3(
        ram[15075]), .S0(n27178), .S1(n26703), .ZN(n23289) );
  MUX41 U9352 ( .I0(n23269), .I1(n23270), .I2(n23271), .I3(n23272), .S0(
        n26232), .S1(n26350), .ZN(n23268) );
  MUX41 U9353 ( .I0(ram[14523]), .I1(ram[14515]), .I2(ram[14507]), .I3(
        ram[14499]), .S0(n27176), .S1(n26701), .ZN(n23270) );
  MUX41 U9354 ( .I0(ram[14491]), .I1(ram[14483]), .I2(ram[14475]), .I3(
        ram[14467]), .S0(n27176), .S1(n26701), .ZN(n23272) );
  MUX41 U9355 ( .I0(ram[14587]), .I1(ram[14579]), .I2(ram[14571]), .I3(
        ram[14563]), .S0(n27177), .S1(n26702), .ZN(n23269) );
  MUX41 U9356 ( .I0(n23244), .I1(n23245), .I2(n23246), .I3(n23247), .S0(
        n26232), .S1(n26350), .ZN(n23243) );
  MUX41 U9357 ( .I0(ram[14011]), .I1(ram[14003]), .I2(ram[13995]), .I3(
        ram[13987]), .S0(n27175), .S1(n26700), .ZN(n23245) );
  MUX41 U9358 ( .I0(ram[13979]), .I1(ram[13971]), .I2(ram[13963]), .I3(
        ram[13955]), .S0(n27175), .S1(n26700), .ZN(n23247) );
  MUX41 U9359 ( .I0(ram[14075]), .I1(ram[14067]), .I2(ram[14059]), .I3(
        ram[14051]), .S0(n27175), .S1(n26700), .ZN(n23244) );
  MUX41 U9360 ( .I0(n23204), .I1(n23205), .I2(n23206), .I3(n23207), .S0(
        n26231), .S1(n26349), .ZN(n23203) );
  MUX41 U9361 ( .I0(ram[12955]), .I1(ram[12947]), .I2(ram[12939]), .I3(
        ram[12931]), .S0(n27173), .S1(n26698), .ZN(n23207) );
  MUX41 U9362 ( .I0(ram[12987]), .I1(ram[12979]), .I2(ram[12971]), .I3(
        ram[12963]), .S0(n27173), .S1(n26698), .ZN(n23205) );
  MUX41 U9363 ( .I0(ram[13051]), .I1(ram[13043]), .I2(ram[13035]), .I3(
        ram[13027]), .S0(n27173), .S1(n26698), .ZN(n23204) );
  MUX41 U9364 ( .I0(n23184), .I1(n23185), .I2(n23186), .I3(n23187), .S0(
        n26231), .S1(n26349), .ZN(n23183) );
  MUX41 U9365 ( .I0(ram[12475]), .I1(ram[12467]), .I2(ram[12459]), .I3(
        ram[12451]), .S0(n27172), .S1(n26697), .ZN(n23185) );
  MUX41 U9366 ( .I0(ram[12443]), .I1(ram[12435]), .I2(ram[12427]), .I3(
        ram[12419]), .S0(n27171), .S1(n26696), .ZN(n23187) );
  MUX41 U9367 ( .I0(ram[12539]), .I1(ram[12531]), .I2(ram[12523]), .I3(
        ram[12515]), .S0(n27172), .S1(n26697), .ZN(n23184) );
  MUX41 U9368 ( .I0(n22987), .I1(n22988), .I2(n22989), .I3(n22990), .S0(
        n26228), .S1(n26346), .ZN(n22986) );
  MUX41 U9369 ( .I0(ram[7867]), .I1(ram[7859]), .I2(ram[7851]), .I3(
        ram[7843]), .S0(n27160), .S1(n26685), .ZN(n22988) );
  MUX41 U9370 ( .I0(ram[7835]), .I1(ram[7827]), .I2(ram[7819]), .I3(
        ram[7811]), .S0(n27160), .S1(n26685), .ZN(n22990) );
  MUX41 U9371 ( .I0(ram[7931]), .I1(ram[7923]), .I2(ram[7915]), .I3(
        ram[7907]), .S0(n27161), .S1(n26686), .ZN(n22987) );
  MUX41 U9372 ( .I0(n22927), .I1(n22928), .I2(n22929), .I3(n22930), .S0(
        n26227), .S1(n26345), .ZN(n22926) );
  MUX41 U9373 ( .I0(ram[6331]), .I1(ram[6323]), .I2(ram[6315]), .I3(
        ram[6307]), .S0(n27157), .S1(n26682), .ZN(n22928) );
  MUX41 U9374 ( .I0(ram[6299]), .I1(ram[6291]), .I2(ram[6283]), .I3(
        ram[6275]), .S0(n27157), .S1(n26682), .ZN(n22930) );
  MUX41 U9375 ( .I0(ram[6395]), .I1(ram[6387]), .I2(ram[6379]), .I3(
        ram[6371]), .S0(n27157), .S1(n26682), .ZN(n22927) );
  MUX41 U9376 ( .I0(n22947), .I1(n22948), .I2(n22949), .I3(n22950), .S0(
        n26227), .S1(n26345), .ZN(n22946) );
  MUX41 U9377 ( .I0(ram[6843]), .I1(ram[6835]), .I2(ram[6827]), .I3(
        ram[6819]), .S0(n27158), .S1(n26683), .ZN(n22948) );
  MUX41 U9378 ( .I0(ram[6811]), .I1(ram[6803]), .I2(ram[6795]), .I3(
        ram[6787]), .S0(n27158), .S1(n26683), .ZN(n22950) );
  MUX41 U9379 ( .I0(ram[6907]), .I1(ram[6899]), .I2(ram[6891]), .I3(
        ram[6883]), .S0(n27158), .S1(n26683), .ZN(n22947) );
  MUX41 U9380 ( .I0(n22902), .I1(n22903), .I2(n22904), .I3(n22905), .S0(
        n26227), .S1(n26345), .ZN(n22901) );
  MUX41 U9381 ( .I0(ram[5819]), .I1(ram[5811]), .I2(ram[5803]), .I3(
        ram[5795]), .S0(n27156), .S1(n26681), .ZN(n22903) );
  MUX41 U9382 ( .I0(ram[5787]), .I1(ram[5779]), .I2(ram[5771]), .I3(
        ram[5763]), .S0(n27155), .S1(n26680), .ZN(n22905) );
  MUX41 U9383 ( .I0(ram[5883]), .I1(ram[5875]), .I2(ram[5867]), .I3(
        ram[5859]), .S0(n27156), .S1(n26681), .ZN(n22902) );
  MUX41 U9384 ( .I0(n23158), .I1(n23159), .I2(n23160), .I3(n23161), .S0(
        n26230), .S1(n26348), .ZN(n23157) );
  MUX41 U9385 ( .I0(ram[11963]), .I1(ram[11955]), .I2(ram[11947]), .I3(
        ram[11939]), .S0(n27170), .S1(n26695), .ZN(n23159) );
  MUX41 U9386 ( .I0(ram[11931]), .I1(ram[11923]), .I2(ram[11915]), .I3(
        ram[11907]), .S0(n27170), .S1(n26695), .ZN(n23161) );
  MUX41 U9387 ( .I0(ram[12027]), .I1(ram[12019]), .I2(ram[12011]), .I3(
        ram[12003]), .S0(n27170), .S1(n26695), .ZN(n23158) );
  MUX41 U9388 ( .I0(n23098), .I1(n23099), .I2(n23100), .I3(n23101), .S0(
        n26230), .S1(n26348), .ZN(n23097) );
  MUX41 U9389 ( .I0(ram[10427]), .I1(ram[10419]), .I2(ram[10411]), .I3(
        ram[10403]), .S0(n27167), .S1(n26692), .ZN(n23099) );
  MUX41 U9390 ( .I0(ram[10395]), .I1(ram[10387]), .I2(ram[10379]), .I3(
        ram[10371]), .S0(n27167), .S1(n26692), .ZN(n23101) );
  MUX41 U9391 ( .I0(ram[10491]), .I1(ram[10483]), .I2(ram[10475]), .I3(
        ram[10467]), .S0(n27167), .S1(n26692), .ZN(n23098) );
  MUX41 U9392 ( .I0(n23118), .I1(n23119), .I2(n23120), .I3(n23121), .S0(
        n26230), .S1(n26348), .ZN(n23117) );
  MUX41 U9393 ( .I0(ram[10939]), .I1(ram[10931]), .I2(ram[10923]), .I3(
        ram[10915]), .S0(n27168), .S1(n26693), .ZN(n23119) );
  MUX41 U9394 ( .I0(ram[10907]), .I1(ram[10899]), .I2(ram[10891]), .I3(
        ram[10883]), .S0(n27168), .S1(n26693), .ZN(n23121) );
  MUX41 U9395 ( .I0(ram[11003]), .I1(ram[10995]), .I2(ram[10987]), .I3(
        ram[10979]), .S0(n27168), .S1(n26693), .ZN(n23118) );
  MUX41 U9396 ( .I0(n23073), .I1(n23074), .I2(n23075), .I3(n23076), .S0(
        n26229), .S1(n26347), .ZN(n23072) );
  MUX41 U9397 ( .I0(ram[9915]), .I1(ram[9907]), .I2(ram[9899]), .I3(
        ram[9891]), .S0(n27165), .S1(n26690), .ZN(n23074) );
  MUX41 U9398 ( .I0(ram[9883]), .I1(ram[9875]), .I2(ram[9867]), .I3(
        ram[9859]), .S0(n27165), .S1(n26690), .ZN(n23076) );
  MUX41 U9399 ( .I0(ram[9979]), .I1(ram[9971]), .I2(ram[9963]), .I3(
        ram[9955]), .S0(n27166), .S1(n26691), .ZN(n23073) );
  MUX41 U9400 ( .I0(n23013), .I1(n23014), .I2(n23015), .I3(n23016), .S0(
        n26228), .S1(n26346), .ZN(n23012) );
  MUX41 U9401 ( .I0(ram[8379]), .I1(ram[8371]), .I2(ram[8363]), .I3(
        ram[8355]), .S0(n27162), .S1(n26687), .ZN(n23014) );
  MUX41 U9402 ( .I0(ram[8347]), .I1(ram[8339]), .I2(ram[8331]), .I3(
        ram[8323]), .S0(n27162), .S1(n26687), .ZN(n23016) );
  MUX41 U9403 ( .I0(ram[8443]), .I1(ram[8435]), .I2(ram[8427]), .I3(
        ram[8419]), .S0(n27162), .S1(n26687), .ZN(n23013) );
  MUX41 U9404 ( .I0(n24013), .I1(n24014), .I2(n24015), .I3(n24016), .S0(
        n26243), .S1(n26361), .ZN(n24012) );
  MUX41 U9405 ( .I0(ram[16060]), .I1(ram[16052]), .I2(ram[16044]), .I3(
        ram[16036]), .S0(n27220), .S1(n26745), .ZN(n24014) );
  MUX41 U9406 ( .I0(ram[16028]), .I1(ram[16020]), .I2(ram[16012]), .I3(
        ram[16004]), .S0(n27219), .S1(n26744), .ZN(n24016) );
  MUX41 U9407 ( .I0(ram[16124]), .I1(ram[16116]), .I2(ram[16108]), .I3(
        ram[16100]), .S0(n27220), .S1(n26745), .ZN(n24013) );
  MUX41 U9408 ( .I0(n23973), .I1(n23974), .I2(n23975), .I3(n23976), .S0(
        n26242), .S1(n26360), .ZN(n23972) );
  MUX41 U9409 ( .I0(ram[15004]), .I1(ram[14996]), .I2(ram[14988]), .I3(
        ram[14980]), .S0(n27217), .S1(n26742), .ZN(n23976) );
  MUX41 U9410 ( .I0(ram[15036]), .I1(ram[15028]), .I2(ram[15020]), .I3(
        ram[15012]), .S0(n27217), .S1(n26742), .ZN(n23974) );
  MUX41 U9411 ( .I0(ram[15100]), .I1(ram[15092]), .I2(ram[15084]), .I3(
        ram[15076]), .S0(n27217), .S1(n26742), .ZN(n23973) );
  MUX41 U9412 ( .I0(n23953), .I1(n23954), .I2(n23955), .I3(n23956), .S0(
        n26242), .S1(n26360), .ZN(n23952) );
  MUX41 U9413 ( .I0(ram[14524]), .I1(ram[14516]), .I2(ram[14508]), .I3(
        ram[14500]), .S0(n27216), .S1(n26741), .ZN(n23954) );
  MUX41 U9414 ( .I0(ram[14492]), .I1(ram[14484]), .I2(ram[14476]), .I3(
        ram[14468]), .S0(n27216), .S1(n26741), .ZN(n23956) );
  MUX41 U9415 ( .I0(ram[14588]), .I1(ram[14580]), .I2(ram[14572]), .I3(
        ram[14564]), .S0(n27216), .S1(n26741), .ZN(n23953) );
  MUX41 U9416 ( .I0(n23928), .I1(n23929), .I2(n23930), .I3(n23931), .S0(
        n26242), .S1(n26360), .ZN(n23927) );
  MUX41 U9417 ( .I0(ram[14012]), .I1(ram[14004]), .I2(ram[13996]), .I3(
        ram[13988]), .S0(n27215), .S1(n26740), .ZN(n23929) );
  MUX41 U9418 ( .I0(ram[13980]), .I1(ram[13972]), .I2(ram[13964]), .I3(
        ram[13956]), .S0(n27215), .S1(n26740), .ZN(n23931) );
  MUX41 U9419 ( .I0(ram[14076]), .I1(ram[14068]), .I2(ram[14060]), .I3(
        ram[14052]), .S0(n27215), .S1(n26740), .ZN(n23928) );
  MUX41 U9420 ( .I0(n23888), .I1(n23889), .I2(n23890), .I3(n23891), .S0(
        n26241), .S1(n26359), .ZN(n23887) );
  MUX41 U9421 ( .I0(ram[12956]), .I1(ram[12948]), .I2(ram[12940]), .I3(
        ram[12932]), .S0(n27212), .S1(n26737), .ZN(n23891) );
  MUX41 U9422 ( .I0(ram[12988]), .I1(ram[12980]), .I2(ram[12972]), .I3(
        ram[12964]), .S0(n27212), .S1(n26737), .ZN(n23889) );
  MUX41 U9423 ( .I0(ram[13052]), .I1(ram[13044]), .I2(ram[13036]), .I3(
        ram[13028]), .S0(n27212), .S1(n26737), .ZN(n23888) );
  MUX41 U9424 ( .I0(n23868), .I1(n23869), .I2(n23870), .I3(n23871), .S0(
        n26241), .S1(n26359), .ZN(n23867) );
  MUX41 U9425 ( .I0(ram[12476]), .I1(ram[12468]), .I2(ram[12460]), .I3(
        ram[12452]), .S0(n27211), .S1(n26736), .ZN(n23869) );
  MUX41 U9426 ( .I0(ram[12444]), .I1(ram[12436]), .I2(ram[12428]), .I3(
        ram[12420]), .S0(n27211), .S1(n26736), .ZN(n23871) );
  MUX41 U9427 ( .I0(ram[12540]), .I1(ram[12532]), .I2(ram[12524]), .I3(
        ram[12516]), .S0(n27211), .S1(n26736), .ZN(n23868) );
  MUX41 U9428 ( .I0(n23671), .I1(n23672), .I2(n23673), .I3(n23674), .S0(
        n26238), .S1(n26356), .ZN(n23670) );
  MUX41 U9429 ( .I0(ram[7868]), .I1(ram[7860]), .I2(ram[7852]), .I3(
        ram[7844]), .S0(n27200), .S1(n26725), .ZN(n23672) );
  MUX41 U9430 ( .I0(ram[7836]), .I1(ram[7828]), .I2(ram[7820]), .I3(
        ram[7812]), .S0(n27200), .S1(n26725), .ZN(n23674) );
  MUX41 U9431 ( .I0(ram[7932]), .I1(ram[7924]), .I2(ram[7916]), .I3(
        ram[7908]), .S0(n27200), .S1(n26725), .ZN(n23671) );
  MUX41 U9432 ( .I0(n23611), .I1(n23612), .I2(n23613), .I3(n23614), .S0(
        n26237), .S1(n26355), .ZN(n23610) );
  MUX41 U9433 ( .I0(ram[6332]), .I1(ram[6324]), .I2(ram[6316]), .I3(
        ram[6308]), .S0(n27196), .S1(n26721), .ZN(n23612) );
  MUX41 U9434 ( .I0(ram[6300]), .I1(ram[6292]), .I2(ram[6284]), .I3(
        ram[6276]), .S0(n27196), .S1(n26721), .ZN(n23614) );
  MUX41 U9435 ( .I0(ram[6396]), .I1(ram[6388]), .I2(ram[6380]), .I3(
        ram[6372]), .S0(n27196), .S1(n26721), .ZN(n23611) );
  MUX41 U9436 ( .I0(n23631), .I1(n23632), .I2(n23633), .I3(n23634), .S0(
        n26237), .S1(n26355), .ZN(n23630) );
  MUX41 U9437 ( .I0(ram[6844]), .I1(ram[6836]), .I2(ram[6828]), .I3(
        ram[6820]), .S0(n27197), .S1(n26722), .ZN(n23632) );
  MUX41 U9438 ( .I0(ram[6812]), .I1(ram[6804]), .I2(ram[6796]), .I3(
        ram[6788]), .S0(n27197), .S1(n26722), .ZN(n23634) );
  MUX41 U9439 ( .I0(ram[6908]), .I1(ram[6900]), .I2(ram[6892]), .I3(
        ram[6884]), .S0(n27198), .S1(n26723), .ZN(n23631) );
  MUX41 U9440 ( .I0(n23586), .I1(n23587), .I2(n23588), .I3(n23589), .S0(
        n26237), .S1(n26355), .ZN(n23585) );
  MUX41 U9441 ( .I0(ram[5820]), .I1(ram[5812]), .I2(ram[5804]), .I3(
        ram[5796]), .S0(n27195), .S1(n26720), .ZN(n23587) );
  MUX41 U9442 ( .I0(ram[5788]), .I1(ram[5780]), .I2(ram[5772]), .I3(
        ram[5764]), .S0(n27195), .S1(n26720), .ZN(n23589) );
  MUX41 U9443 ( .I0(ram[5884]), .I1(ram[5876]), .I2(ram[5868]), .I3(
        ram[5860]), .S0(n27195), .S1(n26720), .ZN(n23586) );
  MUX41 U9444 ( .I0(n23842), .I1(n23843), .I2(n23844), .I3(n23845), .S0(
        n26240), .S1(n26358), .ZN(n23841) );
  MUX41 U9445 ( .I0(ram[11964]), .I1(ram[11956]), .I2(ram[11948]), .I3(
        ram[11940]), .S0(n27210), .S1(n26735), .ZN(n23843) );
  MUX41 U9446 ( .I0(ram[11932]), .I1(ram[11924]), .I2(ram[11916]), .I3(
        ram[11908]), .S0(n27210), .S1(n26735), .ZN(n23845) );
  MUX41 U9447 ( .I0(ram[12028]), .I1(ram[12020]), .I2(ram[12012]), .I3(
        ram[12004]), .S0(n27210), .S1(n26735), .ZN(n23842) );
  MUX41 U9448 ( .I0(n23782), .I1(n23783), .I2(n23784), .I3(n23785), .S0(
        n26239), .S1(n26357), .ZN(n23781) );
  MUX41 U9449 ( .I0(ram[10428]), .I1(ram[10420]), .I2(ram[10412]), .I3(
        ram[10404]), .S0(n27206), .S1(n26731), .ZN(n23783) );
  MUX41 U9450 ( .I0(ram[10396]), .I1(ram[10388]), .I2(ram[10380]), .I3(
        ram[10372]), .S0(n27206), .S1(n26731), .ZN(n23785) );
  MUX41 U9451 ( .I0(ram[10492]), .I1(ram[10484]), .I2(ram[10476]), .I3(
        ram[10468]), .S0(n27206), .S1(n26731), .ZN(n23782) );
  MUX41 U9452 ( .I0(n23802), .I1(n23803), .I2(n23804), .I3(n23805), .S0(
        n26240), .S1(n26358), .ZN(n23801) );
  MUX41 U9453 ( .I0(ram[10940]), .I1(ram[10932]), .I2(ram[10924]), .I3(
        ram[10916]), .S0(n27207), .S1(n26732), .ZN(n23803) );
  MUX41 U9454 ( .I0(ram[10908]), .I1(ram[10900]), .I2(ram[10892]), .I3(
        ram[10884]), .S0(n27207), .S1(n26732), .ZN(n23805) );
  MUX41 U9455 ( .I0(ram[11004]), .I1(ram[10996]), .I2(ram[10988]), .I3(
        ram[10980]), .S0(n27207), .S1(n26732), .ZN(n23802) );
  MUX41 U9456 ( .I0(n23757), .I1(n23758), .I2(n23759), .I3(n23760), .S0(
        n26239), .S1(n26357), .ZN(n23756) );
  MUX41 U9457 ( .I0(ram[9916]), .I1(ram[9908]), .I2(ram[9900]), .I3(
        ram[9892]), .S0(n27205), .S1(n26730), .ZN(n23758) );
  MUX41 U9458 ( .I0(ram[9884]), .I1(ram[9876]), .I2(ram[9868]), .I3(
        ram[9860]), .S0(n27205), .S1(n26730), .ZN(n23760) );
  MUX41 U9459 ( .I0(ram[9980]), .I1(ram[9972]), .I2(ram[9964]), .I3(
        ram[9956]), .S0(n27205), .S1(n26730), .ZN(n23757) );
  MUX41 U9460 ( .I0(n23697), .I1(n23698), .I2(n23699), .I3(n23700), .S0(
        n26238), .S1(n26356), .ZN(n23696) );
  MUX41 U9461 ( .I0(ram[8380]), .I1(ram[8372]), .I2(ram[8364]), .I3(
        ram[8356]), .S0(n27201), .S1(n26726), .ZN(n23698) );
  MUX41 U9462 ( .I0(ram[8348]), .I1(ram[8340]), .I2(ram[8332]), .I3(
        ram[8324]), .S0(n27201), .S1(n26726), .ZN(n23700) );
  MUX41 U9463 ( .I0(ram[8444]), .I1(ram[8436]), .I2(ram[8428]), .I3(
        ram[8420]), .S0(n27201), .S1(n26726), .ZN(n23697) );
  MUX41 U9464 ( .I0(n24697), .I1(n24698), .I2(n24699), .I3(n24700), .S0(
        n26253), .S1(n26371), .ZN(n24696) );
  MUX41 U9465 ( .I0(ram[16061]), .I1(ram[16053]), .I2(ram[16045]), .I3(
        ram[16037]), .S0(n27259), .S1(n26784), .ZN(n24698) );
  MUX41 U9466 ( .I0(ram[16029]), .I1(ram[16021]), .I2(ram[16013]), .I3(
        ram[16005]), .S0(n27259), .S1(n26784), .ZN(n24700) );
  MUX41 U9467 ( .I0(ram[16125]), .I1(ram[16117]), .I2(ram[16109]), .I3(
        ram[16101]), .S0(n27259), .S1(n26784), .ZN(n24697) );
  MUX41 U9468 ( .I0(n24657), .I1(n24658), .I2(n24659), .I3(n24660), .S0(
        n26252), .S1(n26370), .ZN(n24656) );
  MUX41 U9469 ( .I0(ram[15005]), .I1(ram[14997]), .I2(ram[14989]), .I3(
        ram[14981]), .S0(n27256), .S1(n26781), .ZN(n24660) );
  MUX41 U9470 ( .I0(ram[15037]), .I1(ram[15029]), .I2(ram[15021]), .I3(
        ram[15013]), .S0(n27256), .S1(n26781), .ZN(n24658) );
  MUX41 U9471 ( .I0(ram[15101]), .I1(ram[15093]), .I2(ram[15085]), .I3(
        ram[15077]), .S0(n27257), .S1(n26782), .ZN(n24657) );
  MUX41 U9472 ( .I0(n24637), .I1(n24638), .I2(n24639), .I3(n24640), .S0(
        n26252), .S1(n26370), .ZN(n24636) );
  MUX41 U9473 ( .I0(ram[14525]), .I1(ram[14517]), .I2(ram[14509]), .I3(
        ram[14501]), .S0(n27255), .S1(n26780), .ZN(n24638) );
  MUX41 U9474 ( .I0(ram[14493]), .I1(ram[14485]), .I2(ram[14477]), .I3(
        ram[14469]), .S0(n27255), .S1(n26780), .ZN(n24640) );
  MUX41 U9475 ( .I0(ram[14589]), .I1(ram[14581]), .I2(ram[14573]), .I3(
        ram[14565]), .S0(n27255), .S1(n26780), .ZN(n24637) );
  MUX41 U9476 ( .I0(n24612), .I1(n24613), .I2(n24614), .I3(n24615), .S0(
        n26251), .S1(n26369), .ZN(n24611) );
  MUX41 U9477 ( .I0(ram[14013]), .I1(ram[14005]), .I2(ram[13997]), .I3(
        ram[13989]), .S0(n27254), .S1(n26779), .ZN(n24613) );
  MUX41 U9478 ( .I0(ram[13981]), .I1(ram[13973]), .I2(ram[13965]), .I3(
        ram[13957]), .S0(n27254), .S1(n26779), .ZN(n24615) );
  MUX41 U9479 ( .I0(ram[14077]), .I1(ram[14069]), .I2(ram[14061]), .I3(
        ram[14053]), .S0(n27254), .S1(n26779), .ZN(n24612) );
  MUX41 U9480 ( .I0(n24572), .I1(n24573), .I2(n24574), .I3(n24575), .S0(
        n26251), .S1(n26369), .ZN(n24571) );
  MUX41 U9481 ( .I0(ram[12957]), .I1(ram[12949]), .I2(ram[12941]), .I3(
        ram[12933]), .S0(n27251), .S1(n26776), .ZN(n24575) );
  MUX41 U9482 ( .I0(ram[12989]), .I1(ram[12981]), .I2(ram[12973]), .I3(
        ram[12965]), .S0(n27252), .S1(n26777), .ZN(n24573) );
  MUX41 U9483 ( .I0(ram[13053]), .I1(ram[13045]), .I2(ram[13037]), .I3(
        ram[13029]), .S0(n27252), .S1(n26777), .ZN(n24572) );
  MUX41 U9484 ( .I0(n24552), .I1(n24553), .I2(n24554), .I3(n24555), .S0(
        n26250), .S1(n26368), .ZN(n24551) );
  MUX41 U9485 ( .I0(ram[12477]), .I1(ram[12469]), .I2(ram[12461]), .I3(
        ram[12453]), .S0(n27250), .S1(n26775), .ZN(n24553) );
  MUX41 U9486 ( .I0(ram[12445]), .I1(ram[12437]), .I2(ram[12429]), .I3(
        ram[12421]), .S0(n27250), .S1(n26775), .ZN(n24555) );
  MUX41 U9487 ( .I0(ram[12541]), .I1(ram[12533]), .I2(ram[12525]), .I3(
        ram[12517]), .S0(n27250), .S1(n26775), .ZN(n24552) );
  MUX41 U9488 ( .I0(n24355), .I1(n24356), .I2(n24357), .I3(n24358), .S0(
        n26248), .S1(n26366), .ZN(n24354) );
  MUX41 U9489 ( .I0(ram[7869]), .I1(ram[7861]), .I2(ram[7853]), .I3(
        ram[7845]), .S0(n27239), .S1(n26764), .ZN(n24356) );
  MUX41 U9490 ( .I0(ram[7837]), .I1(ram[7829]), .I2(ram[7821]), .I3(
        ram[7813]), .S0(n27239), .S1(n26764), .ZN(n24358) );
  MUX41 U9491 ( .I0(ram[7933]), .I1(ram[7925]), .I2(ram[7917]), .I3(
        ram[7909]), .S0(n27239), .S1(n26764), .ZN(n24355) );
  MUX41 U9492 ( .I0(n24295), .I1(n24296), .I2(n24297), .I3(n24298), .S0(
        n26247), .S1(n26365), .ZN(n24294) );
  MUX41 U9493 ( .I0(ram[6333]), .I1(ram[6325]), .I2(ram[6317]), .I3(
        ram[6309]), .S0(n27236), .S1(n26761), .ZN(n24296) );
  MUX41 U9494 ( .I0(ram[6301]), .I1(ram[6293]), .I2(ram[6285]), .I3(
        ram[6277]), .S0(n27235), .S1(n26760), .ZN(n24298) );
  MUX41 U9495 ( .I0(ram[6397]), .I1(ram[6389]), .I2(ram[6381]), .I3(
        ram[6373]), .S0(n27236), .S1(n26761), .ZN(n24295) );
  MUX41 U9496 ( .I0(n24315), .I1(n24316), .I2(n24317), .I3(n24318), .S0(
        n26247), .S1(n26365), .ZN(n24314) );
  MUX41 U9497 ( .I0(ram[6845]), .I1(ram[6837]), .I2(ram[6829]), .I3(
        ram[6821]), .S0(n27237), .S1(n26762), .ZN(n24316) );
  MUX41 U9498 ( .I0(ram[6813]), .I1(ram[6805]), .I2(ram[6797]), .I3(
        ram[6789]), .S0(n27237), .S1(n26762), .ZN(n24318) );
  MUX41 U9499 ( .I0(ram[6909]), .I1(ram[6901]), .I2(ram[6893]), .I3(
        ram[6885]), .S0(n27237), .S1(n26762), .ZN(n24315) );
  MUX41 U9500 ( .I0(n24270), .I1(n24271), .I2(n24272), .I3(n24273), .S0(
        n26246), .S1(n26364), .ZN(n24269) );
  MUX41 U9501 ( .I0(ram[5821]), .I1(ram[5813]), .I2(ram[5805]), .I3(
        ram[5797]), .S0(n27234), .S1(n26759), .ZN(n24271) );
  MUX41 U9502 ( .I0(ram[5789]), .I1(ram[5781]), .I2(ram[5773]), .I3(
        ram[5765]), .S0(n27234), .S1(n26759), .ZN(n24273) );
  MUX41 U9503 ( .I0(ram[5885]), .I1(ram[5877]), .I2(ram[5869]), .I3(
        ram[5861]), .S0(n27234), .S1(n26759), .ZN(n24270) );
  MUX41 U9504 ( .I0(n24526), .I1(n24527), .I2(n24528), .I3(n24529), .S0(
        n26250), .S1(n26368), .ZN(n24525) );
  MUX41 U9505 ( .I0(ram[11965]), .I1(ram[11957]), .I2(ram[11949]), .I3(
        ram[11941]), .S0(n27249), .S1(n26774), .ZN(n24527) );
  MUX41 U9506 ( .I0(ram[11933]), .I1(ram[11925]), .I2(ram[11917]), .I3(
        ram[11909]), .S0(n27249), .S1(n26774), .ZN(n24529) );
  MUX41 U9507 ( .I0(ram[12029]), .I1(ram[12021]), .I2(ram[12013]), .I3(
        ram[12005]), .S0(n27249), .S1(n26774), .ZN(n24526) );
  MUX41 U9508 ( .I0(n24466), .I1(n24467), .I2(n24468), .I3(n24469), .S0(
        n26249), .S1(n26367), .ZN(n24465) );
  MUX41 U9509 ( .I0(ram[10429]), .I1(ram[10421]), .I2(ram[10413]), .I3(
        ram[10405]), .S0(n27245), .S1(n26770), .ZN(n24467) );
  MUX41 U9510 ( .I0(ram[10397]), .I1(ram[10389]), .I2(ram[10381]), .I3(
        ram[10373]), .S0(n27245), .S1(n26770), .ZN(n24469) );
  MUX41 U9511 ( .I0(ram[10493]), .I1(ram[10485]), .I2(ram[10477]), .I3(
        ram[10469]), .S0(n27246), .S1(n26771), .ZN(n24466) );
  MUX41 U9512 ( .I0(n24486), .I1(n24487), .I2(n24488), .I3(n24489), .S0(
        n26250), .S1(n26368), .ZN(n24485) );
  MUX41 U9513 ( .I0(ram[10941]), .I1(ram[10933]), .I2(ram[10925]), .I3(
        ram[10917]), .S0(n27247), .S1(n26772), .ZN(n24487) );
  MUX41 U9514 ( .I0(ram[10909]), .I1(ram[10901]), .I2(ram[10893]), .I3(
        ram[10885]), .S0(n27247), .S1(n26772), .ZN(n24489) );
  MUX41 U9515 ( .I0(ram[11005]), .I1(ram[10997]), .I2(ram[10989]), .I3(
        ram[10981]), .S0(n27247), .S1(n26772), .ZN(n24486) );
  MUX41 U9516 ( .I0(n24441), .I1(n24442), .I2(n24443), .I3(n24444), .S0(
        n26249), .S1(n26367), .ZN(n24440) );
  MUX41 U9517 ( .I0(ram[9917]), .I1(ram[9909]), .I2(ram[9901]), .I3(
        ram[9893]), .S0(n27244), .S1(n26769), .ZN(n24442) );
  MUX41 U9518 ( .I0(ram[9885]), .I1(ram[9877]), .I2(ram[9869]), .I3(
        ram[9861]), .S0(n27244), .S1(n26769), .ZN(n24444) );
  MUX41 U9519 ( .I0(ram[9981]), .I1(ram[9973]), .I2(ram[9965]), .I3(
        ram[9957]), .S0(n27244), .S1(n26769), .ZN(n24441) );
  MUX41 U9520 ( .I0(n24381), .I1(n24382), .I2(n24383), .I3(n24384), .S0(
        n26248), .S1(n26366), .ZN(n24380) );
  MUX41 U9521 ( .I0(ram[8381]), .I1(ram[8373]), .I2(ram[8365]), .I3(
        ram[8357]), .S0(n27240), .S1(n26765), .ZN(n24382) );
  MUX41 U9522 ( .I0(ram[8349]), .I1(ram[8341]), .I2(ram[8333]), .I3(
        ram[8325]), .S0(n27240), .S1(n26765), .ZN(n24384) );
  MUX41 U9523 ( .I0(ram[8445]), .I1(ram[8437]), .I2(ram[8429]), .I3(
        ram[8421]), .S0(n27241), .S1(n26766), .ZN(n24381) );
  MUX41 U9524 ( .I0(n25381), .I1(n25382), .I2(n25383), .I3(n25384), .S0(
        n26262), .S1(n26380), .ZN(n25380) );
  MUX41 U9525 ( .I0(ram[16062]), .I1(ram[16054]), .I2(ram[16046]), .I3(
        ram[16038]), .S0(n27298), .S1(n26823), .ZN(n25382) );
  MUX41 U9526 ( .I0(ram[16030]), .I1(ram[16022]), .I2(ram[16014]), .I3(
        ram[16006]), .S0(n27298), .S1(n26823), .ZN(n25384) );
  MUX41 U9527 ( .I0(ram[16126]), .I1(ram[16118]), .I2(ram[16110]), .I3(
        ram[16102]), .S0(n27298), .S1(n26823), .ZN(n25381) );
  MUX41 U9528 ( .I0(n25341), .I1(n25342), .I2(n25343), .I3(n25344), .S0(
        n26262), .S1(n26380), .ZN(n25340) );
  MUX41 U9529 ( .I0(ram[15006]), .I1(ram[14998]), .I2(ram[14990]), .I3(
        ram[14982]), .S0(n27296), .S1(n26821), .ZN(n25344) );
  MUX41 U9530 ( .I0(ram[15038]), .I1(ram[15030]), .I2(ram[15022]), .I3(
        ram[15014]), .S0(n27296), .S1(n26821), .ZN(n25342) );
  MUX41 U9531 ( .I0(ram[15102]), .I1(ram[15094]), .I2(ram[15086]), .I3(
        ram[15078]), .S0(n27296), .S1(n26821), .ZN(n25341) );
  MUX41 U9532 ( .I0(n25321), .I1(n25322), .I2(n25323), .I3(n25324), .S0(
        n26262), .S1(n26380), .ZN(n25320) );
  MUX41 U9533 ( .I0(ram[14526]), .I1(ram[14518]), .I2(ram[14510]), .I3(
        ram[14502]), .S0(n27295), .S1(n26820), .ZN(n25322) );
  MUX41 U9534 ( .I0(ram[14494]), .I1(ram[14486]), .I2(ram[14478]), .I3(
        ram[14470]), .S0(n27295), .S1(n26820), .ZN(n25324) );
  MUX41 U9535 ( .I0(ram[14590]), .I1(ram[14582]), .I2(ram[14574]), .I3(
        ram[14566]), .S0(n27295), .S1(n26820), .ZN(n25321) );
  MUX41 U9536 ( .I0(n25296), .I1(n25297), .I2(n25298), .I3(n25299), .S0(
        n26261), .S1(n26379), .ZN(n25295) );
  MUX41 U9537 ( .I0(ram[14014]), .I1(ram[14006]), .I2(ram[13998]), .I3(
        ram[13990]), .S0(n27293), .S1(n26818), .ZN(n25297) );
  MUX41 U9538 ( .I0(ram[13982]), .I1(ram[13974]), .I2(ram[13966]), .I3(
        ram[13958]), .S0(n27293), .S1(n26818), .ZN(n25299) );
  MUX41 U9539 ( .I0(ram[14078]), .I1(ram[14070]), .I2(ram[14062]), .I3(
        ram[14054]), .S0(n27294), .S1(n26819), .ZN(n25296) );
  MUX41 U9540 ( .I0(n25256), .I1(n25257), .I2(n25258), .I3(n25259), .S0(
        n26261), .S1(n26379), .ZN(n25255) );
  MUX41 U9541 ( .I0(ram[12958]), .I1(ram[12950]), .I2(ram[12942]), .I3(
        ram[12934]), .S0(n27291), .S1(n26816), .ZN(n25259) );
  MUX41 U9542 ( .I0(ram[12990]), .I1(ram[12982]), .I2(ram[12974]), .I3(
        ram[12966]), .S0(n27291), .S1(n26816), .ZN(n25257) );
  MUX41 U9543 ( .I0(ram[13054]), .I1(ram[13046]), .I2(ram[13038]), .I3(
        ram[13030]), .S0(n27291), .S1(n26816), .ZN(n25256) );
  MUX41 U9544 ( .I0(n25236), .I1(n25237), .I2(n25238), .I3(n25239), .S0(
        n26260), .S1(n26378), .ZN(n25235) );
  MUX41 U9545 ( .I0(ram[12478]), .I1(ram[12470]), .I2(ram[12462]), .I3(
        ram[12454]), .S0(n27290), .S1(n26815), .ZN(n25237) );
  MUX41 U9546 ( .I0(ram[12446]), .I1(ram[12438]), .I2(ram[12430]), .I3(
        ram[12422]), .S0(n27290), .S1(n26815), .ZN(n25239) );
  MUX41 U9547 ( .I0(ram[12542]), .I1(ram[12534]), .I2(ram[12526]), .I3(
        ram[12518]), .S0(n27290), .S1(n26815), .ZN(n25236) );
  MUX41 U9548 ( .I0(n25039), .I1(n25040), .I2(n25041), .I3(n25042), .S0(
        n26258), .S1(n26376), .ZN(n25038) );
  MUX41 U9549 ( .I0(ram[7870]), .I1(ram[7862]), .I2(ram[7854]), .I3(
        ram[7846]), .S0(n27279), .S1(n26804), .ZN(n25040) );
  MUX41 U9550 ( .I0(ram[7838]), .I1(ram[7830]), .I2(ram[7822]), .I3(
        ram[7814]), .S0(n27279), .S1(n26804), .ZN(n25042) );
  MUX41 U9551 ( .I0(ram[7934]), .I1(ram[7926]), .I2(ram[7918]), .I3(
        ram[7910]), .S0(n27279), .S1(n26804), .ZN(n25039) );
  MUX41 U9552 ( .I0(n24979), .I1(n24980), .I2(n24981), .I3(n24982), .S0(
        n26257), .S1(n26375), .ZN(n24978) );
  MUX41 U9553 ( .I0(ram[6334]), .I1(ram[6326]), .I2(ram[6318]), .I3(
        ram[6310]), .S0(n27275), .S1(n26800), .ZN(n24980) );
  MUX41 U9554 ( .I0(ram[6302]), .I1(ram[6294]), .I2(ram[6286]), .I3(
        ram[6278]), .S0(n27275), .S1(n26800), .ZN(n24982) );
  MUX41 U9555 ( .I0(ram[6398]), .I1(ram[6390]), .I2(ram[6382]), .I3(
        ram[6374]), .S0(n27275), .S1(n26800), .ZN(n24979) );
  MUX41 U9556 ( .I0(n24999), .I1(n25000), .I2(n25001), .I3(n25002), .S0(
        n26257), .S1(n26375), .ZN(n24998) );
  MUX41 U9557 ( .I0(ram[6846]), .I1(ram[6838]), .I2(ram[6830]), .I3(
        ram[6822]), .S0(n27276), .S1(n26801), .ZN(n25000) );
  MUX41 U9558 ( .I0(ram[6814]), .I1(ram[6806]), .I2(ram[6798]), .I3(
        ram[6790]), .S0(n27276), .S1(n26801), .ZN(n25002) );
  MUX41 U9559 ( .I0(ram[6910]), .I1(ram[6902]), .I2(ram[6894]), .I3(
        ram[6886]), .S0(n27276), .S1(n26801), .ZN(n24999) );
  MUX41 U9560 ( .I0(n24954), .I1(n24955), .I2(n24956), .I3(n24957), .S0(
        n26256), .S1(n26374), .ZN(n24953) );
  MUX41 U9561 ( .I0(ram[5822]), .I1(ram[5814]), .I2(ram[5806]), .I3(
        ram[5798]), .S0(n27274), .S1(n26799), .ZN(n24955) );
  MUX41 U9562 ( .I0(ram[5790]), .I1(ram[5782]), .I2(ram[5774]), .I3(
        ram[5766]), .S0(n27274), .S1(n26799), .ZN(n24957) );
  MUX41 U9563 ( .I0(ram[5886]), .I1(ram[5878]), .I2(ram[5870]), .I3(
        ram[5862]), .S0(n27274), .S1(n26799), .ZN(n24954) );
  MUX41 U9564 ( .I0(n25210), .I1(n25211), .I2(n25212), .I3(n25213), .S0(
        n26260), .S1(n26378), .ZN(n25209) );
  MUX41 U9565 ( .I0(ram[11966]), .I1(ram[11958]), .I2(ram[11950]), .I3(
        ram[11942]), .S0(n27288), .S1(n26813), .ZN(n25211) );
  MUX41 U9566 ( .I0(ram[11934]), .I1(ram[11926]), .I2(ram[11918]), .I3(
        ram[11910]), .S0(n27288), .S1(n26813), .ZN(n25213) );
  MUX41 U9567 ( .I0(ram[12030]), .I1(ram[12022]), .I2(ram[12014]), .I3(
        ram[12006]), .S0(n27289), .S1(n26814), .ZN(n25210) );
  MUX41 U9568 ( .I0(n25150), .I1(n25151), .I2(n25152), .I3(n25153), .S0(
        n26259), .S1(n26377), .ZN(n25149) );
  MUX41 U9569 ( .I0(ram[10430]), .I1(ram[10422]), .I2(ram[10414]), .I3(
        ram[10406]), .S0(n27285), .S1(n26810), .ZN(n25151) );
  MUX41 U9570 ( .I0(ram[10398]), .I1(ram[10390]), .I2(ram[10382]), .I3(
        ram[10374]), .S0(n27285), .S1(n26810), .ZN(n25153) );
  MUX41 U9571 ( .I0(ram[10494]), .I1(ram[10486]), .I2(ram[10478]), .I3(
        ram[10470]), .S0(n27285), .S1(n26810), .ZN(n25150) );
  MUX41 U9572 ( .I0(n25170), .I1(n25171), .I2(n25172), .I3(n25173), .S0(
        n26259), .S1(n26377), .ZN(n25169) );
  MUX41 U9573 ( .I0(ram[10942]), .I1(ram[10934]), .I2(ram[10926]), .I3(
        ram[10918]), .S0(n27286), .S1(n26811), .ZN(n25171) );
  MUX41 U9574 ( .I0(ram[10910]), .I1(ram[10902]), .I2(ram[10894]), .I3(
        ram[10886]), .S0(n27286), .S1(n26811), .ZN(n25173) );
  MUX41 U9575 ( .I0(ram[11006]), .I1(ram[10998]), .I2(ram[10990]), .I3(
        ram[10982]), .S0(n27286), .S1(n26811), .ZN(n25170) );
  MUX41 U9576 ( .I0(n25125), .I1(n25126), .I2(n25127), .I3(n25128), .S0(
        n26259), .S1(n26377), .ZN(n25124) );
  MUX41 U9577 ( .I0(ram[9918]), .I1(ram[9910]), .I2(ram[9902]), .I3(
        ram[9894]), .S0(n27284), .S1(n26809), .ZN(n25126) );
  MUX41 U9578 ( .I0(ram[9886]), .I1(ram[9878]), .I2(ram[9870]), .I3(
        ram[9862]), .S0(n27283), .S1(n26808), .ZN(n25128) );
  MUX41 U9579 ( .I0(ram[9982]), .I1(ram[9974]), .I2(ram[9966]), .I3(
        ram[9958]), .S0(n27284), .S1(n26809), .ZN(n25125) );
  MUX41 U9580 ( .I0(n25065), .I1(n25066), .I2(n25067), .I3(n25068), .S0(
        n26258), .S1(n26376), .ZN(n25064) );
  MUX41 U9581 ( .I0(ram[8382]), .I1(ram[8374]), .I2(ram[8366]), .I3(
        ram[8358]), .S0(n27280), .S1(n26805), .ZN(n25066) );
  MUX41 U9582 ( .I0(ram[8350]), .I1(ram[8342]), .I2(ram[8334]), .I3(
        ram[8326]), .S0(n27280), .S1(n26805), .ZN(n25068) );
  MUX41 U9583 ( .I0(ram[8446]), .I1(ram[8438]), .I2(ram[8430]), .I3(
        ram[8422]), .S0(n27280), .S1(n26805), .ZN(n25065) );
  MUX41 U9584 ( .I0(n26065), .I1(n26066), .I2(n26067), .I3(n26068), .S0(
        n26272), .S1(n26390), .ZN(n26064) );
  MUX41 U9585 ( .I0(ram[16063]), .I1(ram[16055]), .I2(ram[16047]), .I3(
        ram[16039]), .S0(n27338), .S1(n26863), .ZN(n26066) );
  MUX41 U9586 ( .I0(ram[16031]), .I1(ram[16023]), .I2(ram[16015]), .I3(
        ram[16007]), .S0(n27338), .S1(n26863), .ZN(n26068) );
  MUX41 U9587 ( .I0(ram[16127]), .I1(ram[16119]), .I2(ram[16111]), .I3(
        ram[16103]), .S0(n27338), .S1(n26863), .ZN(n26065) );
  MUX41 U9588 ( .I0(n26025), .I1(n26026), .I2(n26027), .I3(n26028), .S0(
        n26272), .S1(n26390), .ZN(n26024) );
  MUX41 U9589 ( .I0(ram[15007]), .I1(ram[14999]), .I2(ram[14991]), .I3(
        ram[14983]), .S0(n27335), .S1(n26860), .ZN(n26028) );
  MUX41 U9590 ( .I0(ram[15039]), .I1(ram[15031]), .I2(ram[15023]), .I3(
        ram[15015]), .S0(n27335), .S1(n26860), .ZN(n26026) );
  MUX41 U9591 ( .I0(ram[15103]), .I1(ram[15095]), .I2(ram[15087]), .I3(
        ram[15079]), .S0(n27335), .S1(n26860), .ZN(n26025) );
  MUX41 U9592 ( .I0(n26005), .I1(n26006), .I2(n26007), .I3(n26008), .S0(
        n26271), .S1(n26389), .ZN(n26004) );
  MUX41 U9593 ( .I0(ram[14527]), .I1(ram[14519]), .I2(ram[14511]), .I3(
        ram[14503]), .S0(n27334), .S1(n26859), .ZN(n26006) );
  MUX41 U9594 ( .I0(ram[14495]), .I1(ram[14487]), .I2(ram[14479]), .I3(
        ram[14471]), .S0(n27334), .S1(n26859), .ZN(n26008) );
  MUX41 U9595 ( .I0(ram[14591]), .I1(ram[14583]), .I2(ram[14575]), .I3(
        ram[14567]), .S0(n27334), .S1(n26859), .ZN(n26005) );
  MUX41 U9596 ( .I0(n25980), .I1(n25981), .I2(n25982), .I3(n25983), .S0(
        n26271), .S1(n26389), .ZN(n25979) );
  MUX41 U9597 ( .I0(ram[14015]), .I1(ram[14007]), .I2(ram[13999]), .I3(
        ram[13991]), .S0(n27333), .S1(n26858), .ZN(n25981) );
  MUX41 U9598 ( .I0(ram[13983]), .I1(ram[13975]), .I2(ram[13967]), .I3(
        ram[13959]), .S0(n27333), .S1(n26858), .ZN(n25983) );
  MUX41 U9599 ( .I0(ram[14079]), .I1(ram[14071]), .I2(ram[14063]), .I3(
        ram[14055]), .S0(n27333), .S1(n26858), .ZN(n25980) );
  MUX41 U9600 ( .I0(n25940), .I1(n25941), .I2(n25942), .I3(n25943), .S0(
        n26270), .S1(n26388), .ZN(n25939) );
  MUX41 U9601 ( .I0(ram[12959]), .I1(ram[12951]), .I2(ram[12943]), .I3(
        ram[12935]), .S0(n27330), .S1(n26855), .ZN(n25943) );
  MUX41 U9602 ( .I0(ram[12991]), .I1(ram[12983]), .I2(ram[12975]), .I3(
        ram[12967]), .S0(n27330), .S1(n26855), .ZN(n25941) );
  MUX41 U9603 ( .I0(ram[13055]), .I1(ram[13047]), .I2(ram[13039]), .I3(
        ram[13031]), .S0(n27330), .S1(n26855), .ZN(n25940) );
  MUX41 U9604 ( .I0(n25920), .I1(n25921), .I2(n25922), .I3(n25923), .S0(
        n26270), .S1(n26388), .ZN(n25919) );
  MUX41 U9605 ( .I0(ram[12479]), .I1(ram[12471]), .I2(ram[12463]), .I3(
        ram[12455]), .S0(n27329), .S1(n26854), .ZN(n25921) );
  MUX41 U9606 ( .I0(ram[12447]), .I1(ram[12439]), .I2(ram[12431]), .I3(
        ram[12423]), .S0(n27329), .S1(n26854), .ZN(n25923) );
  MUX41 U9607 ( .I0(ram[12543]), .I1(ram[12535]), .I2(ram[12527]), .I3(
        ram[12519]), .S0(n27329), .S1(n26854), .ZN(n25920) );
  MUX41 U9608 ( .I0(n25723), .I1(n25724), .I2(n25725), .I3(n25726), .S0(
        n26267), .S1(n26385), .ZN(n25722) );
  MUX41 U9609 ( .I0(ram[7871]), .I1(ram[7863]), .I2(ram[7855]), .I3(
        ram[7847]), .S0(n27318), .S1(n26843), .ZN(n25724) );
  MUX41 U9610 ( .I0(ram[7839]), .I1(ram[7831]), .I2(ram[7823]), .I3(
        ram[7815]), .S0(n27318), .S1(n26843), .ZN(n25726) );
  MUX41 U9611 ( .I0(ram[7935]), .I1(ram[7927]), .I2(ram[7919]), .I3(
        ram[7911]), .S0(n27318), .S1(n26843), .ZN(n25723) );
  MUX41 U9612 ( .I0(n25663), .I1(n25664), .I2(n25665), .I3(n25666), .S0(
        n26266), .S1(n26384), .ZN(n25662) );
  MUX41 U9613 ( .I0(ram[6335]), .I1(ram[6327]), .I2(ram[6319]), .I3(
        ram[6311]), .S0(n27314), .S1(n26839), .ZN(n25664) );
  MUX41 U9614 ( .I0(ram[6303]), .I1(ram[6295]), .I2(ram[6287]), .I3(
        ram[6279]), .S0(n27314), .S1(n26839), .ZN(n25666) );
  MUX41 U9615 ( .I0(ram[6399]), .I1(ram[6391]), .I2(ram[6383]), .I3(
        ram[6375]), .S0(n27314), .S1(n26839), .ZN(n25663) );
  MUX41 U9616 ( .I0(n25683), .I1(n25684), .I2(n25685), .I3(n25686), .S0(
        n26267), .S1(n26385), .ZN(n25682) );
  MUX41 U9617 ( .I0(ram[6847]), .I1(ram[6839]), .I2(ram[6831]), .I3(
        ram[6823]), .S0(n27316), .S1(n26841), .ZN(n25684) );
  MUX41 U9618 ( .I0(ram[6815]), .I1(ram[6807]), .I2(ram[6799]), .I3(
        ram[6791]), .S0(n27315), .S1(n26840), .ZN(n25686) );
  MUX41 U9619 ( .I0(ram[6911]), .I1(ram[6903]), .I2(ram[6895]), .I3(
        ram[6887]), .S0(n27316), .S1(n26841), .ZN(n25683) );
  MUX41 U9620 ( .I0(n25638), .I1(n25639), .I2(n25640), .I3(n25641), .S0(
        n26266), .S1(n26384), .ZN(n25637) );
  MUX41 U9621 ( .I0(ram[5823]), .I1(ram[5815]), .I2(ram[5807]), .I3(
        ram[5799]), .S0(n27313), .S1(n26838), .ZN(n25639) );
  MUX41 U9622 ( .I0(ram[5791]), .I1(ram[5783]), .I2(ram[5775]), .I3(
        ram[5767]), .S0(n27313), .S1(n26838), .ZN(n25641) );
  MUX41 U9623 ( .I0(ram[5887]), .I1(ram[5879]), .I2(ram[5871]), .I3(
        ram[5863]), .S0(n27313), .S1(n26838), .ZN(n25638) );
  MUX41 U9624 ( .I0(n25894), .I1(n25895), .I2(n25896), .I3(n25897), .S0(
        n26270), .S1(n26388), .ZN(n25893) );
  MUX41 U9625 ( .I0(ram[11967]), .I1(ram[11959]), .I2(ram[11951]), .I3(
        ram[11943]), .S0(n27328), .S1(n26853), .ZN(n25895) );
  MUX41 U9626 ( .I0(ram[11935]), .I1(ram[11927]), .I2(ram[11919]), .I3(
        ram[11911]), .S0(n27328), .S1(n26853), .ZN(n25897) );
  MUX41 U9627 ( .I0(ram[12031]), .I1(ram[12023]), .I2(ram[12015]), .I3(
        ram[12007]), .S0(n27328), .S1(n26853), .ZN(n25894) );
  MUX41 U9628 ( .I0(n25834), .I1(n25835), .I2(n25836), .I3(n25837), .S0(
        n26269), .S1(n26387), .ZN(n25833) );
  MUX41 U9629 ( .I0(ram[10431]), .I1(ram[10423]), .I2(ram[10415]), .I3(
        ram[10407]), .S0(n27324), .S1(n26849), .ZN(n25835) );
  MUX41 U9630 ( .I0(ram[10399]), .I1(ram[10391]), .I2(ram[10383]), .I3(
        ram[10375]), .S0(n27324), .S1(n26849), .ZN(n25837) );
  MUX41 U9631 ( .I0(ram[10495]), .I1(ram[10487]), .I2(ram[10479]), .I3(
        ram[10471]), .S0(n27324), .S1(n26849), .ZN(n25834) );
  MUX41 U9632 ( .I0(n25854), .I1(n25855), .I2(n25856), .I3(n25857), .S0(
        n26269), .S1(n26387), .ZN(n25853) );
  MUX41 U9633 ( .I0(ram[10943]), .I1(ram[10935]), .I2(ram[10927]), .I3(
        ram[10919]), .S0(n27325), .S1(n26850), .ZN(n25855) );
  MUX41 U9634 ( .I0(ram[10911]), .I1(ram[10903]), .I2(ram[10895]), .I3(
        ram[10887]), .S0(n27325), .S1(n26850), .ZN(n25857) );
  MUX41 U9635 ( .I0(ram[11007]), .I1(ram[10999]), .I2(ram[10991]), .I3(
        ram[10983]), .S0(n27326), .S1(n26851), .ZN(n25854) );
  MUX41 U9636 ( .I0(n25809), .I1(n25810), .I2(n25811), .I3(n25812), .S0(
        n26269), .S1(n26387), .ZN(n25808) );
  MUX41 U9637 ( .I0(ram[9919]), .I1(ram[9911]), .I2(ram[9903]), .I3(
        ram[9895]), .S0(n27323), .S1(n26848), .ZN(n25810) );
  MUX41 U9638 ( .I0(ram[9887]), .I1(ram[9879]), .I2(ram[9871]), .I3(
        ram[9863]), .S0(n27323), .S1(n26848), .ZN(n25812) );
  MUX41 U9639 ( .I0(ram[9983]), .I1(ram[9975]), .I2(ram[9967]), .I3(
        ram[9959]), .S0(n27323), .S1(n26848), .ZN(n25809) );
  MUX41 U9640 ( .I0(n25749), .I1(n25750), .I2(n25751), .I3(n25752), .S0(
        n26268), .S1(n26386), .ZN(n25748) );
  MUX41 U9641 ( .I0(ram[8383]), .I1(ram[8375]), .I2(ram[8367]), .I3(
        ram[8359]), .S0(n27319), .S1(n26844), .ZN(n25750) );
  MUX41 U9642 ( .I0(ram[8351]), .I1(ram[8343]), .I2(ram[8335]), .I3(
        ram[8327]), .S0(n27319), .S1(n26844), .ZN(n25752) );
  MUX41 U9643 ( .I0(ram[8447]), .I1(ram[8439]), .I2(ram[8431]), .I3(
        ram[8423]), .S0(n27319), .S1(n26844), .ZN(n25749) );
  MUX41 U9644 ( .I0(n4098), .I1(n20625), .I2(n20626), .I3(n20627), .S0(
        n26194), .S1(n26312), .ZN(n3969) );
  MUX41 U9645 ( .I0(ram[280]), .I1(ram[272]), .I2(ram[264]), .I3(ram[256]), .S0(n27024), .S1(n26549), .ZN(n20627) );
  MUX41 U9646 ( .I0(ram[312]), .I1(ram[304]), .I2(ram[296]), .I3(ram[288]), .S0(n27024), .S1(n26549), .ZN(n20625) );
  MUX41 U9647 ( .I0(ram[376]), .I1(ram[368]), .I2(ram[360]), .I3(ram[352]), .S0(n27024), .S1(n26549), .ZN(n4098) );
  MUX41 U9648 ( .I0(n20644), .I1(n20645), .I2(n20646), .I3(n20647), .S0(
        n26194), .S1(n26312), .ZN(n20643) );
  MUX41 U9649 ( .I0(ram[792]), .I1(ram[784]), .I2(ram[776]), .I3(ram[768]), .S0(n27025), .S1(n26550), .ZN(n20647) );
  MUX41 U9650 ( .I0(ram[824]), .I1(ram[816]), .I2(ram[808]), .I3(ram[800]), .S0(n27025), .S1(n26550), .ZN(n20645) );
  MUX41 U9651 ( .I0(ram[888]), .I1(ram[880]), .I2(ram[872]), .I3(ram[864]), .S0(n27026), .S1(n26551), .ZN(n20644) );
  MUX41 U9652 ( .I0(ram[3416]), .I1(ram[3408]), .I2(ram[3400]), .I3(
        ram[3392]), .S0(n27032), .S1(n26557), .ZN(n20751) );
  MUX41 U9653 ( .I0(ram[3544]), .I1(ram[3536]), .I2(ram[3528]), .I3(
        ram[3520]), .S0(n27032), .S1(n26557), .ZN(n20756) );
  MUX41 U9654 ( .I0(ram[3288]), .I1(ram[3280]), .I2(ram[3272]), .I3(
        ram[3264]), .S0(n27031), .S1(n26556), .ZN(n20746) );
  MUX41 U9655 ( .I0(ram[3160]), .I1(ram[3152]), .I2(ram[3144]), .I3(
        ram[3136]), .S0(n27031), .S1(n26556), .ZN(n20741) );
  MUX41 U9656 ( .I0(ram[3928]), .I1(ram[3920]), .I2(ram[3912]), .I3(
        ram[3904]), .S0(n27033), .S1(n26558), .ZN(n20771) );
  MUX41 U9657 ( .I0(ram[4056]), .I1(ram[4048]), .I2(ram[4040]), .I3(
        ram[4032]), .S0(n27033), .S1(n26558), .ZN(n20776) );
  MUX41 U9658 ( .I0(ram[3800]), .I1(ram[3792]), .I2(ram[3784]), .I3(
        ram[3776]), .S0(n27033), .S1(n26558), .ZN(n20766) );
  MUX41 U9659 ( .I0(ram[3672]), .I1(ram[3664]), .I2(ram[3656]), .I3(
        ram[3648]), .S0(n27032), .S1(n26557), .ZN(n20761) );
  MUX41 U9660 ( .I0(ram[2392]), .I1(ram[2384]), .I2(ram[2376]), .I3(
        ram[2368]), .S0(n27029), .S1(n26554), .ZN(n20711) );
  MUX41 U9661 ( .I0(ram[2520]), .I1(ram[2512]), .I2(ram[2504]), .I3(
        ram[2496]), .S0(n27029), .S1(n26554), .ZN(n20716) );
  MUX41 U9662 ( .I0(ram[2264]), .I1(ram[2256]), .I2(ram[2248]), .I3(
        ram[2240]), .S0(n27029), .S1(n26554), .ZN(n20706) );
  MUX41 U9663 ( .I0(ram[2136]), .I1(ram[2128]), .I2(ram[2120]), .I3(
        ram[2112]), .S0(n27029), .S1(n26554), .ZN(n20701) );
  MUX41 U9664 ( .I0(ram[2904]), .I1(ram[2896]), .I2(ram[2888]), .I3(
        ram[2880]), .S0(n27030), .S1(n26555), .ZN(n20731) );
  MUX41 U9665 ( .I0(ram[3032]), .I1(ram[3024]), .I2(ram[3016]), .I3(
        ram[3008]), .S0(n27031), .S1(n26556), .ZN(n20736) );
  MUX41 U9666 ( .I0(ram[2776]), .I1(ram[2768]), .I2(ram[2760]), .I3(
        ram[2752]), .S0(n27030), .S1(n26555), .ZN(n20726) );
  MUX41 U9667 ( .I0(ram[2648]), .I1(ram[2640]), .I2(ram[2632]), .I3(
        ram[2624]), .S0(n27030), .S1(n26555), .ZN(n20721) );
  MUX41 U9668 ( .I0(ram[1368]), .I1(ram[1360]), .I2(ram[1352]), .I3(
        ram[1344]), .S0(n27027), .S1(n26552), .ZN(n20666) );
  MUX41 U9669 ( .I0(ram[1496]), .I1(ram[1488]), .I2(ram[1480]), .I3(
        ram[1472]), .S0(n27027), .S1(n26552), .ZN(n20671) );
  MUX41 U9670 ( .I0(ram[1240]), .I1(ram[1232]), .I2(ram[1224]), .I3(
        ram[1216]), .S0(n27026), .S1(n26551), .ZN(n20661) );
  MUX41 U9671 ( .I0(ram[1112]), .I1(ram[1104]), .I2(ram[1096]), .I3(
        ram[1088]), .S0(n27026), .S1(n26551), .ZN(n20656) );
  MUX41 U9672 ( .I0(ram[1880]), .I1(ram[1872]), .I2(ram[1864]), .I3(
        ram[1856]), .S0(n27028), .S1(n26553), .ZN(n20686) );
  MUX41 U9673 ( .I0(ram[2008]), .I1(ram[2000]), .I2(ram[1992]), .I3(
        ram[1984]), .S0(n27028), .S1(n26553), .ZN(n20691) );
  MUX41 U9674 ( .I0(ram[1752]), .I1(ram[1744]), .I2(ram[1736]), .I3(
        ram[1728]), .S0(n27028), .S1(n26553), .ZN(n20681) );
  MUX41 U9675 ( .I0(ram[1624]), .I1(ram[1616]), .I2(ram[1608]), .I3(
        ram[1600]), .S0(n27027), .S1(n26552), .ZN(n20676) );
  MUX41 U9676 ( .I0(ram[344]), .I1(ram[336]), .I2(ram[328]), .I3(ram[320]), .S0(n27024), .S1(n26549), .ZN(n20626) );
  MUX41 U9677 ( .I0(ram[472]), .I1(ram[464]), .I2(ram[456]), .I3(ram[448]), .S0(n27025), .S1(n26550), .ZN(n20631) );
  MUX41 U9678 ( .I0(ram[216]), .I1(ram[208]), .I2(ram[200]), .I3(ram[192]), .S0(n27024), .S1(n26549), .ZN(n3711) );
  MUX41 U9679 ( .I0(ram[88]), .I1(ram[80]), .I2(ram[72]), .I3(ram[64]), 
        .S0(n27024), .S1(n26549), .ZN(n3065) );
  MUX41 U9680 ( .I0(ram[856]), .I1(ram[848]), .I2(ram[840]), .I3(ram[832]), .S0(n27025), .S1(n26550), .ZN(n20646) );
  MUX41 U9681 ( .I0(ram[984]), .I1(ram[976]), .I2(ram[968]), .I3(ram[960]), .S0(n27026), .S1(n26551), .ZN(n20651) );
  MUX41 U9682 ( .I0(ram[3417]), .I1(ram[3409]), .I2(ram[3401]), .I3(
        ram[3393]), .S0(n27071), .S1(n26596), .ZN(n21435) );
  MUX41 U9683 ( .I0(ram[3545]), .I1(ram[3537]), .I2(ram[3529]), .I3(
        ram[3521]), .S0(n27071), .S1(n26596), .ZN(n21440) );
  MUX41 U9684 ( .I0(ram[3289]), .I1(ram[3281]), .I2(ram[3273]), .I3(
        ram[3265]), .S0(n27071), .S1(n26596), .ZN(n21430) );
  MUX41 U9685 ( .I0(ram[3161]), .I1(ram[3153]), .I2(ram[3145]), .I3(
        ram[3137]), .S0(n27070), .S1(n26595), .ZN(n21425) );
  MUX41 U9686 ( .I0(ram[3929]), .I1(ram[3921]), .I2(ram[3913]), .I3(
        ram[3905]), .S0(n27072), .S1(n26597), .ZN(n21455) );
  MUX41 U9687 ( .I0(ram[4057]), .I1(ram[4049]), .I2(ram[4041]), .I3(
        ram[4033]), .S0(n27073), .S1(n26598), .ZN(n21460) );
  MUX41 U9688 ( .I0(ram[3801]), .I1(ram[3793]), .I2(ram[3785]), .I3(
        ram[3777]), .S0(n27072), .S1(n26597), .ZN(n21450) );
  MUX41 U9689 ( .I0(ram[3673]), .I1(ram[3665]), .I2(ram[3657]), .I3(
        ram[3649]), .S0(n27072), .S1(n26597), .ZN(n21445) );
  MUX41 U9690 ( .I0(ram[2393]), .I1(ram[2385]), .I2(ram[2377]), .I3(
        ram[2369]), .S0(n27069), .S1(n26594), .ZN(n21395) );
  MUX41 U9691 ( .I0(ram[2521]), .I1(ram[2513]), .I2(ram[2505]), .I3(
        ram[2497]), .S0(n27069), .S1(n26594), .ZN(n21400) );
  MUX41 U9692 ( .I0(ram[2265]), .I1(ram[2257]), .I2(ram[2249]), .I3(
        ram[2241]), .S0(n27068), .S1(n26593), .ZN(n21390) );
  MUX41 U9693 ( .I0(ram[2137]), .I1(ram[2129]), .I2(ram[2121]), .I3(
        ram[2113]), .S0(n27068), .S1(n26593), .ZN(n21385) );
  MUX41 U9694 ( .I0(ram[2905]), .I1(ram[2897]), .I2(ram[2889]), .I3(
        ram[2881]), .S0(n27070), .S1(n26595), .ZN(n21415) );
  MUX41 U9695 ( .I0(ram[3033]), .I1(ram[3025]), .I2(ram[3017]), .I3(
        ram[3009]), .S0(n27070), .S1(n26595), .ZN(n21420) );
  MUX41 U9696 ( .I0(ram[2777]), .I1(ram[2769]), .I2(ram[2761]), .I3(
        ram[2753]), .S0(n27069), .S1(n26594), .ZN(n21410) );
  MUX41 U9697 ( .I0(ram[2649]), .I1(ram[2641]), .I2(ram[2633]), .I3(
        ram[2625]), .S0(n27069), .S1(n26594), .ZN(n21405) );
  MUX41 U9698 ( .I0(ram[1369]), .I1(ram[1361]), .I2(ram[1353]), .I3(
        ram[1345]), .S0(n27066), .S1(n26591), .ZN(n21350) );
  MUX41 U9699 ( .I0(ram[1497]), .I1(ram[1489]), .I2(ram[1481]), .I3(
        ram[1473]), .S0(n27066), .S1(n26591), .ZN(n21355) );
  MUX41 U9700 ( .I0(ram[1241]), .I1(ram[1233]), .I2(ram[1225]), .I3(
        ram[1217]), .S0(n27066), .S1(n26591), .ZN(n21345) );
  MUX41 U9701 ( .I0(ram[1113]), .I1(ram[1105]), .I2(ram[1097]), .I3(
        ram[1089]), .S0(n27065), .S1(n26590), .ZN(n21340) );
  MUX41 U9702 ( .I0(ram[1881]), .I1(ram[1873]), .I2(ram[1865]), .I3(
        ram[1857]), .S0(n27067), .S1(n26592), .ZN(n21370) );
  MUX41 U9703 ( .I0(ram[2009]), .I1(ram[2001]), .I2(ram[1993]), .I3(
        ram[1985]), .S0(n27068), .S1(n26593), .ZN(n21375) );
  MUX41 U9704 ( .I0(ram[1753]), .I1(ram[1745]), .I2(ram[1737]), .I3(
        ram[1729]), .S0(n27067), .S1(n26592), .ZN(n21365) );
  MUX41 U9705 ( .I0(ram[1625]), .I1(ram[1617]), .I2(ram[1609]), .I3(
        ram[1601]), .S0(n27067), .S1(n26592), .ZN(n21360) );
  MUX41 U9706 ( .I0(ram[345]), .I1(ram[337]), .I2(ram[329]), .I3(ram[321]), .S0(n27064), .S1(n26589), .ZN(n21310) );
  MUX41 U9707 ( .I0(ram[473]), .I1(ram[465]), .I2(ram[457]), .I3(ram[449]), .S0(n27064), .S1(n26589), .ZN(n21315) );
  MUX41 U9708 ( .I0(ram[217]), .I1(ram[209]), .I2(ram[201]), .I3(ram[193]), .S0(n27063), .S1(n26588), .ZN(n21305) );
  MUX41 U9709 ( .I0(ram[89]), .I1(ram[81]), .I2(ram[73]), .I3(ram[65]), 
        .S0(n27063), .S1(n26588), .ZN(n21300) );
  MUX41 U9710 ( .I0(ram[857]), .I1(ram[849]), .I2(ram[841]), .I3(ram[833]), .S0(n27065), .S1(n26590), .ZN(n21330) );
  MUX41 U9711 ( .I0(ram[985]), .I1(ram[977]), .I2(ram[969]), .I3(ram[961]), .S0(n27065), .S1(n26590), .ZN(n21335) );
  MUX41 U9712 ( .I0(ram[729]), .I1(ram[721]), .I2(ram[713]), .I3(ram[705]), .S0(n27065), .S1(n26590), .ZN(n21325) );
  MUX41 U9713 ( .I0(ram[3418]), .I1(ram[3410]), .I2(ram[3402]), .I3(
        ram[3394]), .S0(n27110), .S1(n26635), .ZN(n22119) );
  MUX41 U9714 ( .I0(ram[3546]), .I1(ram[3538]), .I2(ram[3530]), .I3(
        ram[3522]), .S0(n27111), .S1(n26636), .ZN(n22124) );
  MUX41 U9715 ( .I0(ram[3290]), .I1(ram[3282]), .I2(ram[3274]), .I3(
        ram[3266]), .S0(n27110), .S1(n26635), .ZN(n22114) );
  MUX41 U9716 ( .I0(ram[3162]), .I1(ram[3154]), .I2(ram[3146]), .I3(
        ram[3138]), .S0(n27110), .S1(n26635), .ZN(n22109) );
  MUX41 U9717 ( .I0(ram[3930]), .I1(ram[3922]), .I2(ram[3914]), .I3(
        ram[3906]), .S0(n27112), .S1(n26637), .ZN(n22139) );
  MUX41 U9718 ( .I0(ram[4058]), .I1(ram[4050]), .I2(ram[4042]), .I3(
        ram[4034]), .S0(n27112), .S1(n26637), .ZN(n22144) );
  MUX41 U9719 ( .I0(ram[3802]), .I1(ram[3794]), .I2(ram[3786]), .I3(
        ram[3778]), .S0(n27111), .S1(n26636), .ZN(n22134) );
  MUX41 U9720 ( .I0(ram[3674]), .I1(ram[3666]), .I2(ram[3658]), .I3(
        ram[3650]), .S0(n27111), .S1(n26636), .ZN(n22129) );
  MUX41 U9721 ( .I0(ram[2394]), .I1(ram[2386]), .I2(ram[2378]), .I3(
        ram[2370]), .S0(n27108), .S1(n26633), .ZN(n22079) );
  MUX41 U9722 ( .I0(ram[2522]), .I1(ram[2514]), .I2(ram[2506]), .I3(
        ram[2498]), .S0(n27108), .S1(n26633), .ZN(n22084) );
  MUX41 U9723 ( .I0(ram[2266]), .I1(ram[2258]), .I2(ram[2250]), .I3(
        ram[2242]), .S0(n27108), .S1(n26633), .ZN(n22074) );
  MUX41 U9724 ( .I0(ram[2138]), .I1(ram[2130]), .I2(ram[2122]), .I3(
        ram[2114]), .S0(n27107), .S1(n26632), .ZN(n22069) );
  MUX41 U9725 ( .I0(ram[2906]), .I1(ram[2898]), .I2(ram[2890]), .I3(
        ram[2882]), .S0(n27109), .S1(n26634), .ZN(n22099) );
  MUX41 U9726 ( .I0(ram[3034]), .I1(ram[3026]), .I2(ram[3018]), .I3(
        ram[3010]), .S0(n27109), .S1(n26634), .ZN(n22104) );
  MUX41 U9727 ( .I0(ram[2778]), .I1(ram[2770]), .I2(ram[2762]), .I3(
        ram[2754]), .S0(n27109), .S1(n26634), .ZN(n22094) );
  MUX41 U9728 ( .I0(ram[2650]), .I1(ram[2642]), .I2(ram[2634]), .I3(
        ram[2626]), .S0(n27109), .S1(n26634), .ZN(n22089) );
  MUX41 U9729 ( .I0(ram[1370]), .I1(ram[1362]), .I2(ram[1354]), .I3(
        ram[1346]), .S0(n27105), .S1(n26630), .ZN(n22034) );
  MUX41 U9730 ( .I0(ram[1498]), .I1(ram[1490]), .I2(ram[1482]), .I3(
        ram[1474]), .S0(n27106), .S1(n26631), .ZN(n22039) );
  MUX41 U9731 ( .I0(ram[1242]), .I1(ram[1234]), .I2(ram[1226]), .I3(
        ram[1218]), .S0(n27105), .S1(n26630), .ZN(n22029) );
  MUX41 U9732 ( .I0(ram[1114]), .I1(ram[1106]), .I2(ram[1098]), .I3(
        ram[1090]), .S0(n27105), .S1(n26630), .ZN(n22024) );
  MUX41 U9733 ( .I0(ram[1882]), .I1(ram[1874]), .I2(ram[1866]), .I3(
        ram[1858]), .S0(n27107), .S1(n26632), .ZN(n22054) );
  MUX41 U9734 ( .I0(ram[2010]), .I1(ram[2002]), .I2(ram[1994]), .I3(
        ram[1986]), .S0(n27107), .S1(n26632), .ZN(n22059) );
  MUX41 U9735 ( .I0(ram[1754]), .I1(ram[1746]), .I2(ram[1738]), .I3(
        ram[1730]), .S0(n27106), .S1(n26631), .ZN(n22049) );
  MUX41 U9736 ( .I0(ram[1626]), .I1(ram[1618]), .I2(ram[1610]), .I3(
        ram[1602]), .S0(n27106), .S1(n26631), .ZN(n22044) );
  MUX41 U9737 ( .I0(ram[346]), .I1(ram[338]), .I2(ram[330]), .I3(ram[322]), .S0(n27103), .S1(n26628), .ZN(n21994) );
  MUX41 U9738 ( .I0(ram[474]), .I1(ram[466]), .I2(ram[458]), .I3(ram[450]), .S0(n27103), .S1(n26628), .ZN(n21999) );
  MUX41 U9739 ( .I0(ram[218]), .I1(ram[210]), .I2(ram[202]), .I3(ram[194]), .S0(n27103), .S1(n26628), .ZN(n21989) );
  MUX41 U9740 ( .I0(ram[90]), .I1(ram[82]), .I2(ram[74]), .I3(ram[66]), 
        .S0(n27102), .S1(n26627), .ZN(n21984) );
  MUX41 U9741 ( .I0(ram[858]), .I1(ram[850]), .I2(ram[842]), .I3(ram[834]), .S0(n27104), .S1(n26629), .ZN(n22014) );
  MUX41 U9742 ( .I0(ram[986]), .I1(ram[978]), .I2(ram[970]), .I3(ram[962]), .S0(n27105), .S1(n26630), .ZN(n22019) );
  MUX41 U9743 ( .I0(ram[730]), .I1(ram[722]), .I2(ram[714]), .I3(ram[706]), .S0(n27104), .S1(n26629), .ZN(n22009) );
  MUX41 U9744 ( .I0(ram[602]), .I1(ram[594]), .I2(ram[586]), .I3(ram[578]), .S0(n27104), .S1(n26629), .ZN(n22004) );
  MUX41 U9745 ( .I0(ram[3419]), .I1(ram[3411]), .I2(ram[3403]), .I3(
        ram[3395]), .S0(n27150), .S1(n26675), .ZN(n22803) );
  MUX41 U9746 ( .I0(ram[3547]), .I1(ram[3539]), .I2(ram[3531]), .I3(
        ram[3523]), .S0(n27150), .S1(n26675), .ZN(n22808) );
  MUX41 U9747 ( .I0(ram[3291]), .I1(ram[3283]), .I2(ram[3275]), .I3(
        ram[3267]), .S0(n27149), .S1(n26674), .ZN(n22798) );
  MUX41 U9748 ( .I0(ram[3163]), .I1(ram[3155]), .I2(ram[3147]), .I3(
        ram[3139]), .S0(n27149), .S1(n26674), .ZN(n22793) );
  MUX41 U9749 ( .I0(ram[3931]), .I1(ram[3923]), .I2(ram[3915]), .I3(
        ram[3907]), .S0(n27151), .S1(n26676), .ZN(n22823) );
  MUX41 U9750 ( .I0(ram[4059]), .I1(ram[4051]), .I2(ram[4043]), .I3(
        ram[4035]), .S0(n27151), .S1(n26676), .ZN(n22828) );
  MUX41 U9751 ( .I0(ram[3803]), .I1(ram[3795]), .I2(ram[3787]), .I3(
        ram[3779]), .S0(n27151), .S1(n26676), .ZN(n22818) );
  MUX41 U9752 ( .I0(ram[3675]), .I1(ram[3667]), .I2(ram[3659]), .I3(
        ram[3651]), .S0(n27150), .S1(n26675), .ZN(n22813) );
  MUX41 U9753 ( .I0(ram[2395]), .I1(ram[2387]), .I2(ram[2379]), .I3(
        ram[2371]), .S0(n27147), .S1(n26672), .ZN(n22763) );
  MUX41 U9754 ( .I0(ram[2523]), .I1(ram[2515]), .I2(ram[2507]), .I3(
        ram[2499]), .S0(n27148), .S1(n26673), .ZN(n22768) );
  MUX41 U9755 ( .I0(ram[2267]), .I1(ram[2259]), .I2(ram[2251]), .I3(
        ram[2243]), .S0(n27147), .S1(n26672), .ZN(n22758) );
  MUX41 U9756 ( .I0(ram[2139]), .I1(ram[2131]), .I2(ram[2123]), .I3(
        ram[2115]), .S0(n27147), .S1(n26672), .ZN(n22753) );
  MUX41 U9757 ( .I0(ram[2907]), .I1(ram[2899]), .I2(ram[2891]), .I3(
        ram[2883]), .S0(n27149), .S1(n26674), .ZN(n22783) );
  MUX41 U9758 ( .I0(ram[3035]), .I1(ram[3027]), .I2(ram[3019]), .I3(
        ram[3011]), .S0(n27149), .S1(n26674), .ZN(n22788) );
  MUX41 U9759 ( .I0(ram[2779]), .I1(ram[2771]), .I2(ram[2763]), .I3(
        ram[2755]), .S0(n27148), .S1(n26673), .ZN(n22778) );
  MUX41 U9760 ( .I0(ram[2651]), .I1(ram[2643]), .I2(ram[2635]), .I3(
        ram[2627]), .S0(n27148), .S1(n26673), .ZN(n22773) );
  MUX41 U9761 ( .I0(ram[1371]), .I1(ram[1363]), .I2(ram[1355]), .I3(
        ram[1347]), .S0(n27145), .S1(n26670), .ZN(n22718) );
  MUX41 U9762 ( .I0(ram[1499]), .I1(ram[1491]), .I2(ram[1483]), .I3(
        ram[1475]), .S0(n27145), .S1(n26670), .ZN(n22723) );
  MUX41 U9763 ( .I0(ram[1243]), .I1(ram[1235]), .I2(ram[1227]), .I3(
        ram[1219]), .S0(n27145), .S1(n26670), .ZN(n22713) );
  MUX41 U9764 ( .I0(ram[1115]), .I1(ram[1107]), .I2(ram[1099]), .I3(
        ram[1091]), .S0(n27144), .S1(n26669), .ZN(n22708) );
  MUX41 U9765 ( .I0(ram[1883]), .I1(ram[1875]), .I2(ram[1867]), .I3(
        ram[1859]), .S0(n27146), .S1(n26671), .ZN(n22738) );
  MUX41 U9766 ( .I0(ram[2011]), .I1(ram[2003]), .I2(ram[1995]), .I3(
        ram[1987]), .S0(n27146), .S1(n26671), .ZN(n22743) );
  MUX41 U9767 ( .I0(ram[1755]), .I1(ram[1747]), .I2(ram[1739]), .I3(
        ram[1731]), .S0(n27146), .S1(n26671), .ZN(n22733) );
  MUX41 U9768 ( .I0(ram[1627]), .I1(ram[1619]), .I2(ram[1611]), .I3(
        ram[1603]), .S0(n27145), .S1(n26670), .ZN(n22728) );
  MUX41 U9769 ( .I0(ram[347]), .I1(ram[339]), .I2(ram[331]), .I3(ram[323]), .S0(n27142), .S1(n26667), .ZN(n22678) );
  MUX41 U9770 ( .I0(ram[475]), .I1(ram[467]), .I2(ram[459]), .I3(ram[451]), .S0(n27143), .S1(n26668), .ZN(n22683) );
  MUX41 U9771 ( .I0(ram[219]), .I1(ram[211]), .I2(ram[203]), .I3(ram[195]), .S0(n27142), .S1(n26667), .ZN(n22673) );
  MUX41 U9772 ( .I0(ram[91]), .I1(ram[83]), .I2(ram[75]), .I3(ram[67]), 
        .S0(n27142), .S1(n26667), .ZN(n22668) );
  MUX41 U9773 ( .I0(ram[859]), .I1(ram[851]), .I2(ram[843]), .I3(ram[835]), .S0(n27144), .S1(n26669), .ZN(n22698) );
  MUX41 U9774 ( .I0(ram[987]), .I1(ram[979]), .I2(ram[971]), .I3(ram[963]), .S0(n27144), .S1(n26669), .ZN(n22703) );
  MUX41 U9775 ( .I0(ram[731]), .I1(ram[723]), .I2(ram[715]), .I3(ram[707]), .S0(n27143), .S1(n26668), .ZN(n22693) );
  MUX41 U9776 ( .I0(ram[603]), .I1(ram[595]), .I2(ram[587]), .I3(ram[579]), .S0(n27143), .S1(n26668), .ZN(n22688) );
  MUX41 U9777 ( .I0(ram[3420]), .I1(ram[3412]), .I2(ram[3404]), .I3(
        ram[3396]), .S0(n27189), .S1(n26714), .ZN(n23487) );
  MUX41 U9778 ( .I0(ram[3548]), .I1(ram[3540]), .I2(ram[3532]), .I3(
        ram[3524]), .S0(n27189), .S1(n26714), .ZN(n23492) );
  MUX41 U9779 ( .I0(ram[3292]), .I1(ram[3284]), .I2(ram[3276]), .I3(
        ram[3268]), .S0(n27189), .S1(n26714), .ZN(n23482) );
  MUX41 U9780 ( .I0(ram[3164]), .I1(ram[3156]), .I2(ram[3148]), .I3(
        ram[3140]), .S0(n27189), .S1(n26714), .ZN(n23477) );
  MUX41 U9781 ( .I0(ram[3932]), .I1(ram[3924]), .I2(ram[3916]), .I3(
        ram[3908]), .S0(n27190), .S1(n26715), .ZN(n23507) );
  MUX41 U9782 ( .I0(ram[4060]), .I1(ram[4052]), .I2(ram[4044]), .I3(
        ram[4036]), .S0(n27191), .S1(n26716), .ZN(n23512) );
  MUX41 U9783 ( .I0(ram[3804]), .I1(ram[3796]), .I2(ram[3788]), .I3(
        ram[3780]), .S0(n27190), .S1(n26715), .ZN(n23502) );
  MUX41 U9784 ( .I0(ram[3676]), .I1(ram[3668]), .I2(ram[3660]), .I3(
        ram[3652]), .S0(n27190), .S1(n26715), .ZN(n23497) );
  MUX41 U9785 ( .I0(ram[2396]), .I1(ram[2388]), .I2(ram[2380]), .I3(
        ram[2372]), .S0(n27187), .S1(n26712), .ZN(n23447) );
  MUX41 U9786 ( .I0(ram[2524]), .I1(ram[2516]), .I2(ram[2508]), .I3(
        ram[2500]), .S0(n27187), .S1(n26712), .ZN(n23452) );
  MUX41 U9787 ( .I0(ram[2268]), .I1(ram[2260]), .I2(ram[2252]), .I3(
        ram[2244]), .S0(n27186), .S1(n26711), .ZN(n23442) );
  MUX41 U9788 ( .I0(ram[2140]), .I1(ram[2132]), .I2(ram[2124]), .I3(
        ram[2116]), .S0(n27186), .S1(n26711), .ZN(n23437) );
  MUX41 U9789 ( .I0(ram[2908]), .I1(ram[2900]), .I2(ram[2892]), .I3(
        ram[2884]), .S0(n27188), .S1(n26713), .ZN(n23467) );
  MUX41 U9790 ( .I0(ram[3036]), .I1(ram[3028]), .I2(ram[3020]), .I3(
        ram[3012]), .S0(n27188), .S1(n26713), .ZN(n23472) );
  MUX41 U9791 ( .I0(ram[2780]), .I1(ram[2772]), .I2(ram[2764]), .I3(
        ram[2756]), .S0(n27188), .S1(n26713), .ZN(n23462) );
  MUX41 U9792 ( .I0(ram[2652]), .I1(ram[2644]), .I2(ram[2636]), .I3(
        ram[2628]), .S0(n27187), .S1(n26712), .ZN(n23457) );
  MUX41 U9793 ( .I0(ram[1372]), .I1(ram[1364]), .I2(ram[1356]), .I3(
        ram[1348]), .S0(n27184), .S1(n26709), .ZN(n23402) );
  MUX41 U9794 ( .I0(ram[1500]), .I1(ram[1492]), .I2(ram[1484]), .I3(
        ram[1476]), .S0(n27185), .S1(n26710), .ZN(n23407) );
  MUX41 U9795 ( .I0(ram[1244]), .I1(ram[1236]), .I2(ram[1228]), .I3(
        ram[1220]), .S0(n27184), .S1(n26709), .ZN(n23397) );
  MUX41 U9796 ( .I0(ram[1116]), .I1(ram[1108]), .I2(ram[1100]), .I3(
        ram[1092]), .S0(n27184), .S1(n26709), .ZN(n23392) );
  MUX41 U9797 ( .I0(ram[1884]), .I1(ram[1876]), .I2(ram[1868]), .I3(
        ram[1860]), .S0(n27185), .S1(n26710), .ZN(n23422) );
  MUX41 U9798 ( .I0(ram[2012]), .I1(ram[2004]), .I2(ram[1996]), .I3(
        ram[1988]), .S0(n27186), .S1(n26711), .ZN(n23427) );
  MUX41 U9799 ( .I0(ram[1756]), .I1(ram[1748]), .I2(ram[1740]), .I3(
        ram[1732]), .S0(n27185), .S1(n26710), .ZN(n23417) );
  MUX41 U9800 ( .I0(ram[1628]), .I1(ram[1620]), .I2(ram[1612]), .I3(
        ram[1604]), .S0(n27185), .S1(n26710), .ZN(n23412) );
  MUX41 U9801 ( .I0(ram[348]), .I1(ram[340]), .I2(ram[332]), .I3(ram[324]), .S0(n27182), .S1(n26707), .ZN(n23362) );
  MUX41 U9802 ( .I0(ram[476]), .I1(ram[468]), .I2(ram[460]), .I3(ram[452]), .S0(n27182), .S1(n26707), .ZN(n23367) );
  MUX41 U9803 ( .I0(ram[220]), .I1(ram[212]), .I2(ram[204]), .I3(ram[196]), .S0(n27181), .S1(n26706), .ZN(n23357) );
  MUX41 U9804 ( .I0(ram[92]), .I1(ram[84]), .I2(ram[76]), .I3(ram[68]), 
        .S0(n27181), .S1(n26706), .ZN(n23352) );
  MUX41 U9805 ( .I0(ram[860]), .I1(ram[852]), .I2(ram[844]), .I3(ram[836]), .S0(n27183), .S1(n26708), .ZN(n23382) );
  MUX41 U9806 ( .I0(ram[988]), .I1(ram[980]), .I2(ram[972]), .I3(ram[964]), .S0(n27183), .S1(n26708), .ZN(n23387) );
  MUX41 U9807 ( .I0(ram[732]), .I1(ram[724]), .I2(ram[716]), .I3(ram[708]), .S0(n27183), .S1(n26708), .ZN(n23377) );
  MUX41 U9808 ( .I0(ram[604]), .I1(ram[596]), .I2(ram[588]), .I3(ram[580]), .S0(n27182), .S1(n26707), .ZN(n23372) );
  MUX41 U9809 ( .I0(ram[3421]), .I1(ram[3413]), .I2(ram[3405]), .I3(
        ram[3397]), .S0(n27229), .S1(n26754), .ZN(n24171) );
  MUX41 U9810 ( .I0(ram[3549]), .I1(ram[3541]), .I2(ram[3533]), .I3(
        ram[3525]), .S0(n27229), .S1(n26754), .ZN(n24176) );
  MUX41 U9811 ( .I0(ram[3293]), .I1(ram[3285]), .I2(ram[3277]), .I3(
        ram[3269]), .S0(n27228), .S1(n26753), .ZN(n24166) );
  MUX41 U9812 ( .I0(ram[3165]), .I1(ram[3157]), .I2(ram[3149]), .I3(
        ram[3141]), .S0(n27228), .S1(n26753), .ZN(n24161) );
  MUX41 U9813 ( .I0(ram[3933]), .I1(ram[3925]), .I2(ram[3917]), .I3(
        ram[3909]), .S0(n27230), .S1(n26755), .ZN(n24191) );
  MUX41 U9814 ( .I0(ram[4061]), .I1(ram[4053]), .I2(ram[4045]), .I3(
        ram[4037]), .S0(n27230), .S1(n26755), .ZN(n24196) );
  MUX41 U9815 ( .I0(ram[3805]), .I1(ram[3797]), .I2(ram[3789]), .I3(
        ram[3781]), .S0(n27229), .S1(n26754), .ZN(n24186) );
  MUX41 U9816 ( .I0(ram[3677]), .I1(ram[3669]), .I2(ram[3661]), .I3(
        ram[3653]), .S0(n27229), .S1(n26754), .ZN(n24181) );
  MUX41 U9817 ( .I0(ram[2397]), .I1(ram[2389]), .I2(ram[2381]), .I3(
        ram[2373]), .S0(n27226), .S1(n26751), .ZN(n24131) );
  MUX41 U9818 ( .I0(ram[2525]), .I1(ram[2517]), .I2(ram[2509]), .I3(
        ram[2501]), .S0(n27226), .S1(n26751), .ZN(n24136) );
  MUX41 U9819 ( .I0(ram[2269]), .I1(ram[2261]), .I2(ram[2253]), .I3(
        ram[2245]), .S0(n27226), .S1(n26751), .ZN(n24126) );
  MUX41 U9820 ( .I0(ram[2141]), .I1(ram[2133]), .I2(ram[2125]), .I3(
        ram[2117]), .S0(n27225), .S1(n26750), .ZN(n24121) );
  MUX41 U9821 ( .I0(ram[2909]), .I1(ram[2901]), .I2(ram[2893]), .I3(
        ram[2885]), .S0(n27227), .S1(n26752), .ZN(n24151) );
  MUX41 U9822 ( .I0(ram[3037]), .I1(ram[3029]), .I2(ram[3021]), .I3(
        ram[3013]), .S0(n27228), .S1(n26753), .ZN(n24156) );
  MUX41 U9823 ( .I0(ram[2781]), .I1(ram[2773]), .I2(ram[2765]), .I3(
        ram[2757]), .S0(n27227), .S1(n26752), .ZN(n24146) );
  MUX41 U9824 ( .I0(ram[2653]), .I1(ram[2645]), .I2(ram[2637]), .I3(
        ram[2629]), .S0(n27227), .S1(n26752), .ZN(n24141) );
  MUX41 U9825 ( .I0(ram[1373]), .I1(ram[1365]), .I2(ram[1357]), .I3(
        ram[1349]), .S0(n27224), .S1(n26749), .ZN(n24086) );
  MUX41 U9826 ( .I0(ram[1501]), .I1(ram[1493]), .I2(ram[1485]), .I3(
        ram[1477]), .S0(n27224), .S1(n26749), .ZN(n24091) );
  MUX41 U9827 ( .I0(ram[1245]), .I1(ram[1237]), .I2(ram[1229]), .I3(
        ram[1221]), .S0(n27223), .S1(n26748), .ZN(n24081) );
  MUX41 U9828 ( .I0(ram[1117]), .I1(ram[1109]), .I2(ram[1101]), .I3(
        ram[1093]), .S0(n27223), .S1(n26748), .ZN(n24076) );
  MUX41 U9829 ( .I0(ram[1885]), .I1(ram[1877]), .I2(ram[1869]), .I3(
        ram[1861]), .S0(n27225), .S1(n26750), .ZN(n24106) );
  MUX41 U9830 ( .I0(ram[2013]), .I1(ram[2005]), .I2(ram[1997]), .I3(
        ram[1989]), .S0(n27225), .S1(n26750), .ZN(n24111) );
  MUX41 U9831 ( .I0(ram[1757]), .I1(ram[1749]), .I2(ram[1741]), .I3(
        ram[1733]), .S0(n27225), .S1(n26750), .ZN(n24101) );
  MUX41 U9832 ( .I0(ram[1629]), .I1(ram[1621]), .I2(ram[1613]), .I3(
        ram[1605]), .S0(n27224), .S1(n26749), .ZN(n24096) );
  MUX41 U9833 ( .I0(ram[349]), .I1(ram[341]), .I2(ram[333]), .I3(ram[325]), .S0(n27221), .S1(n26746), .ZN(n24046) );
  MUX41 U9834 ( .I0(ram[477]), .I1(ram[469]), .I2(ram[461]), .I3(ram[453]), .S0(n27221), .S1(n26746), .ZN(n24051) );
  MUX41 U9835 ( .I0(ram[221]), .I1(ram[213]), .I2(ram[205]), .I3(ram[197]), .S0(n27221), .S1(n26746), .ZN(n24041) );
  MUX41 U9836 ( .I0(ram[93]), .I1(ram[85]), .I2(ram[77]), .I3(ram[69]), 
        .S0(n27221), .S1(n26746), .ZN(n24036) );
  MUX41 U9837 ( .I0(ram[861]), .I1(ram[853]), .I2(ram[845]), .I3(ram[837]), .S0(n27222), .S1(n26747), .ZN(n24066) );
  MUX41 U9838 ( .I0(ram[989]), .I1(ram[981]), .I2(ram[973]), .I3(ram[965]), .S0(n27223), .S1(n26748), .ZN(n24071) );
  MUX41 U9839 ( .I0(ram[733]), .I1(ram[725]), .I2(ram[717]), .I3(ram[709]), .S0(n27222), .S1(n26747), .ZN(n24061) );
  MUX41 U9840 ( .I0(ram[605]), .I1(ram[597]), .I2(ram[589]), .I3(ram[581]), .S0(n27222), .S1(n26747), .ZN(n24056) );
  MUX41 U9841 ( .I0(ram[3422]), .I1(ram[3414]), .I2(ram[3406]), .I3(
        ram[3398]), .S0(n27268), .S1(n26793), .ZN(n24855) );
  MUX41 U9842 ( .I0(ram[3550]), .I1(ram[3542]), .I2(ram[3534]), .I3(
        ram[3526]), .S0(n27268), .S1(n26793), .ZN(n24860) );
  MUX41 U9843 ( .I0(ram[3294]), .I1(ram[3286]), .I2(ram[3278]), .I3(
        ram[3270]), .S0(n27268), .S1(n26793), .ZN(n24850) );
  MUX41 U9844 ( .I0(ram[3166]), .I1(ram[3158]), .I2(ram[3150]), .I3(
        ram[3142]), .S0(n27267), .S1(n26792), .ZN(n24845) );
  MUX41 U9845 ( .I0(ram[3934]), .I1(ram[3926]), .I2(ram[3918]), .I3(
        ram[3910]), .S0(n27269), .S1(n26794), .ZN(n24875) );
  MUX41 U9846 ( .I0(ram[4062]), .I1(ram[4054]), .I2(ram[4046]), .I3(
        ram[4038]), .S0(n27269), .S1(n26794), .ZN(n24880) );
  MUX41 U9847 ( .I0(ram[3806]), .I1(ram[3798]), .I2(ram[3790]), .I3(
        ram[3782]), .S0(n27269), .S1(n26794), .ZN(n24870) );
  MUX41 U9848 ( .I0(ram[3678]), .I1(ram[3670]), .I2(ram[3662]), .I3(
        ram[3654]), .S0(n27269), .S1(n26794), .ZN(n24865) );
  MUX41 U9849 ( .I0(ram[2398]), .I1(ram[2390]), .I2(ram[2382]), .I3(
        ram[2374]), .S0(n27265), .S1(n26790), .ZN(n24815) );
  MUX41 U9850 ( .I0(ram[2526]), .I1(ram[2518]), .I2(ram[2510]), .I3(
        ram[2502]), .S0(n27266), .S1(n26791), .ZN(n24820) );
  MUX41 U9851 ( .I0(ram[2270]), .I1(ram[2262]), .I2(ram[2254]), .I3(
        ram[2246]), .S0(n27265), .S1(n26790), .ZN(n24810) );
  MUX41 U9852 ( .I0(ram[2142]), .I1(ram[2134]), .I2(ram[2126]), .I3(
        ram[2118]), .S0(n27265), .S1(n26790), .ZN(n24805) );
  MUX41 U9853 ( .I0(ram[2910]), .I1(ram[2902]), .I2(ram[2894]), .I3(
        ram[2886]), .S0(n27267), .S1(n26792), .ZN(n24835) );
  MUX41 U9854 ( .I0(ram[3038]), .I1(ram[3030]), .I2(ram[3022]), .I3(
        ram[3014]), .S0(n27267), .S1(n26792), .ZN(n24840) );
  MUX41 U9855 ( .I0(ram[2782]), .I1(ram[2774]), .I2(ram[2766]), .I3(
        ram[2758]), .S0(n27266), .S1(n26791), .ZN(n24830) );
  MUX41 U9856 ( .I0(ram[2654]), .I1(ram[2646]), .I2(ram[2638]), .I3(
        ram[2630]), .S0(n27266), .S1(n26791), .ZN(n24825) );
  MUX41 U9857 ( .I0(ram[1374]), .I1(ram[1366]), .I2(ram[1358]), .I3(
        ram[1350]), .S0(n27263), .S1(n26788), .ZN(n24770) );
  MUX41 U9858 ( .I0(ram[1502]), .I1(ram[1494]), .I2(ram[1486]), .I3(
        ram[1478]), .S0(n27263), .S1(n26788), .ZN(n24775) );
  MUX41 U9859 ( .I0(ram[1246]), .I1(ram[1238]), .I2(ram[1230]), .I3(
        ram[1222]), .S0(n27263), .S1(n26788), .ZN(n24765) );
  MUX41 U9860 ( .I0(ram[1118]), .I1(ram[1110]), .I2(ram[1102]), .I3(
        ram[1094]), .S0(n27262), .S1(n26787), .ZN(n24760) );
  MUX41 U9861 ( .I0(ram[1886]), .I1(ram[1878]), .I2(ram[1870]), .I3(
        ram[1862]), .S0(n27264), .S1(n26789), .ZN(n24790) );
  MUX41 U9862 ( .I0(ram[2014]), .I1(ram[2006]), .I2(ram[1998]), .I3(
        ram[1990]), .S0(n27265), .S1(n26790), .ZN(n24795) );
  MUX41 U9863 ( .I0(ram[1758]), .I1(ram[1750]), .I2(ram[1742]), .I3(
        ram[1734]), .S0(n27264), .S1(n26789), .ZN(n24785) );
  MUX41 U9864 ( .I0(ram[1630]), .I1(ram[1622]), .I2(ram[1614]), .I3(
        ram[1606]), .S0(n27264), .S1(n26789), .ZN(n24780) );
  MUX41 U9865 ( .I0(ram[350]), .I1(ram[342]), .I2(ram[334]), .I3(ram[326]), .S0(n27261), .S1(n26786), .ZN(n24730) );
  MUX41 U9866 ( .I0(ram[478]), .I1(ram[470]), .I2(ram[462]), .I3(ram[454]), .S0(n27261), .S1(n26786), .ZN(n24735) );
  MUX41 U9867 ( .I0(ram[222]), .I1(ram[214]), .I2(ram[206]), .I3(ram[198]), .S0(n27260), .S1(n26785), .ZN(n24725) );
  MUX41 U9868 ( .I0(ram[94]), .I1(ram[86]), .I2(ram[78]), .I3(ram[70]), 
        .S0(n27260), .S1(n26785), .ZN(n24720) );
  MUX41 U9869 ( .I0(ram[862]), .I1(ram[854]), .I2(ram[846]), .I3(ram[838]), .S0(n27262), .S1(n26787), .ZN(n24750) );
  MUX41 U9870 ( .I0(ram[990]), .I1(ram[982]), .I2(ram[974]), .I3(ram[966]), .S0(n27262), .S1(n26787), .ZN(n24755) );
  MUX41 U9871 ( .I0(ram[734]), .I1(ram[726]), .I2(ram[718]), .I3(ram[710]), .S0(n27261), .S1(n26786), .ZN(n24745) );
  MUX41 U9872 ( .I0(ram[606]), .I1(ram[598]), .I2(ram[590]), .I3(ram[582]), .S0(n27261), .S1(n26786), .ZN(n24740) );
  MUX41 U9873 ( .I0(ram[3423]), .I1(ram[3415]), .I2(ram[3407]), .I3(
        ram[3399]), .S0(n27307), .S1(n26832), .ZN(n25539) );
  MUX41 U9874 ( .I0(ram[3551]), .I1(ram[3543]), .I2(ram[3535]), .I3(
        ram[3527]), .S0(n27308), .S1(n26833), .ZN(n25544) );
  MUX41 U9875 ( .I0(ram[3295]), .I1(ram[3287]), .I2(ram[3279]), .I3(
        ram[3271]), .S0(n27307), .S1(n26832), .ZN(n25534) );
  MUX41 U9876 ( .I0(ram[3167]), .I1(ram[3159]), .I2(ram[3151]), .I3(
        ram[3143]), .S0(n27307), .S1(n26832), .ZN(n25529) );
  MUX41 U9877 ( .I0(ram[3935]), .I1(ram[3927]), .I2(ram[3919]), .I3(
        ram[3911]), .S0(n27309), .S1(n26834), .ZN(n25559) );
  MUX41 U9878 ( .I0(ram[4063]), .I1(ram[4055]), .I2(ram[4047]), .I3(
        ram[4039]), .S0(n27309), .S1(n26834), .ZN(n25564) );
  MUX41 U9879 ( .I0(ram[3807]), .I1(ram[3799]), .I2(ram[3791]), .I3(
        ram[3783]), .S0(n27308), .S1(n26833), .ZN(n25554) );
  MUX41 U9880 ( .I0(ram[3679]), .I1(ram[3671]), .I2(ram[3663]), .I3(
        ram[3655]), .S0(n27308), .S1(n26833), .ZN(n25549) );
  MUX41 U9881 ( .I0(ram[2399]), .I1(ram[2391]), .I2(ram[2383]), .I3(
        ram[2375]), .S0(n27305), .S1(n26830), .ZN(n25499) );
  MUX41 U9882 ( .I0(ram[2527]), .I1(ram[2519]), .I2(ram[2511]), .I3(
        ram[2503]), .S0(n27305), .S1(n26830), .ZN(n25504) );
  MUX41 U9883 ( .I0(ram[2271]), .I1(ram[2263]), .I2(ram[2255]), .I3(
        ram[2247]), .S0(n27305), .S1(n26830), .ZN(n25494) );
  MUX41 U9884 ( .I0(ram[2143]), .I1(ram[2135]), .I2(ram[2127]), .I3(
        ram[2119]), .S0(n27304), .S1(n26829), .ZN(n25489) );
  MUX41 U9885 ( .I0(ram[2911]), .I1(ram[2903]), .I2(ram[2895]), .I3(
        ram[2887]), .S0(n27306), .S1(n26831), .ZN(n25519) );
  MUX41 U9886 ( .I0(ram[3039]), .I1(ram[3031]), .I2(ram[3023]), .I3(
        ram[3015]), .S0(n27306), .S1(n26831), .ZN(n25524) );
  MUX41 U9887 ( .I0(ram[2783]), .I1(ram[2775]), .I2(ram[2767]), .I3(
        ram[2759]), .S0(n27306), .S1(n26831), .ZN(n25514) );
  MUX41 U9888 ( .I0(ram[2655]), .I1(ram[2647]), .I2(ram[2639]), .I3(
        ram[2631]), .S0(n27305), .S1(n26830), .ZN(n25509) );
  MUX41 U9889 ( .I0(ram[1375]), .I1(ram[1367]), .I2(ram[1359]), .I3(
        ram[1351]), .S0(n27302), .S1(n26827), .ZN(n25454) );
  MUX41 U9890 ( .I0(ram[1503]), .I1(ram[1495]), .I2(ram[1487]), .I3(
        ram[1479]), .S0(n27303), .S1(n26828), .ZN(n25459) );
  MUX41 U9891 ( .I0(ram[1247]), .I1(ram[1239]), .I2(ram[1231]), .I3(
        ram[1223]), .S0(n27302), .S1(n26827), .ZN(n25449) );
  MUX41 U9892 ( .I0(ram[1119]), .I1(ram[1111]), .I2(ram[1103]), .I3(
        ram[1095]), .S0(n27302), .S1(n26827), .ZN(n25444) );
  MUX41 U9893 ( .I0(ram[1887]), .I1(ram[1879]), .I2(ram[1871]), .I3(
        ram[1863]), .S0(n27304), .S1(n26829), .ZN(n25474) );
  MUX41 U9894 ( .I0(ram[2015]), .I1(ram[2007]), .I2(ram[1999]), .I3(
        ram[1991]), .S0(n27304), .S1(n26829), .ZN(n25479) );
  MUX41 U9895 ( .I0(ram[1759]), .I1(ram[1751]), .I2(ram[1743]), .I3(
        ram[1735]), .S0(n27303), .S1(n26828), .ZN(n25469) );
  MUX41 U9896 ( .I0(ram[1631]), .I1(ram[1623]), .I2(ram[1615]), .I3(
        ram[1607]), .S0(n27303), .S1(n26828), .ZN(n25464) );
  MUX41 U9897 ( .I0(ram[351]), .I1(ram[343]), .I2(ram[335]), .I3(ram[327]), .S0(n27300), .S1(n26825), .ZN(n25414) );
  MUX41 U9898 ( .I0(ram[479]), .I1(ram[471]), .I2(ram[463]), .I3(ram[455]), .S0(n27300), .S1(n26825), .ZN(n25419) );
  MUX41 U9899 ( .I0(ram[223]), .I1(ram[215]), .I2(ram[207]), .I3(ram[199]), .S0(n27300), .S1(n26825), .ZN(n25409) );
  MUX41 U9900 ( .I0(ram[95]), .I1(ram[87]), .I2(ram[79]), .I3(ram[71]), 
        .S0(n27299), .S1(n26824), .ZN(n25404) );
  MUX41 U9901 ( .I0(ram[863]), .I1(ram[855]), .I2(ram[847]), .I3(ram[839]), .S0(n27301), .S1(n26826), .ZN(n25434) );
  MUX41 U9902 ( .I0(ram[991]), .I1(ram[983]), .I2(ram[975]), .I3(ram[967]), .S0(n27301), .S1(n26826), .ZN(n25439) );
  MUX41 U9903 ( .I0(ram[735]), .I1(ram[727]), .I2(ram[719]), .I3(ram[711]), .S0(n27301), .S1(n26826), .ZN(n25429) );
  MUX41 U9904 ( .I0(ram[607]), .I1(ram[599]), .I2(ram[591]), .I3(ram[583]), .S0(n27301), .S1(n26826), .ZN(n25424) );
  MUX41 U9905 ( .I0(ram[15704]), .I1(ram[15696]), .I2(ram[15688]), .I3(
        ram[15680]), .S0(n27061), .S1(n26586), .ZN(n21264) );
  MUX41 U9906 ( .I0(ram[15832]), .I1(ram[15824]), .I2(ram[15816]), .I3(
        ram[15808]), .S0(n27061), .S1(n26586), .ZN(n21269) );
  MUX41 U9907 ( .I0(ram[15576]), .I1(ram[15568]), .I2(ram[15560]), .I3(
        ram[15552]), .S0(n27061), .S1(n26586), .ZN(n21259) );
  MUX41 U9908 ( .I0(ram[15448]), .I1(ram[15440]), .I2(ram[15432]), .I3(
        ram[15424]), .S0(n27061), .S1(n26586), .ZN(n21254) );
  MUX41 U9909 ( .I0(ram[16216]), .I1(ram[16208]), .I2(ram[16200]), .I3(
        ram[16192]), .S0(n27062), .S1(n26587), .ZN(n21284) );
  MUX41 U9910 ( .I0(ram[16344]), .I1(ram[16336]), .I2(ram[16328]), .I3(
        ram[16320]), .S0(n27063), .S1(n26588), .ZN(n21289) );
  MUX41 U9911 ( .I0(ram[16088]), .I1(ram[16080]), .I2(ram[16072]), .I3(
        ram[16064]), .S0(n27062), .S1(n26587), .ZN(n21279) );
  MUX41 U9912 ( .I0(ram[15960]), .I1(ram[15952]), .I2(ram[15944]), .I3(
        ram[15936]), .S0(n27062), .S1(n26587), .ZN(n21274) );
  MUX41 U9913 ( .I0(ram[15192]), .I1(ram[15184]), .I2(ram[15176]), .I3(
        ram[15168]), .S0(n27060), .S1(n26585), .ZN(n21244) );
  MUX41 U9914 ( .I0(ram[15320]), .I1(ram[15312]), .I2(ram[15304]), .I3(
        ram[15296]), .S0(n27060), .S1(n26585), .ZN(n21249) );
  MUX41 U9915 ( .I0(ram[15064]), .I1(ram[15056]), .I2(ram[15048]), .I3(
        ram[15040]), .S0(n27060), .S1(n26585), .ZN(n21239) );
  MUX41 U9916 ( .I0(ram[14936]), .I1(ram[14928]), .I2(ram[14920]), .I3(
        ram[14912]), .S0(n27059), .S1(n26584), .ZN(n21234) );
  MUX41 U9917 ( .I0(ram[14680]), .I1(ram[14672]), .I2(ram[14664]), .I3(
        ram[14656]), .S0(n27059), .S1(n26584), .ZN(n21224) );
  MUX41 U9918 ( .I0(ram[14808]), .I1(ram[14800]), .I2(ram[14792]), .I3(
        ram[14784]), .S0(n27059), .S1(n26584), .ZN(n21229) );
  MUX41 U9919 ( .I0(ram[14552]), .I1(ram[14544]), .I2(ram[14536]), .I3(
        ram[14528]), .S0(n27058), .S1(n26583), .ZN(n21219) );
  MUX41 U9920 ( .I0(ram[14424]), .I1(ram[14416]), .I2(ram[14408]), .I3(
        ram[14400]), .S0(n27058), .S1(n26583), .ZN(n21214) );
  MUX41 U9921 ( .I0(ram[13656]), .I1(ram[13648]), .I2(ram[13640]), .I3(
        ram[13632]), .S0(n27056), .S1(n26581), .ZN(n21179) );
  MUX41 U9922 ( .I0(ram[13784]), .I1(ram[13776]), .I2(ram[13768]), .I3(
        ram[13760]), .S0(n27057), .S1(n26582), .ZN(n21184) );
  MUX41 U9923 ( .I0(ram[13528]), .I1(ram[13520]), .I2(ram[13512]), .I3(
        ram[13504]), .S0(n27056), .S1(n26581), .ZN(n21174) );
  MUX41 U9924 ( .I0(ram[13400]), .I1(ram[13392]), .I2(ram[13384]), .I3(
        ram[13376]), .S0(n27056), .S1(n26581), .ZN(n21169) );
  MUX41 U9925 ( .I0(ram[14168]), .I1(ram[14160]), .I2(ram[14152]), .I3(
        ram[14144]), .S0(n27057), .S1(n26582), .ZN(n21199) );
  MUX41 U9926 ( .I0(ram[14296]), .I1(ram[14288]), .I2(ram[14280]), .I3(
        ram[14272]), .S0(n27058), .S1(n26583), .ZN(n21204) );
  MUX41 U9927 ( .I0(ram[14040]), .I1(ram[14032]), .I2(ram[14024]), .I3(
        ram[14016]), .S0(n27057), .S1(n26582), .ZN(n21194) );
  MUX41 U9928 ( .I0(ram[13912]), .I1(ram[13904]), .I2(ram[13896]), .I3(
        ram[13888]), .S0(n27057), .S1(n26582), .ZN(n21189) );
  MUX41 U9929 ( .I0(ram[13144]), .I1(ram[13136]), .I2(ram[13128]), .I3(
        ram[13120]), .S0(n27055), .S1(n26580), .ZN(n21159) );
  MUX41 U9930 ( .I0(ram[13272]), .I1(ram[13264]), .I2(ram[13256]), .I3(
        ram[13248]), .S0(n27055), .S1(n26580), .ZN(n21164) );
  MUX41 U9931 ( .I0(ram[13016]), .I1(ram[13008]), .I2(ram[13000]), .I3(
        ram[12992]), .S0(n27055), .S1(n26580), .ZN(n21154) );
  MUX41 U9932 ( .I0(ram[12888]), .I1(ram[12880]), .I2(ram[12872]), .I3(
        ram[12864]), .S0(n27054), .S1(n26579), .ZN(n21149) );
  MUX41 U9933 ( .I0(ram[12632]), .I1(ram[12624]), .I2(ram[12616]), .I3(
        ram[12608]), .S0(n27054), .S1(n26579), .ZN(n21139) );
  MUX41 U9934 ( .I0(ram[12760]), .I1(ram[12752]), .I2(ram[12744]), .I3(
        ram[12736]), .S0(n27054), .S1(n26579), .ZN(n21144) );
  MUX41 U9935 ( .I0(ram[12504]), .I1(ram[12496]), .I2(ram[12488]), .I3(
        ram[12480]), .S0(n27053), .S1(n26578), .ZN(n21134) );
  MUX41 U9936 ( .I0(ram[12376]), .I1(ram[12368]), .I2(ram[12360]), .I3(
        ram[12352]), .S0(n27053), .S1(n26578), .ZN(n21129) );
  MUX41 U9937 ( .I0(n20749), .I1(n20750), .I2(n20751), .I3(n20752), .S0(
        n26196), .S1(n26314), .ZN(n20748) );
  MUX41 U9938 ( .I0(ram[3384]), .I1(ram[3376]), .I2(ram[3368]), .I3(
        ram[3360]), .S0(n27032), .S1(n26557), .ZN(n20750) );
  MUX41 U9939 ( .I0(ram[3352]), .I1(ram[3344]), .I2(ram[3336]), .I3(
        ram[3328]), .S0(n27031), .S1(n26556), .ZN(n20752) );
  MUX41 U9940 ( .I0(ram[3448]), .I1(ram[3440]), .I2(ram[3432]), .I3(
        ram[3424]), .S0(n27032), .S1(n26557), .ZN(n20749) );
  MUX41 U9941 ( .I0(n20769), .I1(n20770), .I2(n20771), .I3(n20772), .S0(
        n26196), .S1(n26314), .ZN(n20768) );
  MUX41 U9942 ( .I0(ram[3896]), .I1(ram[3888]), .I2(ram[3880]), .I3(
        ram[3872]), .S0(n27033), .S1(n26558), .ZN(n20770) );
  MUX41 U9943 ( .I0(ram[3864]), .I1(ram[3856]), .I2(ram[3848]), .I3(
        ram[3840]), .S0(n27033), .S1(n26558), .ZN(n20772) );
  MUX41 U9944 ( .I0(ram[3960]), .I1(ram[3952]), .I2(ram[3944]), .I3(
        ram[3936]), .S0(n27033), .S1(n26558), .ZN(n20769) );
  MUX41 U9945 ( .I0(n20709), .I1(n20710), .I2(n20711), .I3(n20712), .S0(
        n26195), .S1(n26313), .ZN(n20708) );
  MUX41 U9946 ( .I0(ram[2328]), .I1(ram[2320]), .I2(ram[2312]), .I3(
        ram[2304]), .S0(n27029), .S1(n26554), .ZN(n20712) );
  MUX41 U9947 ( .I0(ram[2360]), .I1(ram[2352]), .I2(ram[2344]), .I3(
        ram[2336]), .S0(n27029), .S1(n26554), .ZN(n20710) );
  MUX41 U9948 ( .I0(ram[2424]), .I1(ram[2416]), .I2(ram[2408]), .I3(
        ram[2400]), .S0(n27029), .S1(n26554), .ZN(n20709) );
  MUX41 U9949 ( .I0(n20729), .I1(n20730), .I2(n20731), .I3(n20732), .S0(
        n26195), .S1(n26313), .ZN(n20728) );
  MUX41 U9950 ( .I0(ram[2840]), .I1(ram[2832]), .I2(ram[2824]), .I3(
        ram[2816]), .S0(n27030), .S1(n26555), .ZN(n20732) );
  MUX41 U9951 ( .I0(ram[2872]), .I1(ram[2864]), .I2(ram[2856]), .I3(
        ram[2848]), .S0(n27030), .S1(n26555), .ZN(n20730) );
  MUX41 U9952 ( .I0(ram[2936]), .I1(ram[2928]), .I2(ram[2920]), .I3(
        ram[2912]), .S0(n27030), .S1(n26555), .ZN(n20729) );
  MUX41 U9953 ( .I0(n20664), .I1(n20665), .I2(n20666), .I3(n20667), .S0(
        n26195), .S1(n26313), .ZN(n20663) );
  MUX41 U9954 ( .I0(ram[1336]), .I1(ram[1328]), .I2(ram[1320]), .I3(
        ram[1312]), .S0(n27027), .S1(n26552), .ZN(n20665) );
  MUX41 U9955 ( .I0(ram[1304]), .I1(ram[1296]), .I2(ram[1288]), .I3(
        ram[1280]), .S0(n27027), .S1(n26552), .ZN(n20667) );
  MUX41 U9956 ( .I0(ram[1400]), .I1(ram[1392]), .I2(ram[1384]), .I3(
        ram[1376]), .S0(n27027), .S1(n26552), .ZN(n20664) );
  MUX41 U9957 ( .I0(n20684), .I1(n20685), .I2(n20686), .I3(n20687), .S0(
        n26195), .S1(n26313), .ZN(n20683) );
  MUX41 U9958 ( .I0(ram[1816]), .I1(ram[1808]), .I2(ram[1800]), .I3(
        ram[1792]), .S0(n27028), .S1(n26553), .ZN(n20687) );
  MUX41 U9959 ( .I0(ram[1848]), .I1(ram[1840]), .I2(ram[1832]), .I3(
        ram[1824]), .S0(n27028), .S1(n26553), .ZN(n20685) );
  MUX41 U9960 ( .I0(ram[1912]), .I1(ram[1904]), .I2(ram[1896]), .I3(
        ram[1888]), .S0(n27028), .S1(n26553), .ZN(n20684) );
  MUX41 U9961 ( .I0(ram[7512]), .I1(ram[7504]), .I2(ram[7496]), .I3(
        ram[7488]), .S0(n27041), .S1(n26566), .ZN(n20922) );
  MUX41 U9962 ( .I0(ram[7640]), .I1(ram[7632]), .I2(ram[7624]), .I3(
        ram[7616]), .S0(n27042), .S1(n26567), .ZN(n20927) );
  MUX41 U9963 ( .I0(ram[7384]), .I1(ram[7376]), .I2(ram[7368]), .I3(
        ram[7360]), .S0(n27041), .S1(n26566), .ZN(n20917) );
  MUX41 U9964 ( .I0(ram[7256]), .I1(ram[7248]), .I2(ram[7240]), .I3(
        ram[7232]), .S0(n27041), .S1(n26566), .ZN(n20912) );
  MUX41 U9965 ( .I0(ram[8024]), .I1(ram[8016]), .I2(ram[8008]), .I3(
        ram[8000]), .S0(n27043), .S1(n26568), .ZN(n20942) );
  MUX41 U9966 ( .I0(ram[8152]), .I1(ram[8144]), .I2(ram[8136]), .I3(
        ram[8128]), .S0(n27043), .S1(n26568), .ZN(n20947) );
  MUX41 U9967 ( .I0(ram[7896]), .I1(ram[7888]), .I2(ram[7880]), .I3(
        ram[7872]), .S0(n27042), .S1(n26567), .ZN(n20937) );
  MUX41 U9968 ( .I0(ram[7768]), .I1(ram[7760]), .I2(ram[7752]), .I3(
        ram[7744]), .S0(n27042), .S1(n26567), .ZN(n20932) );
  MUX41 U9969 ( .I0(ram[6488]), .I1(ram[6480]), .I2(ram[6472]), .I3(
        ram[6464]), .S0(n27039), .S1(n26564), .ZN(n20882) );
  MUX41 U9970 ( .I0(ram[6616]), .I1(ram[6608]), .I2(ram[6600]), .I3(
        ram[6592]), .S0(n27039), .S1(n26564), .ZN(n20887) );
  MUX41 U9971 ( .I0(ram[6360]), .I1(ram[6352]), .I2(ram[6344]), .I3(
        ram[6336]), .S0(n27039), .S1(n26564), .ZN(n20877) );
  MUX41 U9972 ( .I0(ram[6232]), .I1(ram[6224]), .I2(ram[6216]), .I3(
        ram[6208]), .S0(n27038), .S1(n26563), .ZN(n20872) );
  MUX41 U9973 ( .I0(ram[7000]), .I1(ram[6992]), .I2(ram[6984]), .I3(
        ram[6976]), .S0(n27040), .S1(n26565), .ZN(n20902) );
  MUX41 U9974 ( .I0(ram[7128]), .I1(ram[7120]), .I2(ram[7112]), .I3(
        ram[7104]), .S0(n27041), .S1(n26566), .ZN(n20907) );
  MUX41 U9975 ( .I0(ram[6872]), .I1(ram[6864]), .I2(ram[6856]), .I3(
        ram[6848]), .S0(n27040), .S1(n26565), .ZN(n20897) );
  MUX41 U9976 ( .I0(ram[5464]), .I1(ram[5456]), .I2(ram[5448]), .I3(
        ram[5440]), .S0(n27037), .S1(n26562), .ZN(n20837) );
  MUX41 U9977 ( .I0(ram[5592]), .I1(ram[5584]), .I2(ram[5576]), .I3(
        ram[5568]), .S0(n27037), .S1(n26562), .ZN(n20842) );
  MUX41 U9978 ( .I0(ram[5336]), .I1(ram[5328]), .I2(ram[5320]), .I3(
        ram[5312]), .S0(n27036), .S1(n26561), .ZN(n20832) );
  MUX41 U9979 ( .I0(ram[5208]), .I1(ram[5200]), .I2(ram[5192]), .I3(
        ram[5184]), .S0(n27036), .S1(n26561), .ZN(n20827) );
  MUX41 U9980 ( .I0(ram[5976]), .I1(ram[5968]), .I2(ram[5960]), .I3(
        ram[5952]), .S0(n27038), .S1(n26563), .ZN(n20857) );
  MUX41 U9981 ( .I0(ram[6104]), .I1(ram[6096]), .I2(ram[6088]), .I3(
        ram[6080]), .S0(n27038), .S1(n26563), .ZN(n20862) );
  MUX41 U9982 ( .I0(ram[5848]), .I1(ram[5840]), .I2(ram[5832]), .I3(
        ram[5824]), .S0(n27037), .S1(n26562), .ZN(n20852) );
  MUX41 U9983 ( .I0(ram[5720]), .I1(ram[5712]), .I2(ram[5704]), .I3(
        ram[5696]), .S0(n27037), .S1(n26562), .ZN(n20847) );
  MUX41 U9984 ( .I0(ram[4440]), .I1(ram[4432]), .I2(ram[4424]), .I3(
        ram[4416]), .S0(n27034), .S1(n26559), .ZN(n20797) );
  MUX41 U9985 ( .I0(ram[4568]), .I1(ram[4560]), .I2(ram[4552]), .I3(
        ram[4544]), .S0(n27034), .S1(n26559), .ZN(n20802) );
  MUX41 U9986 ( .I0(ram[4952]), .I1(ram[4944]), .I2(ram[4936]), .I3(
        ram[4928]), .S0(n27035), .S1(n26560), .ZN(n20817) );
  MUX41 U9987 ( .I0(ram[11608]), .I1(ram[11600]), .I2(ram[11592]), .I3(
        ram[11584]), .S0(n27051), .S1(n26576), .ZN(n21093) );
  MUX41 U9988 ( .I0(ram[11736]), .I1(ram[11728]), .I2(ram[11720]), .I3(
        ram[11712]), .S0(n27052), .S1(n26577), .ZN(n21098) );
  MUX41 U9989 ( .I0(ram[11480]), .I1(ram[11472]), .I2(ram[11464]), .I3(
        ram[11456]), .S0(n27051), .S1(n26576), .ZN(n21088) );
  MUX41 U9990 ( .I0(ram[11352]), .I1(ram[11344]), .I2(ram[11336]), .I3(
        ram[11328]), .S0(n27051), .S1(n26576), .ZN(n21083) );
  MUX41 U9991 ( .I0(ram[12120]), .I1(ram[12112]), .I2(ram[12104]), .I3(
        ram[12096]), .S0(n27053), .S1(n26578), .ZN(n21113) );
  MUX41 U9992 ( .I0(ram[12248]), .I1(ram[12240]), .I2(ram[12232]), .I3(
        ram[12224]), .S0(n27053), .S1(n26578), .ZN(n21118) );
  MUX41 U9993 ( .I0(ram[11992]), .I1(ram[11984]), .I2(ram[11976]), .I3(
        ram[11968]), .S0(n27052), .S1(n26577), .ZN(n21108) );
  MUX41 U9994 ( .I0(ram[11864]), .I1(ram[11856]), .I2(ram[11848]), .I3(
        ram[11840]), .S0(n27052), .S1(n26577), .ZN(n21103) );
  MUX41 U9995 ( .I0(ram[10584]), .I1(ram[10576]), .I2(ram[10568]), .I3(
        ram[10560]), .S0(n27049), .S1(n26574), .ZN(n21053) );
  MUX41 U9996 ( .I0(ram[10712]), .I1(ram[10704]), .I2(ram[10696]), .I3(
        ram[10688]), .S0(n27049), .S1(n26574), .ZN(n21058) );
  MUX41 U9997 ( .I0(ram[10456]), .I1(ram[10448]), .I2(ram[10440]), .I3(
        ram[10432]), .S0(n27049), .S1(n26574), .ZN(n21048) );
  MUX41 U9998 ( .I0(ram[10328]), .I1(ram[10320]), .I2(ram[10312]), .I3(
        ram[10304]), .S0(n27048), .S1(n26573), .ZN(n21043) );
  MUX41 U9999 ( .I0(ram[11096]), .I1(ram[11088]), .I2(ram[11080]), .I3(
        ram[11072]), .S0(n27050), .S1(n26575), .ZN(n21073) );
  MUX41 U10000 ( .I0(ram[11224]), .I1(ram[11216]), .I2(ram[11208]), .I3(
        ram[11200]), .S0(n27050), .S1(n26575), .ZN(n21078) );
  MUX41 U10001 ( .I0(ram[9560]), .I1(ram[9552]), .I2(ram[9544]), .I3(
        ram[9536]), .S0(n27046), .S1(n26571), .ZN(n21008) );
  MUX41 U10002 ( .I0(ram[9688]), .I1(ram[9680]), .I2(ram[9672]), .I3(
        ram[9664]), .S0(n27047), .S1(n26572), .ZN(n21013) );
  MUX41 U10003 ( .I0(ram[9432]), .I1(ram[9424]), .I2(ram[9416]), .I3(
        ram[9408]), .S0(n27046), .S1(n26571), .ZN(n21003) );
  MUX41 U10004 ( .I0(ram[9304]), .I1(ram[9296]), .I2(ram[9288]), .I3(
        ram[9280]), .S0(n27046), .S1(n26571), .ZN(n20998) );
  MUX41 U10005 ( .I0(ram[10072]), .I1(ram[10064]), .I2(ram[10056]), .I3(
        ram[10048]), .S0(n27048), .S1(n26573), .ZN(n21028) );
  MUX41 U10006 ( .I0(ram[10200]), .I1(ram[10192]), .I2(ram[10184]), .I3(
        ram[10176]), .S0(n27048), .S1(n26573), .ZN(n21033) );
  MUX41 U10007 ( .I0(ram[9944]), .I1(ram[9936]), .I2(ram[9928]), .I3(
        ram[9920]), .S0(n27047), .S1(n26572), .ZN(n21023) );
  MUX41 U10008 ( .I0(ram[9816]), .I1(ram[9808]), .I2(ram[9800]), .I3(
        ram[9792]), .S0(n27047), .S1(n26572), .ZN(n21018) );
  MUX41 U10009 ( .I0(ram[8536]), .I1(ram[8528]), .I2(ram[8520]), .I3(
        ram[8512]), .S0(n27044), .S1(n26569), .ZN(n20968) );
  MUX41 U10010 ( .I0(ram[8664]), .I1(ram[8656]), .I2(ram[8648]), .I3(
        ram[8640]), .S0(n27044), .S1(n26569), .ZN(n20973) );
  MUX41 U10011 ( .I0(ram[8408]), .I1(ram[8400]), .I2(ram[8392]), .I3(
        ram[8384]), .S0(n27044), .S1(n26569), .ZN(n20963) );
  MUX41 U10012 ( .I0(ram[9048]), .I1(ram[9040]), .I2(ram[9032]), .I3(
        ram[9024]), .S0(n27045), .S1(n26570), .ZN(n20988) );
  MUX41 U10013 ( .I0(ram[9176]), .I1(ram[9168]), .I2(ram[9160]), .I3(
        ram[9152]), .S0(n27045), .S1(n26570), .ZN(n20993) );
  MUX41 U10014 ( .I0(ram[15705]), .I1(ram[15697]), .I2(ram[15689]), .I3(
        ram[15681]), .S0(n27101), .S1(n26626), .ZN(n21948) );
  MUX41 U10015 ( .I0(ram[15833]), .I1(ram[15825]), .I2(ram[15817]), .I3(
        ram[15809]), .S0(n27101), .S1(n26626), .ZN(n21953) );
  MUX41 U10016 ( .I0(ram[15577]), .I1(ram[15569]), .I2(ram[15561]), .I3(
        ram[15553]), .S0(n27100), .S1(n26625), .ZN(n21943) );
  MUX41 U10017 ( .I0(ram[15449]), .I1(ram[15441]), .I2(ram[15433]), .I3(
        ram[15425]), .S0(n27100), .S1(n26625), .ZN(n21938) );
  MUX41 U10018 ( .I0(ram[16217]), .I1(ram[16209]), .I2(ram[16201]), .I3(
        ram[16193]), .S0(n27102), .S1(n26627), .ZN(n21968) );
  MUX41 U10019 ( .I0(ram[16345]), .I1(ram[16337]), .I2(ram[16329]), .I3(
        ram[16321]), .S0(n27102), .S1(n26627), .ZN(n21973) );
  MUX41 U10020 ( .I0(ram[16089]), .I1(ram[16081]), .I2(ram[16073]), .I3(
        ram[16065]), .S0(n27101), .S1(n26626), .ZN(n21963) );
  MUX41 U10021 ( .I0(ram[15961]), .I1(ram[15953]), .I2(ram[15945]), .I3(
        ram[15937]), .S0(n27101), .S1(n26626), .ZN(n21958) );
  MUX41 U10022 ( .I0(ram[15193]), .I1(ram[15185]), .I2(ram[15177]), .I3(
        ram[15169]), .S0(n27099), .S1(n26624), .ZN(n21928) );
  MUX41 U10023 ( .I0(ram[15321]), .I1(ram[15313]), .I2(ram[15305]), .I3(
        ram[15297]), .S0(n27100), .S1(n26625), .ZN(n21933) );
  MUX41 U10024 ( .I0(ram[15065]), .I1(ram[15057]), .I2(ram[15049]), .I3(
        ram[15041]), .S0(n27099), .S1(n26624), .ZN(n21923) );
  MUX41 U10025 ( .I0(ram[14937]), .I1(ram[14929]), .I2(ram[14921]), .I3(
        ram[14913]), .S0(n27099), .S1(n26624), .ZN(n21918) );
  MUX41 U10026 ( .I0(ram[14681]), .I1(ram[14673]), .I2(ram[14665]), .I3(
        ram[14657]), .S0(n27098), .S1(n26623), .ZN(n21908) );
  MUX41 U10027 ( .I0(ram[14809]), .I1(ram[14801]), .I2(ram[14793]), .I3(
        ram[14785]), .S0(n27098), .S1(n26623), .ZN(n21913) );
  MUX41 U10028 ( .I0(ram[14553]), .I1(ram[14545]), .I2(ram[14537]), .I3(
        ram[14529]), .S0(n27098), .S1(n26623), .ZN(n21903) );
  MUX41 U10029 ( .I0(ram[14425]), .I1(ram[14417]), .I2(ram[14409]), .I3(
        ram[14401]), .S0(n27097), .S1(n26622), .ZN(n21898) );
  MUX41 U10030 ( .I0(ram[13657]), .I1(ram[13649]), .I2(ram[13641]), .I3(
        ram[13633]), .S0(n27096), .S1(n26621), .ZN(n21863) );
  MUX41 U10031 ( .I0(ram[13785]), .I1(ram[13777]), .I2(ram[13769]), .I3(
        ram[13761]), .S0(n27096), .S1(n26621), .ZN(n21868) );
  MUX41 U10032 ( .I0(ram[13529]), .I1(ram[13521]), .I2(ram[13513]), .I3(
        ram[13505]), .S0(n27095), .S1(n26620), .ZN(n21858) );
  MUX41 U10033 ( .I0(ram[13401]), .I1(ram[13393]), .I2(ram[13385]), .I3(
        ram[13377]), .S0(n27095), .S1(n26620), .ZN(n21853) );
  MUX41 U10034 ( .I0(ram[14169]), .I1(ram[14161]), .I2(ram[14153]), .I3(
        ram[14145]), .S0(n27097), .S1(n26622), .ZN(n21883) );
  MUX41 U10035 ( .I0(ram[14297]), .I1(ram[14289]), .I2(ram[14281]), .I3(
        ram[14273]), .S0(n27097), .S1(n26622), .ZN(n21888) );
  MUX41 U10036 ( .I0(ram[14041]), .I1(ram[14033]), .I2(ram[14025]), .I3(
        ram[14017]), .S0(n27097), .S1(n26622), .ZN(n21878) );
  MUX41 U10037 ( .I0(ram[13913]), .I1(ram[13905]), .I2(ram[13897]), .I3(
        ram[13889]), .S0(n27096), .S1(n26621), .ZN(n21873) );
  MUX41 U10038 ( .I0(ram[13145]), .I1(ram[13137]), .I2(ram[13129]), .I3(
        ram[13121]), .S0(n27094), .S1(n26619), .ZN(n21843) );
  MUX41 U10039 ( .I0(ram[13273]), .I1(ram[13265]), .I2(ram[13257]), .I3(
        ram[13249]), .S0(n27095), .S1(n26620), .ZN(n21848) );
  MUX41 U10040 ( .I0(ram[13017]), .I1(ram[13009]), .I2(ram[13001]), .I3(
        ram[12993]), .S0(n27094), .S1(n26619), .ZN(n21838) );
  MUX41 U10041 ( .I0(ram[12889]), .I1(ram[12881]), .I2(ram[12873]), .I3(
        ram[12865]), .S0(n27094), .S1(n26619), .ZN(n21833) );
  MUX41 U10042 ( .I0(ram[12633]), .I1(ram[12625]), .I2(ram[12617]), .I3(
        ram[12609]), .S0(n27093), .S1(n26618), .ZN(n21823) );
  MUX41 U10043 ( .I0(ram[12761]), .I1(ram[12753]), .I2(ram[12745]), .I3(
        ram[12737]), .S0(n27093), .S1(n26618), .ZN(n21828) );
  MUX41 U10044 ( .I0(ram[12505]), .I1(ram[12497]), .I2(ram[12489]), .I3(
        ram[12481]), .S0(n27093), .S1(n26618), .ZN(n21818) );
  MUX41 U10045 ( .I0(ram[12377]), .I1(ram[12369]), .I2(ram[12361]), .I3(
        ram[12353]), .S0(n27093), .S1(n26618), .ZN(n21813) );
  MUX41 U10046 ( .I0(n21433), .I1(n21434), .I2(n21435), .I3(n21436), .S0(
        n26206), .S1(n26324), .ZN(n21432) );
  MUX41 U10047 ( .I0(ram[3385]), .I1(ram[3377]), .I2(ram[3369]), .I3(
        ram[3361]), .S0(n27071), .S1(n26596), .ZN(n21434) );
  MUX41 U10048 ( .I0(ram[3353]), .I1(ram[3345]), .I2(ram[3337]), .I3(
        ram[3329]), .S0(n27071), .S1(n26596), .ZN(n21436) );
  MUX41 U10049 ( .I0(ram[3449]), .I1(ram[3441]), .I2(ram[3433]), .I3(
        ram[3425]), .S0(n27071), .S1(n26596), .ZN(n21433) );
  MUX41 U10050 ( .I0(n21453), .I1(n21454), .I2(n21455), .I3(n21456), .S0(
        n26206), .S1(n26324), .ZN(n21452) );
  MUX41 U10051 ( .I0(ram[3897]), .I1(ram[3889]), .I2(ram[3881]), .I3(
        ram[3873]), .S0(n27072), .S1(n26597), .ZN(n21454) );
  MUX41 U10052 ( .I0(ram[3865]), .I1(ram[3857]), .I2(ram[3849]), .I3(
        ram[3841]), .S0(n27072), .S1(n26597), .ZN(n21456) );
  MUX41 U10053 ( .I0(ram[3961]), .I1(ram[3953]), .I2(ram[3945]), .I3(
        ram[3937]), .S0(n27072), .S1(n26597), .ZN(n21453) );
  MUX41 U10054 ( .I0(n21393), .I1(n21394), .I2(n21395), .I3(n21396), .S0(
        n26205), .S1(n26323), .ZN(n21392) );
  MUX41 U10055 ( .I0(ram[2329]), .I1(ram[2321]), .I2(ram[2313]), .I3(
        ram[2305]), .S0(n27068), .S1(n26593), .ZN(n21396) );
  MUX41 U10056 ( .I0(ram[2361]), .I1(ram[2353]), .I2(ram[2345]), .I3(
        ram[2337]), .S0(n27068), .S1(n26593), .ZN(n21394) );
  MUX41 U10057 ( .I0(ram[2425]), .I1(ram[2417]), .I2(ram[2409]), .I3(
        ram[2401]), .S0(n27069), .S1(n26594), .ZN(n21393) );
  MUX41 U10058 ( .I0(n21413), .I1(n21414), .I2(n21415), .I3(n21416), .S0(
        n26205), .S1(n26323), .ZN(n21412) );
  MUX41 U10059 ( .I0(ram[2841]), .I1(ram[2833]), .I2(ram[2825]), .I3(
        ram[2817]), .S0(n27070), .S1(n26595), .ZN(n21416) );
  MUX41 U10060 ( .I0(ram[2873]), .I1(ram[2865]), .I2(ram[2857]), .I3(
        ram[2849]), .S0(n27070), .S1(n26595), .ZN(n21414) );
  MUX41 U10061 ( .I0(ram[2937]), .I1(ram[2929]), .I2(ram[2921]), .I3(
        ram[2913]), .S0(n27070), .S1(n26595), .ZN(n21413) );
  MUX41 U10062 ( .I0(n21348), .I1(n21349), .I2(n21350), .I3(n21351), .S0(
        n26204), .S1(n26322), .ZN(n21347) );
  MUX41 U10063 ( .I0(ram[1337]), .I1(ram[1329]), .I2(ram[1321]), .I3(
        ram[1313]), .S0(n27066), .S1(n26591), .ZN(n21349) );
  MUX41 U10064 ( .I0(ram[1305]), .I1(ram[1297]), .I2(ram[1289]), .I3(
        ram[1281]), .S0(n27066), .S1(n26591), .ZN(n21351) );
  MUX41 U10065 ( .I0(ram[1401]), .I1(ram[1393]), .I2(ram[1385]), .I3(
        ram[1377]), .S0(n27066), .S1(n26591), .ZN(n21348) );
  MUX41 U10066 ( .I0(n21368), .I1(n21369), .I2(n21370), .I3(n21371), .S0(
        n26205), .S1(n26323), .ZN(n21367) );
  MUX41 U10067 ( .I0(ram[1817]), .I1(ram[1809]), .I2(ram[1801]), .I3(
        ram[1793]), .S0(n27067), .S1(n26592), .ZN(n21371) );
  MUX41 U10068 ( .I0(ram[1849]), .I1(ram[1841]), .I2(ram[1833]), .I3(
        ram[1825]), .S0(n27067), .S1(n26592), .ZN(n21369) );
  MUX41 U10069 ( .I0(ram[1913]), .I1(ram[1905]), .I2(ram[1897]), .I3(
        ram[1889]), .S0(n27067), .S1(n26592), .ZN(n21368) );
  MUX41 U10070 ( .I0(n21308), .I1(n21309), .I2(n21310), .I3(n21311), .S0(
        n26204), .S1(n26322), .ZN(n21307) );
  MUX41 U10071 ( .I0(ram[281]), .I1(ram[273]), .I2(ram[265]), .I3(
        ram[257]), .S0(n27063), .S1(n26588), .ZN(n21311) );
  MUX41 U10072 ( .I0(ram[313]), .I1(ram[305]), .I2(ram[297]), .I3(
        ram[289]), .S0(n27064), .S1(n26589), .ZN(n21309) );
  MUX41 U10073 ( .I0(ram[377]), .I1(ram[369]), .I2(ram[361]), .I3(
        ram[353]), .S0(n27064), .S1(n26589), .ZN(n21308) );
  MUX41 U10074 ( .I0(n21328), .I1(n21329), .I2(n21330), .I3(n21331), .S0(
        n26204), .S1(n26322), .ZN(n21327) );
  MUX41 U10075 ( .I0(ram[793]), .I1(ram[785]), .I2(ram[777]), .I3(
        ram[769]), .S0(n27065), .S1(n26590), .ZN(n21331) );
  MUX41 U10076 ( .I0(ram[825]), .I1(ram[817]), .I2(ram[809]), .I3(
        ram[801]), .S0(n27065), .S1(n26590), .ZN(n21329) );
  MUX41 U10077 ( .I0(ram[889]), .I1(ram[881]), .I2(ram[873]), .I3(
        ram[865]), .S0(n27065), .S1(n26590), .ZN(n21328) );
  MUX41 U10078 ( .I0(ram[7513]), .I1(ram[7505]), .I2(ram[7497]), .I3(
        ram[7489]), .S0(n27081), .S1(n26606), .ZN(n21606) );
  MUX41 U10079 ( .I0(ram[7641]), .I1(ram[7633]), .I2(ram[7625]), .I3(
        ram[7617]), .S0(n27081), .S1(n26606), .ZN(n21611) );
  MUX41 U10080 ( .I0(ram[7385]), .I1(ram[7377]), .I2(ram[7369]), .I3(
        ram[7361]), .S0(n27081), .S1(n26606), .ZN(n21601) );
  MUX41 U10081 ( .I0(ram[7257]), .I1(ram[7249]), .I2(ram[7241]), .I3(
        ram[7233]), .S0(n27080), .S1(n26605), .ZN(n21596) );
  MUX41 U10082 ( .I0(ram[8025]), .I1(ram[8017]), .I2(ram[8009]), .I3(
        ram[8001]), .S0(n27082), .S1(n26607), .ZN(n21626) );
  MUX41 U10083 ( .I0(ram[8153]), .I1(ram[8145]), .I2(ram[8137]), .I3(
        ram[8129]), .S0(n27082), .S1(n26607), .ZN(n21631) );
  MUX41 U10084 ( .I0(ram[7897]), .I1(ram[7889]), .I2(ram[7881]), .I3(
        ram[7873]), .S0(n27082), .S1(n26607), .ZN(n21621) );
  MUX41 U10085 ( .I0(ram[7769]), .I1(ram[7761]), .I2(ram[7753]), .I3(
        ram[7745]), .S0(n27081), .S1(n26606), .ZN(n21616) );
  MUX41 U10086 ( .I0(ram[6489]), .I1(ram[6481]), .I2(ram[6473]), .I3(
        ram[6465]), .S0(n27078), .S1(n26603), .ZN(n21566) );
  MUX41 U10087 ( .I0(ram[6617]), .I1(ram[6609]), .I2(ram[6601]), .I3(
        ram[6593]), .S0(n27079), .S1(n26604), .ZN(n21571) );
  MUX41 U10088 ( .I0(ram[6361]), .I1(ram[6353]), .I2(ram[6345]), .I3(
        ram[6337]), .S0(n27078), .S1(n26603), .ZN(n21561) );
  MUX41 U10089 ( .I0(ram[6233]), .I1(ram[6225]), .I2(ram[6217]), .I3(
        ram[6209]), .S0(n27078), .S1(n26603), .ZN(n21556) );
  MUX41 U10090 ( .I0(ram[7001]), .I1(ram[6993]), .I2(ram[6985]), .I3(
        ram[6977]), .S0(n27080), .S1(n26605), .ZN(n21586) );
  MUX41 U10091 ( .I0(ram[7129]), .I1(ram[7121]), .I2(ram[7113]), .I3(
        ram[7105]), .S0(n27080), .S1(n26605), .ZN(n21591) );
  MUX41 U10092 ( .I0(ram[6873]), .I1(ram[6865]), .I2(ram[6857]), .I3(
        ram[6849]), .S0(n27079), .S1(n26604), .ZN(n21581) );
  MUX41 U10093 ( .I0(ram[5465]), .I1(ram[5457]), .I2(ram[5449]), .I3(
        ram[5441]), .S0(n27076), .S1(n26601), .ZN(n21521) );
  MUX41 U10094 ( .I0(ram[5593]), .I1(ram[5585]), .I2(ram[5577]), .I3(
        ram[5569]), .S0(n27076), .S1(n26601), .ZN(n21526) );
  MUX41 U10095 ( .I0(ram[5337]), .I1(ram[5329]), .I2(ram[5321]), .I3(
        ram[5313]), .S0(n27076), .S1(n26601), .ZN(n21516) );
  MUX41 U10096 ( .I0(ram[5209]), .I1(ram[5201]), .I2(ram[5193]), .I3(
        ram[5185]), .S0(n27075), .S1(n26600), .ZN(n21511) );
  MUX41 U10097 ( .I0(ram[5977]), .I1(ram[5969]), .I2(ram[5961]), .I3(
        ram[5953]), .S0(n27077), .S1(n26602), .ZN(n21541) );
  MUX41 U10098 ( .I0(ram[6105]), .I1(ram[6097]), .I2(ram[6089]), .I3(
        ram[6081]), .S0(n27077), .S1(n26602), .ZN(n21546) );
  MUX41 U10099 ( .I0(ram[5849]), .I1(ram[5841]), .I2(ram[5833]), .I3(
        ram[5825]), .S0(n27077), .S1(n26602), .ZN(n21536) );
  MUX41 U10100 ( .I0(ram[5721]), .I1(ram[5713]), .I2(ram[5705]), .I3(
        ram[5697]), .S0(n27077), .S1(n26602), .ZN(n21531) );
  MUX41 U10101 ( .I0(ram[4441]), .I1(ram[4433]), .I2(ram[4425]), .I3(
        ram[4417]), .S0(n27073), .S1(n26598), .ZN(n21481) );
  MUX41 U10102 ( .I0(ram[4569]), .I1(ram[4561]), .I2(ram[4553]), .I3(
        ram[4545]), .S0(n27074), .S1(n26599), .ZN(n21486) );
  MUX41 U10103 ( .I0(ram[4953]), .I1(ram[4945]), .I2(ram[4937]), .I3(
        ram[4929]), .S0(n27075), .S1(n26600), .ZN(n21501) );
  MUX41 U10104 ( .I0(ram[11609]), .I1(ram[11601]), .I2(ram[11593]), .I3(
        ram[11585]), .S0(n27091), .S1(n26616), .ZN(n21777) );
  MUX41 U10105 ( .I0(ram[11737]), .I1(ram[11729]), .I2(ram[11721]), .I3(
        ram[11713]), .S0(n27091), .S1(n26616), .ZN(n21782) );
  MUX41 U10106 ( .I0(ram[11481]), .I1(ram[11473]), .I2(ram[11465]), .I3(
        ram[11457]), .S0(n27090), .S1(n26615), .ZN(n21772) );
  MUX41 U10107 ( .I0(ram[11353]), .I1(ram[11345]), .I2(ram[11337]), .I3(
        ram[11329]), .S0(n27090), .S1(n26615), .ZN(n21767) );
  MUX41 U10108 ( .I0(ram[12121]), .I1(ram[12113]), .I2(ram[12105]), .I3(
        ram[12097]), .S0(n27092), .S1(n26617), .ZN(n21797) );
  MUX41 U10109 ( .I0(ram[12249]), .I1(ram[12241]), .I2(ram[12233]), .I3(
        ram[12225]), .S0(n27092), .S1(n26617), .ZN(n21802) );
  MUX41 U10110 ( .I0(ram[11993]), .I1(ram[11985]), .I2(ram[11977]), .I3(
        ram[11969]), .S0(n27092), .S1(n26617), .ZN(n21792) );
  MUX41 U10111 ( .I0(ram[11865]), .I1(ram[11857]), .I2(ram[11849]), .I3(
        ram[11841]), .S0(n27091), .S1(n26616), .ZN(n21787) );
  MUX41 U10112 ( .I0(ram[10585]), .I1(ram[10577]), .I2(ram[10569]), .I3(
        ram[10561]), .S0(n27088), .S1(n26613), .ZN(n21737) );
  MUX41 U10113 ( .I0(ram[10713]), .I1(ram[10705]), .I2(ram[10697]), .I3(
        ram[10689]), .S0(n27089), .S1(n26614), .ZN(n21742) );
  MUX41 U10114 ( .I0(ram[10457]), .I1(ram[10449]), .I2(ram[10441]), .I3(
        ram[10433]), .S0(n27088), .S1(n26613), .ZN(n21732) );
  MUX41 U10115 ( .I0(ram[10329]), .I1(ram[10321]), .I2(ram[10313]), .I3(
        ram[10305]), .S0(n27088), .S1(n26613), .ZN(n21727) );
  MUX41 U10116 ( .I0(ram[11097]), .I1(ram[11089]), .I2(ram[11081]), .I3(
        ram[11073]), .S0(n27089), .S1(n26614), .ZN(n21757) );
  MUX41 U10117 ( .I0(ram[11225]), .I1(ram[11217]), .I2(ram[11209]), .I3(
        ram[11201]), .S0(n27090), .S1(n26615), .ZN(n21762) );
  MUX41 U10118 ( .I0(ram[9561]), .I1(ram[9553]), .I2(ram[9545]), .I3(
        ram[9537]), .S0(n27086), .S1(n26611), .ZN(n21692) );
  MUX41 U10119 ( .I0(ram[9689]), .I1(ram[9681]), .I2(ram[9673]), .I3(
        ram[9665]), .S0(n27086), .S1(n26611), .ZN(n21697) );
  MUX41 U10120 ( .I0(ram[9433]), .I1(ram[9425]), .I2(ram[9417]), .I3(
        ram[9409]), .S0(n27085), .S1(n26610), .ZN(n21687) );
  MUX41 U10121 ( .I0(ram[9305]), .I1(ram[9297]), .I2(ram[9289]), .I3(
        ram[9281]), .S0(n27085), .S1(n26610), .ZN(n21682) );
  MUX41 U10122 ( .I0(ram[10073]), .I1(ram[10065]), .I2(ram[10057]), .I3(
        ram[10049]), .S0(n27087), .S1(n26612), .ZN(n21712) );
  MUX41 U10123 ( .I0(ram[10201]), .I1(ram[10193]), .I2(ram[10185]), .I3(
        ram[10177]), .S0(n27087), .S1(n26612), .ZN(n21717) );
  MUX41 U10124 ( .I0(ram[9945]), .I1(ram[9937]), .I2(ram[9929]), .I3(
        ram[9921]), .S0(n27087), .S1(n26612), .ZN(n21707) );
  MUX41 U10125 ( .I0(ram[9817]), .I1(ram[9809]), .I2(ram[9801]), .I3(
        ram[9793]), .S0(n27086), .S1(n26611), .ZN(n21702) );
  MUX41 U10126 ( .I0(ram[8537]), .I1(ram[8529]), .I2(ram[8521]), .I3(
        ram[8513]), .S0(n27083), .S1(n26608), .ZN(n21652) );
  MUX41 U10127 ( .I0(ram[8665]), .I1(ram[8657]), .I2(ram[8649]), .I3(
        ram[8641]), .S0(n27084), .S1(n26609), .ZN(n21657) );
  MUX41 U10128 ( .I0(ram[8409]), .I1(ram[8401]), .I2(ram[8393]), .I3(
        ram[8385]), .S0(n27083), .S1(n26608), .ZN(n21647) );
  MUX41 U10129 ( .I0(ram[9049]), .I1(ram[9041]), .I2(ram[9033]), .I3(
        ram[9025]), .S0(n27085), .S1(n26610), .ZN(n21672) );
  MUX41 U10130 ( .I0(ram[9177]), .I1(ram[9169]), .I2(ram[9161]), .I3(
        ram[9153]), .S0(n27085), .S1(n26610), .ZN(n21677) );
  MUX41 U10131 ( .I0(ram[15706]), .I1(ram[15698]), .I2(ram[15690]), .I3(
        ram[15682]), .S0(n27140), .S1(n26665), .ZN(n22632) );
  MUX41 U10132 ( .I0(ram[15834]), .I1(ram[15826]), .I2(ram[15818]), .I3(
        ram[15810]), .S0(n27140), .S1(n26665), .ZN(n22637) );
  MUX41 U10133 ( .I0(ram[15578]), .I1(ram[15570]), .I2(ram[15562]), .I3(
        ram[15554]), .S0(n27140), .S1(n26665), .ZN(n22627) );
  MUX41 U10134 ( .I0(ram[15450]), .I1(ram[15442]), .I2(ram[15434]), .I3(
        ram[15426]), .S0(n27139), .S1(n26664), .ZN(n22622) );
  MUX41 U10135 ( .I0(ram[16218]), .I1(ram[16210]), .I2(ram[16202]), .I3(
        ram[16194]), .S0(n27141), .S1(n26666), .ZN(n22652) );
  MUX41 U10136 ( .I0(ram[16346]), .I1(ram[16338]), .I2(ram[16330]), .I3(
        ram[16322]), .S0(n27141), .S1(n26666), .ZN(n22657) );
  MUX41 U10137 ( .I0(ram[16090]), .I1(ram[16082]), .I2(ram[16074]), .I3(
        ram[16066]), .S0(n27141), .S1(n26666), .ZN(n22647) );
  MUX41 U10138 ( .I0(ram[15962]), .I1(ram[15954]), .I2(ram[15946]), .I3(
        ram[15938]), .S0(n27141), .S1(n26666), .ZN(n22642) );
  MUX41 U10139 ( .I0(ram[15194]), .I1(ram[15186]), .I2(ram[15178]), .I3(
        ram[15170]), .S0(n27139), .S1(n26664), .ZN(n22612) );
  MUX41 U10140 ( .I0(ram[15322]), .I1(ram[15314]), .I2(ram[15306]), .I3(
        ram[15298]), .S0(n27139), .S1(n26664), .ZN(n22617) );
  MUX41 U10141 ( .I0(ram[15066]), .I1(ram[15058]), .I2(ram[15050]), .I3(
        ram[15042]), .S0(n27138), .S1(n26663), .ZN(n22607) );
  MUX41 U10142 ( .I0(ram[14938]), .I1(ram[14930]), .I2(ram[14922]), .I3(
        ram[14914]), .S0(n27138), .S1(n26663), .ZN(n22602) );
  MUX41 U10143 ( .I0(ram[14682]), .I1(ram[14674]), .I2(ram[14666]), .I3(
        ram[14658]), .S0(n27137), .S1(n26662), .ZN(n22592) );
  MUX41 U10144 ( .I0(ram[14810]), .I1(ram[14802]), .I2(ram[14794]), .I3(
        ram[14786]), .S0(n27138), .S1(n26663), .ZN(n22597) );
  MUX41 U10145 ( .I0(ram[14554]), .I1(ram[14546]), .I2(ram[14538]), .I3(
        ram[14530]), .S0(n27137), .S1(n26662), .ZN(n22587) );
  MUX41 U10146 ( .I0(ram[14426]), .I1(ram[14418]), .I2(ram[14410]), .I3(
        ram[14402]), .S0(n27137), .S1(n26662), .ZN(n22582) );
  MUX41 U10147 ( .I0(ram[13658]), .I1(ram[13650]), .I2(ram[13642]), .I3(
        ram[13634]), .S0(n27135), .S1(n26660), .ZN(n22547) );
  MUX41 U10148 ( .I0(ram[13786]), .I1(ram[13778]), .I2(ram[13770]), .I3(
        ram[13762]), .S0(n27135), .S1(n26660), .ZN(n22552) );
  MUX41 U10149 ( .I0(ram[13530]), .I1(ram[13522]), .I2(ram[13514]), .I3(
        ram[13506]), .S0(n27135), .S1(n26660), .ZN(n22542) );
  MUX41 U10150 ( .I0(ram[13402]), .I1(ram[13394]), .I2(ram[13386]), .I3(
        ram[13378]), .S0(n27134), .S1(n26659), .ZN(n22537) );
  MUX41 U10151 ( .I0(ram[14170]), .I1(ram[14162]), .I2(ram[14154]), .I3(
        ram[14146]), .S0(n27136), .S1(n26661), .ZN(n22567) );
  MUX41 U10152 ( .I0(ram[14298]), .I1(ram[14290]), .I2(ram[14282]), .I3(
        ram[14274]), .S0(n27137), .S1(n26662), .ZN(n22572) );
  MUX41 U10153 ( .I0(ram[14042]), .I1(ram[14034]), .I2(ram[14026]), .I3(
        ram[14018]), .S0(n27136), .S1(n26661), .ZN(n22562) );
  MUX41 U10154 ( .I0(ram[13914]), .I1(ram[13906]), .I2(ram[13898]), .I3(
        ram[13890]), .S0(n27136), .S1(n26661), .ZN(n22557) );
  MUX41 U10155 ( .I0(ram[13146]), .I1(ram[13138]), .I2(ram[13130]), .I3(
        ram[13122]), .S0(n27134), .S1(n26659), .ZN(n22527) );
  MUX41 U10156 ( .I0(ram[13274]), .I1(ram[13266]), .I2(ram[13258]), .I3(
        ram[13250]), .S0(n27134), .S1(n26659), .ZN(n22532) );
  MUX41 U10157 ( .I0(ram[13018]), .I1(ram[13010]), .I2(ram[13002]), .I3(
        ram[12994]), .S0(n27133), .S1(n26658), .ZN(n22522) );
  MUX41 U10158 ( .I0(ram[12890]), .I1(ram[12882]), .I2(ram[12874]), .I3(
        ram[12866]), .S0(n27133), .S1(n26658), .ZN(n22517) );
  MUX41 U10159 ( .I0(ram[12634]), .I1(ram[12626]), .I2(ram[12618]), .I3(
        ram[12610]), .S0(n27133), .S1(n26658), .ZN(n22507) );
  MUX41 U10160 ( .I0(ram[12762]), .I1(ram[12754]), .I2(ram[12746]), .I3(
        ram[12738]), .S0(n27133), .S1(n26658), .ZN(n22512) );
  MUX41 U10161 ( .I0(ram[12506]), .I1(ram[12498]), .I2(ram[12490]), .I3(
        ram[12482]), .S0(n27132), .S1(n26657), .ZN(n22502) );
  MUX41 U10162 ( .I0(ram[12378]), .I1(ram[12370]), .I2(ram[12362]), .I3(
        ram[12354]), .S0(n27132), .S1(n26657), .ZN(n22497) );
  MUX41 U10163 ( .I0(n22117), .I1(n22118), .I2(n22119), .I3(n22120), .S0(
        n26215), .S1(n26333), .ZN(n22116) );
  MUX41 U10164 ( .I0(ram[3386]), .I1(ram[3378]), .I2(ram[3370]), .I3(
        ram[3362]), .S0(n27110), .S1(n26635), .ZN(n22118) );
  MUX41 U10165 ( .I0(ram[3354]), .I1(ram[3346]), .I2(ram[3338]), .I3(
        ram[3330]), .S0(n27110), .S1(n26635), .ZN(n22120) );
  MUX41 U10166 ( .I0(ram[3450]), .I1(ram[3442]), .I2(ram[3434]), .I3(
        ram[3426]), .S0(n27110), .S1(n26635), .ZN(n22117) );
  MUX41 U10167 ( .I0(n22137), .I1(n22138), .I2(n22139), .I3(n22140), .S0(
        n26216), .S1(n26334), .ZN(n22136) );
  MUX41 U10168 ( .I0(ram[3898]), .I1(ram[3890]), .I2(ram[3882]), .I3(
        ram[3874]), .S0(n27112), .S1(n26637), .ZN(n22138) );
  MUX41 U10169 ( .I0(ram[3866]), .I1(ram[3858]), .I2(ram[3850]), .I3(
        ram[3842]), .S0(n27111), .S1(n26636), .ZN(n22140) );
  MUX41 U10170 ( .I0(ram[3962]), .I1(ram[3954]), .I2(ram[3946]), .I3(
        ram[3938]), .S0(n27112), .S1(n26637), .ZN(n22137) );
  MUX41 U10171 ( .I0(n22077), .I1(n22078), .I2(n22079), .I3(n22080), .S0(
        n26215), .S1(n26333), .ZN(n22076) );
  MUX41 U10172 ( .I0(ram[2330]), .I1(ram[2322]), .I2(ram[2314]), .I3(
        ram[2306]), .S0(n27108), .S1(n26633), .ZN(n22080) );
  MUX41 U10173 ( .I0(ram[2362]), .I1(ram[2354]), .I2(ram[2346]), .I3(
        ram[2338]), .S0(n27108), .S1(n26633), .ZN(n22078) );
  MUX41 U10174 ( .I0(ram[2426]), .I1(ram[2418]), .I2(ram[2410]), .I3(
        ram[2402]), .S0(n27108), .S1(n26633), .ZN(n22077) );
  MUX41 U10175 ( .I0(n22097), .I1(n22098), .I2(n22099), .I3(n22100), .S0(
        n26215), .S1(n26333), .ZN(n22096) );
  MUX41 U10176 ( .I0(ram[2842]), .I1(ram[2834]), .I2(ram[2826]), .I3(
        ram[2818]), .S0(n27109), .S1(n26634), .ZN(n22100) );
  MUX41 U10177 ( .I0(ram[2874]), .I1(ram[2866]), .I2(ram[2858]), .I3(
        ram[2850]), .S0(n27109), .S1(n26634), .ZN(n22098) );
  MUX41 U10178 ( .I0(ram[2938]), .I1(ram[2930]), .I2(ram[2922]), .I3(
        ram[2914]), .S0(n27109), .S1(n26634), .ZN(n22097) );
  MUX41 U10179 ( .I0(n22032), .I1(n22033), .I2(n22034), .I3(n22035), .S0(
        n26214), .S1(n26332), .ZN(n22031) );
  MUX41 U10180 ( .I0(ram[1338]), .I1(ram[1330]), .I2(ram[1322]), .I3(
        ram[1314]), .S0(n27105), .S1(n26630), .ZN(n22033) );
  MUX41 U10181 ( .I0(ram[1306]), .I1(ram[1298]), .I2(ram[1290]), .I3(
        ram[1282]), .S0(n27105), .S1(n26630), .ZN(n22035) );
  MUX41 U10182 ( .I0(ram[1402]), .I1(ram[1394]), .I2(ram[1386]), .I3(
        ram[1378]), .S0(n27106), .S1(n26631), .ZN(n22032) );
  MUX41 U10183 ( .I0(n22052), .I1(n22053), .I2(n22054), .I3(n22055), .S0(
        n26215), .S1(n26333), .ZN(n22051) );
  MUX41 U10184 ( .I0(ram[1818]), .I1(ram[1810]), .I2(ram[1802]), .I3(
        ram[1794]), .S0(n27107), .S1(n26632), .ZN(n22055) );
  MUX41 U10185 ( .I0(ram[1850]), .I1(ram[1842]), .I2(ram[1834]), .I3(
        ram[1826]), .S0(n27107), .S1(n26632), .ZN(n22053) );
  MUX41 U10186 ( .I0(ram[1914]), .I1(ram[1906]), .I2(ram[1898]), .I3(
        ram[1890]), .S0(n27107), .S1(n26632), .ZN(n22052) );
  MUX41 U10187 ( .I0(n21992), .I1(n21993), .I2(n21994), .I3(n21995), .S0(
        n26214), .S1(n26332), .ZN(n21991) );
  MUX41 U10188 ( .I0(ram[282]), .I1(ram[274]), .I2(ram[266]), .I3(
        ram[258]), .S0(n27103), .S1(n26628), .ZN(n21995) );
  MUX41 U10189 ( .I0(ram[314]), .I1(ram[306]), .I2(ram[298]), .I3(
        ram[290]), .S0(n27103), .S1(n26628), .ZN(n21993) );
  MUX41 U10190 ( .I0(ram[378]), .I1(ram[370]), .I2(ram[362]), .I3(
        ram[354]), .S0(n27103), .S1(n26628), .ZN(n21992) );
  MUX41 U10191 ( .I0(n22012), .I1(n22013), .I2(n22014), .I3(n22015), .S0(
        n26214), .S1(n26332), .ZN(n22011) );
  MUX41 U10192 ( .I0(ram[794]), .I1(ram[786]), .I2(ram[778]), .I3(
        ram[770]), .S0(n27104), .S1(n26629), .ZN(n22015) );
  MUX41 U10193 ( .I0(ram[826]), .I1(ram[818]), .I2(ram[810]), .I3(
        ram[802]), .S0(n27104), .S1(n26629), .ZN(n22013) );
  MUX41 U10194 ( .I0(ram[890]), .I1(ram[882]), .I2(ram[874]), .I3(
        ram[866]), .S0(n27104), .S1(n26629), .ZN(n22012) );
  MUX41 U10195 ( .I0(ram[7514]), .I1(ram[7506]), .I2(ram[7498]), .I3(
        ram[7490]), .S0(n27120), .S1(n26645), .ZN(n22290) );
  MUX41 U10196 ( .I0(ram[7642]), .I1(ram[7634]), .I2(ram[7626]), .I3(
        ram[7618]), .S0(n27121), .S1(n26646), .ZN(n22295) );
  MUX41 U10197 ( .I0(ram[7386]), .I1(ram[7378]), .I2(ram[7370]), .I3(
        ram[7362]), .S0(n27120), .S1(n26645), .ZN(n22285) );
  MUX41 U10198 ( .I0(ram[7258]), .I1(ram[7250]), .I2(ram[7242]), .I3(
        ram[7234]), .S0(n27120), .S1(n26645), .ZN(n22280) );
  MUX41 U10199 ( .I0(ram[8026]), .I1(ram[8018]), .I2(ram[8010]), .I3(
        ram[8002]), .S0(n27121), .S1(n26646), .ZN(n22310) );
  MUX41 U10200 ( .I0(ram[8154]), .I1(ram[8146]), .I2(ram[8138]), .I3(
        ram[8130]), .S0(n27122), .S1(n26647), .ZN(n22315) );
  MUX41 U10201 ( .I0(ram[7898]), .I1(ram[7890]), .I2(ram[7882]), .I3(
        ram[7874]), .S0(n27121), .S1(n26646), .ZN(n22305) );
  MUX41 U10202 ( .I0(ram[7770]), .I1(ram[7762]), .I2(ram[7754]), .I3(
        ram[7746]), .S0(n27121), .S1(n26646), .ZN(n22300) );
  MUX41 U10203 ( .I0(ram[6490]), .I1(ram[6482]), .I2(ram[6474]), .I3(
        ram[6466]), .S0(n27118), .S1(n26643), .ZN(n22250) );
  MUX41 U10204 ( .I0(ram[6618]), .I1(ram[6610]), .I2(ram[6602]), .I3(
        ram[6594]), .S0(n27118), .S1(n26643), .ZN(n22255) );
  MUX41 U10205 ( .I0(ram[6362]), .I1(ram[6354]), .I2(ram[6346]), .I3(
        ram[6338]), .S0(n27117), .S1(n26642), .ZN(n22245) );
  MUX41 U10206 ( .I0(ram[6234]), .I1(ram[6226]), .I2(ram[6218]), .I3(
        ram[6210]), .S0(n27117), .S1(n26642), .ZN(n22240) );
  MUX41 U10207 ( .I0(ram[7002]), .I1(ram[6994]), .I2(ram[6986]), .I3(
        ram[6978]), .S0(n27119), .S1(n26644), .ZN(n22270) );
  MUX41 U10208 ( .I0(ram[7130]), .I1(ram[7122]), .I2(ram[7114]), .I3(
        ram[7106]), .S0(n27119), .S1(n26644), .ZN(n22275) );
  MUX41 U10209 ( .I0(ram[6874]), .I1(ram[6866]), .I2(ram[6858]), .I3(
        ram[6850]), .S0(n27119), .S1(n26644), .ZN(n22265) );
  MUX41 U10210 ( .I0(ram[6746]), .I1(ram[6738]), .I2(ram[6730]), .I3(
        ram[6722]), .S0(n27118), .S1(n26643), .ZN(n22260) );
  MUX41 U10211 ( .I0(ram[5466]), .I1(ram[5458]), .I2(ram[5450]), .I3(
        ram[5442]), .S0(n27115), .S1(n26640), .ZN(n22205) );
  MUX41 U10212 ( .I0(ram[5594]), .I1(ram[5586]), .I2(ram[5578]), .I3(
        ram[5570]), .S0(n27116), .S1(n26641), .ZN(n22210) );
  MUX41 U10213 ( .I0(ram[5338]), .I1(ram[5330]), .I2(ram[5322]), .I3(
        ram[5314]), .S0(n27115), .S1(n26640), .ZN(n22200) );
  MUX41 U10214 ( .I0(ram[5210]), .I1(ram[5202]), .I2(ram[5194]), .I3(
        ram[5186]), .S0(n27115), .S1(n26640), .ZN(n22195) );
  MUX41 U10215 ( .I0(ram[5978]), .I1(ram[5970]), .I2(ram[5962]), .I3(
        ram[5954]), .S0(n27117), .S1(n26642), .ZN(n22225) );
  MUX41 U10216 ( .I0(ram[6106]), .I1(ram[6098]), .I2(ram[6090]), .I3(
        ram[6082]), .S0(n27117), .S1(n26642), .ZN(n22230) );
  MUX41 U10217 ( .I0(ram[5850]), .I1(ram[5842]), .I2(ram[5834]), .I3(
        ram[5826]), .S0(n27116), .S1(n26641), .ZN(n22220) );
  MUX41 U10218 ( .I0(ram[5722]), .I1(ram[5714]), .I2(ram[5706]), .I3(
        ram[5698]), .S0(n27116), .S1(n26641), .ZN(n22215) );
  MUX41 U10219 ( .I0(ram[4442]), .I1(ram[4434]), .I2(ram[4426]), .I3(
        ram[4418]), .S0(n27113), .S1(n26638), .ZN(n22165) );
  MUX41 U10220 ( .I0(ram[4570]), .I1(ram[4562]), .I2(ram[4554]), .I3(
        ram[4546]), .S0(n27113), .S1(n26638), .ZN(n22170) );
  MUX41 U10221 ( .I0(ram[4954]), .I1(ram[4946]), .I2(ram[4938]), .I3(
        ram[4930]), .S0(n27114), .S1(n26639), .ZN(n22185) );
  MUX41 U10222 ( .I0(ram[11610]), .I1(ram[11602]), .I2(ram[11594]), .I3(
        ram[11586]), .S0(n27130), .S1(n26655), .ZN(n22461) );
  MUX41 U10223 ( .I0(ram[11738]), .I1(ram[11730]), .I2(ram[11722]), .I3(
        ram[11714]), .S0(n27130), .S1(n26655), .ZN(n22466) );
  MUX41 U10224 ( .I0(ram[11482]), .I1(ram[11474]), .I2(ram[11466]), .I3(
        ram[11458]), .S0(n27130), .S1(n26655), .ZN(n22456) );
  MUX41 U10225 ( .I0(ram[11354]), .I1(ram[11346]), .I2(ram[11338]), .I3(
        ram[11330]), .S0(n27129), .S1(n26654), .ZN(n22451) );
  MUX41 U10226 ( .I0(ram[12122]), .I1(ram[12114]), .I2(ram[12106]), .I3(
        ram[12098]), .S0(n27131), .S1(n26656), .ZN(n22481) );
  MUX41 U10227 ( .I0(ram[12250]), .I1(ram[12242]), .I2(ram[12234]), .I3(
        ram[12226]), .S0(n27132), .S1(n26657), .ZN(n22486) );
  MUX41 U10228 ( .I0(ram[11994]), .I1(ram[11986]), .I2(ram[11978]), .I3(
        ram[11970]), .S0(n27131), .S1(n26656), .ZN(n22476) );
  MUX41 U10229 ( .I0(ram[11866]), .I1(ram[11858]), .I2(ram[11850]), .I3(
        ram[11842]), .S0(n27131), .S1(n26656), .ZN(n22471) );
  MUX41 U10230 ( .I0(ram[10586]), .I1(ram[10578]), .I2(ram[10570]), .I3(
        ram[10562]), .S0(n27128), .S1(n26653), .ZN(n22421) );
  MUX41 U10231 ( .I0(ram[10714]), .I1(ram[10706]), .I2(ram[10698]), .I3(
        ram[10690]), .S0(n27128), .S1(n26653), .ZN(n22426) );
  MUX41 U10232 ( .I0(ram[10458]), .I1(ram[10450]), .I2(ram[10442]), .I3(
        ram[10434]), .S0(n27127), .S1(n26652), .ZN(n22416) );
  MUX41 U10233 ( .I0(ram[10330]), .I1(ram[10322]), .I2(ram[10314]), .I3(
        ram[10306]), .S0(n27127), .S1(n26652), .ZN(n22411) );
  MUX41 U10234 ( .I0(ram[11098]), .I1(ram[11090]), .I2(ram[11082]), .I3(
        ram[11074]), .S0(n27129), .S1(n26654), .ZN(n22441) );
  MUX41 U10235 ( .I0(ram[11226]), .I1(ram[11218]), .I2(ram[11210]), .I3(
        ram[11202]), .S0(n27129), .S1(n26654), .ZN(n22446) );
  MUX41 U10236 ( .I0(ram[10970]), .I1(ram[10962]), .I2(ram[10954]), .I3(
        ram[10946]), .S0(n27129), .S1(n26654), .ZN(n22436) );
  MUX41 U10237 ( .I0(ram[9562]), .I1(ram[9554]), .I2(ram[9546]), .I3(
        ram[9538]), .S0(n27125), .S1(n26650), .ZN(n22376) );
  MUX41 U10238 ( .I0(ram[9690]), .I1(ram[9682]), .I2(ram[9674]), .I3(
        ram[9666]), .S0(n27125), .S1(n26650), .ZN(n22381) );
  MUX41 U10239 ( .I0(ram[9434]), .I1(ram[9426]), .I2(ram[9418]), .I3(
        ram[9410]), .S0(n27125), .S1(n26650), .ZN(n22371) );
  MUX41 U10240 ( .I0(ram[9306]), .I1(ram[9298]), .I2(ram[9290]), .I3(
        ram[9282]), .S0(n27125), .S1(n26650), .ZN(n22366) );
  MUX41 U10241 ( .I0(ram[10074]), .I1(ram[10066]), .I2(ram[10058]), .I3(
        ram[10050]), .S0(n27126), .S1(n26651), .ZN(n22396) );
  MUX41 U10242 ( .I0(ram[10202]), .I1(ram[10194]), .I2(ram[10186]), .I3(
        ram[10178]), .S0(n27127), .S1(n26652), .ZN(n22401) );
  MUX41 U10243 ( .I0(ram[9946]), .I1(ram[9938]), .I2(ram[9930]), .I3(
        ram[9922]), .S0(n27126), .S1(n26651), .ZN(n22391) );
  MUX41 U10244 ( .I0(ram[9818]), .I1(ram[9810]), .I2(ram[9802]), .I3(
        ram[9794]), .S0(n27126), .S1(n26651), .ZN(n22386) );
  MUX41 U10245 ( .I0(ram[8538]), .I1(ram[8530]), .I2(ram[8522]), .I3(
        ram[8514]), .S0(n27123), .S1(n26648), .ZN(n22336) );
  MUX41 U10246 ( .I0(ram[8666]), .I1(ram[8658]), .I2(ram[8650]), .I3(
        ram[8642]), .S0(n27123), .S1(n26648), .ZN(n22341) );
  MUX41 U10247 ( .I0(ram[8410]), .I1(ram[8402]), .I2(ram[8394]), .I3(
        ram[8386]), .S0(n27122), .S1(n26647), .ZN(n22331) );
  MUX41 U10248 ( .I0(ram[8282]), .I1(ram[8274]), .I2(ram[8266]), .I3(
        ram[8258]), .S0(n27122), .S1(n26647), .ZN(n22326) );
  MUX41 U10249 ( .I0(ram[9050]), .I1(ram[9042]), .I2(ram[9034]), .I3(
        ram[9026]), .S0(n27124), .S1(n26649), .ZN(n22356) );
  MUX41 U10250 ( .I0(ram[9178]), .I1(ram[9170]), .I2(ram[9162]), .I3(
        ram[9154]), .S0(n27124), .S1(n26649), .ZN(n22361) );
  MUX41 U10251 ( .I0(ram[15707]), .I1(ram[15699]), .I2(ram[15691]), .I3(
        ram[15683]), .S0(n27179), .S1(n26704), .ZN(n23316) );
  MUX41 U10252 ( .I0(ram[15835]), .I1(ram[15827]), .I2(ram[15819]), .I3(
        ram[15811]), .S0(n27180), .S1(n26705), .ZN(n23321) );
  MUX41 U10253 ( .I0(ram[15579]), .I1(ram[15571]), .I2(ram[15563]), .I3(
        ram[15555]), .S0(n27179), .S1(n26704), .ZN(n23311) );
  MUX41 U10254 ( .I0(ram[15451]), .I1(ram[15443]), .I2(ram[15435]), .I3(
        ram[15427]), .S0(n27179), .S1(n26704), .ZN(n23306) );
  MUX41 U10255 ( .I0(ram[16219]), .I1(ram[16211]), .I2(ram[16203]), .I3(
        ram[16195]), .S0(n27181), .S1(n26706), .ZN(n23336) );
  MUX41 U10256 ( .I0(ram[16347]), .I1(ram[16339]), .I2(ram[16331]), .I3(
        ram[16323]), .S0(n27181), .S1(n26706), .ZN(n23341) );
  MUX41 U10257 ( .I0(ram[16091]), .I1(ram[16083]), .I2(ram[16075]), .I3(
        ram[16067]), .S0(n27180), .S1(n26705), .ZN(n23331) );
  MUX41 U10258 ( .I0(ram[15963]), .I1(ram[15955]), .I2(ram[15947]), .I3(
        ram[15939]), .S0(n27180), .S1(n26705), .ZN(n23326) );
  MUX41 U10259 ( .I0(ram[15195]), .I1(ram[15187]), .I2(ram[15179]), .I3(
        ram[15171]), .S0(n27178), .S1(n26703), .ZN(n23296) );
  MUX41 U10260 ( .I0(ram[15323]), .I1(ram[15315]), .I2(ram[15307]), .I3(
        ram[15299]), .S0(n27178), .S1(n26703), .ZN(n23301) );
  MUX41 U10261 ( .I0(ram[15067]), .I1(ram[15059]), .I2(ram[15051]), .I3(
        ram[15043]), .S0(n27178), .S1(n26703), .ZN(n23291) );
  MUX41 U10262 ( .I0(ram[14939]), .I1(ram[14931]), .I2(ram[14923]), .I3(
        ram[14915]), .S0(n27177), .S1(n26702), .ZN(n23286) );
  MUX41 U10263 ( .I0(ram[14683]), .I1(ram[14675]), .I2(ram[14667]), .I3(
        ram[14659]), .S0(n27177), .S1(n26702), .ZN(n23276) );
  MUX41 U10264 ( .I0(ram[14811]), .I1(ram[14803]), .I2(ram[14795]), .I3(
        ram[14787]), .S0(n27177), .S1(n26702), .ZN(n23281) );
  MUX41 U10265 ( .I0(ram[14555]), .I1(ram[14547]), .I2(ram[14539]), .I3(
        ram[14531]), .S0(n27177), .S1(n26702), .ZN(n23271) );
  MUX41 U10266 ( .I0(ram[14427]), .I1(ram[14419]), .I2(ram[14411]), .I3(
        ram[14403]), .S0(n27176), .S1(n26701), .ZN(n23266) );
  MUX41 U10267 ( .I0(ram[13659]), .I1(ram[13651]), .I2(ram[13643]), .I3(
        ram[13635]), .S0(n27174), .S1(n26699), .ZN(n23231) );
  MUX41 U10268 ( .I0(ram[13787]), .I1(ram[13779]), .I2(ram[13771]), .I3(
        ram[13763]), .S0(n27175), .S1(n26700), .ZN(n23236) );
  MUX41 U10269 ( .I0(ram[13531]), .I1(ram[13523]), .I2(ram[13515]), .I3(
        ram[13507]), .S0(n27174), .S1(n26699), .ZN(n23226) );
  MUX41 U10270 ( .I0(ram[13403]), .I1(ram[13395]), .I2(ram[13387]), .I3(
        ram[13379]), .S0(n27174), .S1(n26699), .ZN(n23221) );
  MUX41 U10271 ( .I0(ram[14171]), .I1(ram[14163]), .I2(ram[14155]), .I3(
        ram[14147]), .S0(n27176), .S1(n26701), .ZN(n23251) );
  MUX41 U10272 ( .I0(ram[14299]), .I1(ram[14291]), .I2(ram[14283]), .I3(
        ram[14275]), .S0(n27176), .S1(n26701), .ZN(n23256) );
  MUX41 U10273 ( .I0(ram[14043]), .I1(ram[14035]), .I2(ram[14027]), .I3(
        ram[14019]), .S0(n27175), .S1(n26700), .ZN(n23246) );
  MUX41 U10274 ( .I0(ram[13915]), .I1(ram[13907]), .I2(ram[13899]), .I3(
        ram[13891]), .S0(n27175), .S1(n26700), .ZN(n23241) );
  MUX41 U10275 ( .I0(ram[13147]), .I1(ram[13139]), .I2(ram[13131]), .I3(
        ram[13123]), .S0(n27173), .S1(n26698), .ZN(n23211) );
  MUX41 U10276 ( .I0(ram[13275]), .I1(ram[13267]), .I2(ram[13259]), .I3(
        ram[13251]), .S0(n27173), .S1(n26698), .ZN(n23216) );
  MUX41 U10277 ( .I0(ram[13019]), .I1(ram[13011]), .I2(ram[13003]), .I3(
        ram[12995]), .S0(n27173), .S1(n26698), .ZN(n23206) );
  MUX41 U10278 ( .I0(ram[12891]), .I1(ram[12883]), .I2(ram[12875]), .I3(
        ram[12867]), .S0(n27173), .S1(n26698), .ZN(n23201) );
  MUX41 U10279 ( .I0(ram[12635]), .I1(ram[12627]), .I2(ram[12619]), .I3(
        ram[12611]), .S0(n27172), .S1(n26697), .ZN(n23191) );
  MUX41 U10280 ( .I0(ram[12763]), .I1(ram[12755]), .I2(ram[12747]), .I3(
        ram[12739]), .S0(n27172), .S1(n26697), .ZN(n23196) );
  MUX41 U10281 ( .I0(ram[12507]), .I1(ram[12499]), .I2(ram[12491]), .I3(
        ram[12483]), .S0(n27172), .S1(n26697), .ZN(n23186) );
  MUX41 U10282 ( .I0(ram[12379]), .I1(ram[12371]), .I2(ram[12363]), .I3(
        ram[12355]), .S0(n27171), .S1(n26696), .ZN(n23181) );
  MUX41 U10283 ( .I0(n22801), .I1(n22802), .I2(n22803), .I3(n22804), .S0(
        n26225), .S1(n26343), .ZN(n22800) );
  MUX41 U10284 ( .I0(ram[3387]), .I1(ram[3379]), .I2(ram[3371]), .I3(
        ram[3363]), .S0(n27150), .S1(n26675), .ZN(n22802) );
  MUX41 U10285 ( .I0(ram[3355]), .I1(ram[3347]), .I2(ram[3339]), .I3(
        ram[3331]), .S0(n27150), .S1(n26675), .ZN(n22804) );
  MUX41 U10286 ( .I0(ram[3451]), .I1(ram[3443]), .I2(ram[3435]), .I3(
        ram[3427]), .S0(n27150), .S1(n26675), .ZN(n22801) );
  MUX41 U10287 ( .I0(n22821), .I1(n22822), .I2(n22823), .I3(n22824), .S0(
        n26226), .S1(n26344), .ZN(n22820) );
  MUX41 U10288 ( .I0(ram[3899]), .I1(ram[3891]), .I2(ram[3883]), .I3(
        ram[3875]), .S0(n27151), .S1(n26676), .ZN(n22822) );
  MUX41 U10289 ( .I0(ram[3867]), .I1(ram[3859]), .I2(ram[3851]), .I3(
        ram[3843]), .S0(n27151), .S1(n26676), .ZN(n22824) );
  MUX41 U10290 ( .I0(ram[3963]), .I1(ram[3955]), .I2(ram[3947]), .I3(
        ram[3939]), .S0(n27151), .S1(n26676), .ZN(n22821) );
  MUX41 U10291 ( .I0(n22761), .I1(n22762), .I2(n22763), .I3(n22764), .S0(
        n26225), .S1(n26343), .ZN(n22760) );
  MUX41 U10292 ( .I0(ram[2331]), .I1(ram[2323]), .I2(ram[2315]), .I3(
        ram[2307]), .S0(n27147), .S1(n26672), .ZN(n22764) );
  MUX41 U10293 ( .I0(ram[2363]), .I1(ram[2355]), .I2(ram[2347]), .I3(
        ram[2339]), .S0(n27147), .S1(n26672), .ZN(n22762) );
  MUX41 U10294 ( .I0(ram[2427]), .I1(ram[2419]), .I2(ram[2411]), .I3(
        ram[2403]), .S0(n27147), .S1(n26672), .ZN(n22761) );
  MUX41 U10295 ( .I0(n22781), .I1(n22782), .I2(n22783), .I3(n22784), .S0(
        n26225), .S1(n26343), .ZN(n22780) );
  MUX41 U10296 ( .I0(ram[2843]), .I1(ram[2835]), .I2(ram[2827]), .I3(
        ram[2819]), .S0(n27148), .S1(n26673), .ZN(n22784) );
  MUX41 U10297 ( .I0(ram[2875]), .I1(ram[2867]), .I2(ram[2859]), .I3(
        ram[2851]), .S0(n27148), .S1(n26673), .ZN(n22782) );
  MUX41 U10298 ( .I0(ram[2939]), .I1(ram[2931]), .I2(ram[2923]), .I3(
        ram[2915]), .S0(n27149), .S1(n26674), .ZN(n22781) );
  MUX41 U10299 ( .I0(n22716), .I1(n22717), .I2(n22718), .I3(n22719), .S0(
        n26224), .S1(n26342), .ZN(n22715) );
  MUX41 U10300 ( .I0(ram[1339]), .I1(ram[1331]), .I2(ram[1323]), .I3(
        ram[1315]), .S0(n27145), .S1(n26670), .ZN(n22717) );
  MUX41 U10301 ( .I0(ram[1307]), .I1(ram[1299]), .I2(ram[1291]), .I3(
        ram[1283]), .S0(n27145), .S1(n26670), .ZN(n22719) );
  MUX41 U10302 ( .I0(ram[1403]), .I1(ram[1395]), .I2(ram[1387]), .I3(
        ram[1379]), .S0(n27145), .S1(n26670), .ZN(n22716) );
  MUX41 U10303 ( .I0(n22736), .I1(n22737), .I2(n22738), .I3(n22739), .S0(
        n26224), .S1(n26342), .ZN(n22735) );
  MUX41 U10304 ( .I0(ram[1819]), .I1(ram[1811]), .I2(ram[1803]), .I3(
        ram[1795]), .S0(n27146), .S1(n26671), .ZN(n22739) );
  MUX41 U10305 ( .I0(ram[1851]), .I1(ram[1843]), .I2(ram[1835]), .I3(
        ram[1827]), .S0(n27146), .S1(n26671), .ZN(n22737) );
  MUX41 U10306 ( .I0(ram[1915]), .I1(ram[1907]), .I2(ram[1899]), .I3(
        ram[1891]), .S0(n27146), .S1(n26671), .ZN(n22736) );
  MUX41 U10307 ( .I0(n22676), .I1(n22677), .I2(n22678), .I3(n22679), .S0(
        n26223), .S1(n26341), .ZN(n22675) );
  MUX41 U10308 ( .I0(ram[283]), .I1(ram[275]), .I2(ram[267]), .I3(
        ram[259]), .S0(n27142), .S1(n26667), .ZN(n22679) );
  MUX41 U10309 ( .I0(ram[315]), .I1(ram[307]), .I2(ram[299]), .I3(
        ram[291]), .S0(n27142), .S1(n26667), .ZN(n22677) );
  MUX41 U10310 ( .I0(ram[379]), .I1(ram[371]), .I2(ram[363]), .I3(
        ram[355]), .S0(n27142), .S1(n26667), .ZN(n22676) );
  MUX41 U10311 ( .I0(n22696), .I1(n22697), .I2(n22698), .I3(n22699), .S0(
        n26224), .S1(n26342), .ZN(n22695) );
  MUX41 U10312 ( .I0(ram[795]), .I1(ram[787]), .I2(ram[779]), .I3(
        ram[771]), .S0(n27143), .S1(n26668), .ZN(n22699) );
  MUX41 U10313 ( .I0(ram[827]), .I1(ram[819]), .I2(ram[811]), .I3(
        ram[803]), .S0(n27144), .S1(n26669), .ZN(n22697) );
  MUX41 U10314 ( .I0(ram[891]), .I1(ram[883]), .I2(ram[875]), .I3(
        ram[867]), .S0(n27144), .S1(n26669), .ZN(n22696) );
  MUX41 U10315 ( .I0(ram[7515]), .I1(ram[7507]), .I2(ram[7499]), .I3(
        ram[7491]), .S0(n27160), .S1(n26685), .ZN(n22974) );
  MUX41 U10316 ( .I0(ram[7643]), .I1(ram[7635]), .I2(ram[7627]), .I3(
        ram[7619]), .S0(n27160), .S1(n26685), .ZN(n22979) );
  MUX41 U10317 ( .I0(ram[7387]), .I1(ram[7379]), .I2(ram[7371]), .I3(
        ram[7363]), .S0(n27159), .S1(n26684), .ZN(n22969) );
  MUX41 U10318 ( .I0(ram[7259]), .I1(ram[7251]), .I2(ram[7243]), .I3(
        ram[7235]), .S0(n27159), .S1(n26684), .ZN(n22964) );
  MUX41 U10319 ( .I0(ram[8027]), .I1(ram[8019]), .I2(ram[8011]), .I3(
        ram[8003]), .S0(n27161), .S1(n26686), .ZN(n22994) );
  MUX41 U10320 ( .I0(ram[8155]), .I1(ram[8147]), .I2(ram[8139]), .I3(
        ram[8131]), .S0(n27161), .S1(n26686), .ZN(n22999) );
  MUX41 U10321 ( .I0(ram[7899]), .I1(ram[7891]), .I2(ram[7883]), .I3(
        ram[7875]), .S0(n27161), .S1(n26686), .ZN(n22989) );
  MUX41 U10322 ( .I0(ram[7771]), .I1(ram[7763]), .I2(ram[7755]), .I3(
        ram[7747]), .S0(n27160), .S1(n26685), .ZN(n22984) );
  MUX41 U10323 ( .I0(ram[6491]), .I1(ram[6483]), .I2(ram[6475]), .I3(
        ram[6467]), .S0(n27157), .S1(n26682), .ZN(n22934) );
  MUX41 U10324 ( .I0(ram[6619]), .I1(ram[6611]), .I2(ram[6603]), .I3(
        ram[6595]), .S0(n27157), .S1(n26682), .ZN(n22939) );
  MUX41 U10325 ( .I0(ram[6363]), .I1(ram[6355]), .I2(ram[6347]), .I3(
        ram[6339]), .S0(n27157), .S1(n26682), .ZN(n22929) );
  MUX41 U10326 ( .I0(ram[6235]), .I1(ram[6227]), .I2(ram[6219]), .I3(
        ram[6211]), .S0(n27157), .S1(n26682), .ZN(n22924) );
  MUX41 U10327 ( .I0(ram[7003]), .I1(ram[6995]), .I2(ram[6987]), .I3(
        ram[6979]), .S0(n27158), .S1(n26683), .ZN(n22954) );
  MUX41 U10328 ( .I0(ram[7131]), .I1(ram[7123]), .I2(ram[7115]), .I3(
        ram[7107]), .S0(n27159), .S1(n26684), .ZN(n22959) );
  MUX41 U10329 ( .I0(ram[6875]), .I1(ram[6867]), .I2(ram[6859]), .I3(
        ram[6851]), .S0(n27158), .S1(n26683), .ZN(n22949) );
  MUX41 U10330 ( .I0(ram[6747]), .I1(ram[6739]), .I2(ram[6731]), .I3(
        ram[6723]), .S0(n27158), .S1(n26683), .ZN(n22944) );
  MUX41 U10331 ( .I0(ram[5467]), .I1(ram[5459]), .I2(ram[5451]), .I3(
        ram[5443]), .S0(n27155), .S1(n26680), .ZN(n22889) );
  MUX41 U10332 ( .I0(ram[5595]), .I1(ram[5587]), .I2(ram[5579]), .I3(
        ram[5571]), .S0(n27155), .S1(n26680), .ZN(n22894) );
  MUX41 U10333 ( .I0(ram[5339]), .I1(ram[5331]), .I2(ram[5323]), .I3(
        ram[5315]), .S0(n27154), .S1(n26679), .ZN(n22884) );
  MUX41 U10334 ( .I0(ram[5211]), .I1(ram[5203]), .I2(ram[5195]), .I3(
        ram[5187]), .S0(n27154), .S1(n26679), .ZN(n22879) );
  MUX41 U10335 ( .I0(ram[5979]), .I1(ram[5971]), .I2(ram[5963]), .I3(
        ram[5955]), .S0(n27156), .S1(n26681), .ZN(n22909) );
  MUX41 U10336 ( .I0(ram[6107]), .I1(ram[6099]), .I2(ram[6091]), .I3(
        ram[6083]), .S0(n27156), .S1(n26681), .ZN(n22914) );
  MUX41 U10337 ( .I0(ram[5851]), .I1(ram[5843]), .I2(ram[5835]), .I3(
        ram[5827]), .S0(n27156), .S1(n26681), .ZN(n22904) );
  MUX41 U10338 ( .I0(ram[5723]), .I1(ram[5715]), .I2(ram[5707]), .I3(
        ram[5699]), .S0(n27155), .S1(n26680), .ZN(n22899) );
  MUX41 U10339 ( .I0(ram[4443]), .I1(ram[4435]), .I2(ram[4427]), .I3(
        ram[4419]), .S0(n27152), .S1(n26677), .ZN(n22849) );
  MUX41 U10340 ( .I0(ram[4571]), .I1(ram[4563]), .I2(ram[4555]), .I3(
        ram[4547]), .S0(n27153), .S1(n26678), .ZN(n22854) );
  MUX41 U10341 ( .I0(ram[4955]), .I1(ram[4947]), .I2(ram[4939]), .I3(
        ram[4931]), .S0(n27153), .S1(n26678), .ZN(n22869) );
  MUX41 U10342 ( .I0(ram[11611]), .I1(ram[11603]), .I2(ram[11595]), .I3(
        ram[11587]), .S0(n27169), .S1(n26694), .ZN(n23145) );
  MUX41 U10343 ( .I0(ram[11739]), .I1(ram[11731]), .I2(ram[11723]), .I3(
        ram[11715]), .S0(n27170), .S1(n26695), .ZN(n23150) );
  MUX41 U10344 ( .I0(ram[11483]), .I1(ram[11475]), .I2(ram[11467]), .I3(
        ram[11459]), .S0(n27169), .S1(n26694), .ZN(n23140) );
  MUX41 U10345 ( .I0(ram[11355]), .I1(ram[11347]), .I2(ram[11339]), .I3(
        ram[11331]), .S0(n27169), .S1(n26694), .ZN(n23135) );
  MUX41 U10346 ( .I0(ram[12123]), .I1(ram[12115]), .I2(ram[12107]), .I3(
        ram[12099]), .S0(n27171), .S1(n26696), .ZN(n23165) );
  MUX41 U10347 ( .I0(ram[12251]), .I1(ram[12243]), .I2(ram[12235]), .I3(
        ram[12227]), .S0(n27171), .S1(n26696), .ZN(n23170) );
  MUX41 U10348 ( .I0(ram[11995]), .I1(ram[11987]), .I2(ram[11979]), .I3(
        ram[11971]), .S0(n27170), .S1(n26695), .ZN(n23160) );
  MUX41 U10349 ( .I0(ram[11867]), .I1(ram[11859]), .I2(ram[11851]), .I3(
        ram[11843]), .S0(n27170), .S1(n26695), .ZN(n23155) );
  MUX41 U10350 ( .I0(ram[10587]), .I1(ram[10579]), .I2(ram[10571]), .I3(
        ram[10563]), .S0(n27167), .S1(n26692), .ZN(n23105) );
  MUX41 U10351 ( .I0(ram[10715]), .I1(ram[10707]), .I2(ram[10699]), .I3(
        ram[10691]), .S0(n27167), .S1(n26692), .ZN(n23110) );
  MUX41 U10352 ( .I0(ram[10459]), .I1(ram[10451]), .I2(ram[10443]), .I3(
        ram[10435]), .S0(n27167), .S1(n26692), .ZN(n23100) );
  MUX41 U10353 ( .I0(ram[10331]), .I1(ram[10323]), .I2(ram[10315]), .I3(
        ram[10307]), .S0(n27166), .S1(n26691), .ZN(n23095) );
  MUX41 U10354 ( .I0(ram[11099]), .I1(ram[11091]), .I2(ram[11083]), .I3(
        ram[11075]), .S0(n27168), .S1(n26693), .ZN(n23125) );
  MUX41 U10355 ( .I0(ram[11227]), .I1(ram[11219]), .I2(ram[11211]), .I3(
        ram[11203]), .S0(n27169), .S1(n26694), .ZN(n23130) );
  MUX41 U10356 ( .I0(ram[10971]), .I1(ram[10963]), .I2(ram[10955]), .I3(
        ram[10947]), .S0(n27168), .S1(n26693), .ZN(n23120) );
  MUX41 U10357 ( .I0(ram[9563]), .I1(ram[9555]), .I2(ram[9547]), .I3(
        ram[9539]), .S0(n27165), .S1(n26690), .ZN(n23060) );
  MUX41 U10358 ( .I0(ram[9691]), .I1(ram[9683]), .I2(ram[9675]), .I3(
        ram[9667]), .S0(n27165), .S1(n26690), .ZN(n23065) );
  MUX41 U10359 ( .I0(ram[9435]), .I1(ram[9427]), .I2(ram[9419]), .I3(
        ram[9411]), .S0(n27164), .S1(n26689), .ZN(n23055) );
  MUX41 U10360 ( .I0(ram[9307]), .I1(ram[9299]), .I2(ram[9291]), .I3(
        ram[9283]), .S0(n27164), .S1(n26689), .ZN(n23050) );
  MUX41 U10361 ( .I0(ram[10075]), .I1(ram[10067]), .I2(ram[10059]), .I3(
        ram[10051]), .S0(n27166), .S1(n26691), .ZN(n23080) );
  MUX41 U10362 ( .I0(ram[10203]), .I1(ram[10195]), .I2(ram[10187]), .I3(
        ram[10179]), .S0(n27166), .S1(n26691), .ZN(n23085) );
  MUX41 U10363 ( .I0(ram[9947]), .I1(ram[9939]), .I2(ram[9931]), .I3(
        ram[9923]), .S0(n27165), .S1(n26690), .ZN(n23075) );
  MUX41 U10364 ( .I0(ram[9819]), .I1(ram[9811]), .I2(ram[9803]), .I3(
        ram[9795]), .S0(n27165), .S1(n26690), .ZN(n23070) );
  MUX41 U10365 ( .I0(ram[8539]), .I1(ram[8531]), .I2(ram[8523]), .I3(
        ram[8515]), .S0(n27162), .S1(n26687), .ZN(n23020) );
  MUX41 U10366 ( .I0(ram[8667]), .I1(ram[8659]), .I2(ram[8651]), .I3(
        ram[8643]), .S0(n27162), .S1(n26687), .ZN(n23025) );
  MUX41 U10367 ( .I0(ram[8411]), .I1(ram[8403]), .I2(ram[8395]), .I3(
        ram[8387]), .S0(n27162), .S1(n26687), .ZN(n23015) );
  MUX41 U10368 ( .I0(ram[8283]), .I1(ram[8275]), .I2(ram[8267]), .I3(
        ram[8259]), .S0(n27161), .S1(n26686), .ZN(n23010) );
  MUX41 U10369 ( .I0(ram[9051]), .I1(ram[9043]), .I2(ram[9035]), .I3(
        ram[9027]), .S0(n27163), .S1(n26688), .ZN(n23040) );
  MUX41 U10370 ( .I0(ram[9179]), .I1(ram[9171]), .I2(ram[9163]), .I3(
        ram[9155]), .S0(n27164), .S1(n26689), .ZN(n23045) );
  MUX41 U10371 ( .I0(ram[15708]), .I1(ram[15700]), .I2(ram[15692]), .I3(
        ram[15684]), .S0(n27219), .S1(n26744), .ZN(n24000) );
  MUX41 U10372 ( .I0(ram[15836]), .I1(ram[15828]), .I2(ram[15820]), .I3(
        ram[15812]), .S0(n27219), .S1(n26744), .ZN(n24005) );
  MUX41 U10373 ( .I0(ram[15580]), .I1(ram[15572]), .I2(ram[15564]), .I3(
        ram[15556]), .S0(n27218), .S1(n26743), .ZN(n23995) );
  MUX41 U10374 ( .I0(ram[15452]), .I1(ram[15444]), .I2(ram[15436]), .I3(
        ram[15428]), .S0(n27218), .S1(n26743), .ZN(n23990) );
  MUX41 U10375 ( .I0(ram[16220]), .I1(ram[16212]), .I2(ram[16204]), .I3(
        ram[16196]), .S0(n27220), .S1(n26745), .ZN(n24020) );
  MUX41 U10376 ( .I0(ram[16348]), .I1(ram[16340]), .I2(ram[16332]), .I3(
        ram[16324]), .S0(n27220), .S1(n26745), .ZN(n24025) );
  MUX41 U10377 ( .I0(ram[16092]), .I1(ram[16084]), .I2(ram[16076]), .I3(
        ram[16068]), .S0(n27220), .S1(n26745), .ZN(n24015) );
  MUX41 U10378 ( .I0(ram[15964]), .I1(ram[15956]), .I2(ram[15948]), .I3(
        ram[15940]), .S0(n27219), .S1(n26744), .ZN(n24010) );
  MUX41 U10379 ( .I0(ram[15196]), .I1(ram[15188]), .I2(ram[15180]), .I3(
        ram[15172]), .S0(n27217), .S1(n26742), .ZN(n23980) );
  MUX41 U10380 ( .I0(ram[15324]), .I1(ram[15316]), .I2(ram[15308]), .I3(
        ram[15300]), .S0(n27218), .S1(n26743), .ZN(n23985) );
  MUX41 U10381 ( .I0(ram[15068]), .I1(ram[15060]), .I2(ram[15052]), .I3(
        ram[15044]), .S0(n27217), .S1(n26742), .ZN(n23975) );
  MUX41 U10382 ( .I0(ram[14940]), .I1(ram[14932]), .I2(ram[14924]), .I3(
        ram[14916]), .S0(n27217), .S1(n26742), .ZN(n23970) );
  MUX41 U10383 ( .I0(ram[14684]), .I1(ram[14676]), .I2(ram[14668]), .I3(
        ram[14660]), .S0(n27216), .S1(n26741), .ZN(n23960) );
  MUX41 U10384 ( .I0(ram[14812]), .I1(ram[14804]), .I2(ram[14796]), .I3(
        ram[14788]), .S0(n27217), .S1(n26742), .ZN(n23965) );
  MUX41 U10385 ( .I0(ram[14556]), .I1(ram[14548]), .I2(ram[14540]), .I3(
        ram[14532]), .S0(n27216), .S1(n26741), .ZN(n23955) );
  MUX41 U10386 ( .I0(ram[14428]), .I1(ram[14420]), .I2(ram[14412]), .I3(
        ram[14404]), .S0(n27216), .S1(n26741), .ZN(n23950) );
  MUX41 U10387 ( .I0(ram[13660]), .I1(ram[13652]), .I2(ram[13644]), .I3(
        ram[13636]), .S0(n27214), .S1(n26739), .ZN(n23915) );
  MUX41 U10388 ( .I0(ram[13788]), .I1(ram[13780]), .I2(ram[13772]), .I3(
        ram[13764]), .S0(n27214), .S1(n26739), .ZN(n23920) );
  MUX41 U10389 ( .I0(ram[13532]), .I1(ram[13524]), .I2(ram[13516]), .I3(
        ram[13508]), .S0(n27213), .S1(n26738), .ZN(n23910) );
  MUX41 U10390 ( .I0(ram[13404]), .I1(ram[13396]), .I2(ram[13388]), .I3(
        ram[13380]), .S0(n27213), .S1(n26738), .ZN(n23905) );
  MUX41 U10391 ( .I0(ram[14172]), .I1(ram[14164]), .I2(ram[14156]), .I3(
        ram[14148]), .S0(n27215), .S1(n26740), .ZN(n23935) );
  MUX41 U10392 ( .I0(ram[14300]), .I1(ram[14292]), .I2(ram[14284]), .I3(
        ram[14276]), .S0(n27215), .S1(n26740), .ZN(n23940) );
  MUX41 U10393 ( .I0(ram[14044]), .I1(ram[14036]), .I2(ram[14028]), .I3(
        ram[14020]), .S0(n27215), .S1(n26740), .ZN(n23930) );
  MUX41 U10394 ( .I0(ram[13916]), .I1(ram[13908]), .I2(ram[13900]), .I3(
        ram[13892]), .S0(n27214), .S1(n26739), .ZN(n23925) );
  MUX41 U10395 ( .I0(ram[13148]), .I1(ram[13140]), .I2(ram[13132]), .I3(
        ram[13124]), .S0(n27213), .S1(n26738), .ZN(n23895) );
  MUX41 U10396 ( .I0(ram[13276]), .I1(ram[13268]), .I2(ram[13260]), .I3(
        ram[13252]), .S0(n27213), .S1(n26738), .ZN(n23900) );
  MUX41 U10397 ( .I0(ram[13020]), .I1(ram[13012]), .I2(ram[13004]), .I3(
        ram[12996]), .S0(n27212), .S1(n26737), .ZN(n23890) );
  MUX41 U10398 ( .I0(ram[12892]), .I1(ram[12884]), .I2(ram[12876]), .I3(
        ram[12868]), .S0(n27212), .S1(n26737), .ZN(n23885) );
  MUX41 U10399 ( .I0(ram[12636]), .I1(ram[12628]), .I2(ram[12620]), .I3(
        ram[12612]), .S0(n27211), .S1(n26736), .ZN(n23875) );
  MUX41 U10400 ( .I0(ram[12764]), .I1(ram[12756]), .I2(ram[12748]), .I3(
        ram[12740]), .S0(n27212), .S1(n26737), .ZN(n23880) );
  MUX41 U10401 ( .I0(ram[12508]), .I1(ram[12500]), .I2(ram[12492]), .I3(
        ram[12484]), .S0(n27211), .S1(n26736), .ZN(n23870) );
  MUX41 U10402 ( .I0(ram[12380]), .I1(ram[12372]), .I2(ram[12364]), .I3(
        ram[12356]), .S0(n27211), .S1(n26736), .ZN(n23865) );
  MUX41 U10403 ( .I0(n23485), .I1(n23486), .I2(n23487), .I3(n23488), .S0(
        n26235), .S1(n26353), .ZN(n23484) );
  MUX41 U10404 ( .I0(ram[3388]), .I1(ram[3380]), .I2(ram[3372]), .I3(
        ram[3364]), .S0(n27189), .S1(n26714), .ZN(n23486) );
  MUX41 U10405 ( .I0(ram[3356]), .I1(ram[3348]), .I2(ram[3340]), .I3(
        ram[3332]), .S0(n27189), .S1(n26714), .ZN(n23488) );
  MUX41 U10406 ( .I0(ram[3452]), .I1(ram[3444]), .I2(ram[3436]), .I3(
        ram[3428]), .S0(n27189), .S1(n26714), .ZN(n23485) );
  MUX41 U10407 ( .I0(n23505), .I1(n23506), .I2(n23507), .I3(n23508), .S0(
        n26235), .S1(n26353), .ZN(n23504) );
  MUX41 U10408 ( .I0(ram[3900]), .I1(ram[3892]), .I2(ram[3884]), .I3(
        ram[3876]), .S0(n27190), .S1(n26715), .ZN(n23506) );
  MUX41 U10409 ( .I0(ram[3868]), .I1(ram[3860]), .I2(ram[3852]), .I3(
        ram[3844]), .S0(n27190), .S1(n26715), .ZN(n23508) );
  MUX41 U10410 ( .I0(ram[3964]), .I1(ram[3956]), .I2(ram[3948]), .I3(
        ram[3940]), .S0(n27190), .S1(n26715), .ZN(n23505) );
  MUX41 U10411 ( .I0(n23445), .I1(n23446), .I2(n23447), .I3(n23448), .S0(
        n26235), .S1(n26353), .ZN(n23444) );
  MUX41 U10412 ( .I0(ram[2332]), .I1(ram[2324]), .I2(ram[2316]), .I3(
        ram[2308]), .S0(n27187), .S1(n26712), .ZN(n23448) );
  MUX41 U10413 ( .I0(ram[2364]), .I1(ram[2356]), .I2(ram[2348]), .I3(
        ram[2340]), .S0(n27187), .S1(n26712), .ZN(n23446) );
  MUX41 U10414 ( .I0(ram[2428]), .I1(ram[2420]), .I2(ram[2412]), .I3(
        ram[2404]), .S0(n27187), .S1(n26712), .ZN(n23445) );
  MUX41 U10415 ( .I0(n23465), .I1(n23466), .I2(n23467), .I3(n23468), .S0(
        n26235), .S1(n26353), .ZN(n23464) );
  MUX41 U10416 ( .I0(ram[2844]), .I1(ram[2836]), .I2(ram[2828]), .I3(
        ram[2820]), .S0(n27188), .S1(n26713), .ZN(n23468) );
  MUX41 U10417 ( .I0(ram[2876]), .I1(ram[2868]), .I2(ram[2860]), .I3(
        ram[2852]), .S0(n27188), .S1(n26713), .ZN(n23466) );
  MUX41 U10418 ( .I0(ram[2940]), .I1(ram[2932]), .I2(ram[2924]), .I3(
        ram[2916]), .S0(n27188), .S1(n26713), .ZN(n23465) );
  MUX41 U10419 ( .I0(n23400), .I1(n23401), .I2(n23402), .I3(n23403), .S0(
        n26234), .S1(n26352), .ZN(n23399) );
  MUX41 U10420 ( .I0(ram[1340]), .I1(ram[1332]), .I2(ram[1324]), .I3(
        ram[1316]), .S0(n27184), .S1(n26709), .ZN(n23401) );
  MUX41 U10421 ( .I0(ram[1308]), .I1(ram[1300]), .I2(ram[1292]), .I3(
        ram[1284]), .S0(n27184), .S1(n26709), .ZN(n23403) );
  MUX41 U10422 ( .I0(ram[1404]), .I1(ram[1396]), .I2(ram[1388]), .I3(
        ram[1380]), .S0(n27184), .S1(n26709), .ZN(n23400) );
  MUX41 U10423 ( .I0(n23420), .I1(n23421), .I2(n23422), .I3(n23423), .S0(
        n26234), .S1(n26352), .ZN(n23419) );
  MUX41 U10424 ( .I0(ram[1820]), .I1(ram[1812]), .I2(ram[1804]), .I3(
        ram[1796]), .S0(n27185), .S1(n26710), .ZN(n23423) );
  MUX41 U10425 ( .I0(ram[1852]), .I1(ram[1844]), .I2(ram[1836]), .I3(
        ram[1828]), .S0(n27185), .S1(n26710), .ZN(n23421) );
  MUX41 U10426 ( .I0(ram[1916]), .I1(ram[1908]), .I2(ram[1900]), .I3(
        ram[1892]), .S0(n27186), .S1(n26711), .ZN(n23420) );
  MUX41 U10427 ( .I0(n23360), .I1(n23361), .I2(n23362), .I3(n23363), .S0(
        n26233), .S1(n26351), .ZN(n23359) );
  MUX41 U10428 ( .I0(ram[284]), .I1(ram[276]), .I2(ram[268]), .I3(
        ram[260]), .S0(n27182), .S1(n26707), .ZN(n23363) );
  MUX41 U10429 ( .I0(ram[316]), .I1(ram[308]), .I2(ram[300]), .I3(
        ram[292]), .S0(n27182), .S1(n26707), .ZN(n23361) );
  MUX41 U10430 ( .I0(ram[380]), .I1(ram[372]), .I2(ram[364]), .I3(
        ram[356]), .S0(n27182), .S1(n26707), .ZN(n23360) );
  MUX41 U10431 ( .I0(n23380), .I1(n23381), .I2(n23382), .I3(n23383), .S0(
        n26234), .S1(n26352), .ZN(n23379) );
  MUX41 U10432 ( .I0(ram[796]), .I1(ram[788]), .I2(ram[780]), .I3(
        ram[772]), .S0(n27183), .S1(n26708), .ZN(n23383) );
  MUX41 U10433 ( .I0(ram[828]), .I1(ram[820]), .I2(ram[812]), .I3(
        ram[804]), .S0(n27183), .S1(n26708), .ZN(n23381) );
  MUX41 U10434 ( .I0(ram[892]), .I1(ram[884]), .I2(ram[876]), .I3(
        ram[868]), .S0(n27183), .S1(n26708), .ZN(n23380) );
  MUX41 U10435 ( .I0(ram[7516]), .I1(ram[7508]), .I2(ram[7500]), .I3(
        ram[7492]), .S0(n27199), .S1(n26724), .ZN(n23658) );
  MUX41 U10436 ( .I0(ram[7644]), .I1(ram[7636]), .I2(ram[7628]), .I3(
        ram[7620]), .S0(n27199), .S1(n26724), .ZN(n23663) );
  MUX41 U10437 ( .I0(ram[7388]), .I1(ram[7380]), .I2(ram[7372]), .I3(
        ram[7364]), .S0(n27199), .S1(n26724), .ZN(n23653) );
  MUX41 U10438 ( .I0(ram[7260]), .I1(ram[7252]), .I2(ram[7244]), .I3(
        ram[7236]), .S0(n27198), .S1(n26723), .ZN(n23648) );
  MUX41 U10439 ( .I0(ram[8028]), .I1(ram[8020]), .I2(ram[8012]), .I3(
        ram[8004]), .S0(n27200), .S1(n26725), .ZN(n23678) );
  MUX41 U10440 ( .I0(ram[8156]), .I1(ram[8148]), .I2(ram[8140]), .I3(
        ram[8132]), .S0(n27201), .S1(n26726), .ZN(n23683) );
  MUX41 U10441 ( .I0(ram[7900]), .I1(ram[7892]), .I2(ram[7884]), .I3(
        ram[7876]), .S0(n27200), .S1(n26725), .ZN(n23673) );
  MUX41 U10442 ( .I0(ram[7772]), .I1(ram[7764]), .I2(ram[7756]), .I3(
        ram[7748]), .S0(n27200), .S1(n26725), .ZN(n23668) );
  MUX41 U10443 ( .I0(ram[6492]), .I1(ram[6484]), .I2(ram[6476]), .I3(
        ram[6468]), .S0(n27197), .S1(n26722), .ZN(n23618) );
  MUX41 U10444 ( .I0(ram[6620]), .I1(ram[6612]), .I2(ram[6604]), .I3(
        ram[6596]), .S0(n27197), .S1(n26722), .ZN(n23623) );
  MUX41 U10445 ( .I0(ram[6364]), .I1(ram[6356]), .I2(ram[6348]), .I3(
        ram[6340]), .S0(n27196), .S1(n26721), .ZN(n23613) );
  MUX41 U10446 ( .I0(ram[6236]), .I1(ram[6228]), .I2(ram[6220]), .I3(
        ram[6212]), .S0(n27196), .S1(n26721), .ZN(n23608) );
  MUX41 U10447 ( .I0(ram[7004]), .I1(ram[6996]), .I2(ram[6988]), .I3(
        ram[6980]), .S0(n27198), .S1(n26723), .ZN(n23638) );
  MUX41 U10448 ( .I0(ram[7132]), .I1(ram[7124]), .I2(ram[7116]), .I3(
        ram[7108]), .S0(n27198), .S1(n26723), .ZN(n23643) );
  MUX41 U10449 ( .I0(ram[6876]), .I1(ram[6868]), .I2(ram[6860]), .I3(
        ram[6852]), .S0(n27197), .S1(n26722), .ZN(n23633) );
  MUX41 U10450 ( .I0(ram[6748]), .I1(ram[6740]), .I2(ram[6732]), .I3(
        ram[6724]), .S0(n27197), .S1(n26722), .ZN(n23628) );
  MUX41 U10451 ( .I0(ram[5468]), .I1(ram[5460]), .I2(ram[5452]), .I3(
        ram[5444]), .S0(n27194), .S1(n26719), .ZN(n23573) );
  MUX41 U10452 ( .I0(ram[5596]), .I1(ram[5588]), .I2(ram[5580]), .I3(
        ram[5572]), .S0(n27194), .S1(n26719), .ZN(n23578) );
  MUX41 U10453 ( .I0(ram[5340]), .I1(ram[5332]), .I2(ram[5324]), .I3(
        ram[5316]), .S0(n27194), .S1(n26719), .ZN(n23568) );
  MUX41 U10454 ( .I0(ram[5212]), .I1(ram[5204]), .I2(ram[5196]), .I3(
        ram[5188]), .S0(n27193), .S1(n26718), .ZN(n23563) );
  MUX41 U10455 ( .I0(ram[5980]), .I1(ram[5972]), .I2(ram[5964]), .I3(
        ram[5956]), .S0(n27195), .S1(n26720), .ZN(n23593) );
  MUX41 U10456 ( .I0(ram[6108]), .I1(ram[6100]), .I2(ram[6092]), .I3(
        ram[6084]), .S0(n27196), .S1(n26721), .ZN(n23598) );
  MUX41 U10457 ( .I0(ram[5852]), .I1(ram[5844]), .I2(ram[5836]), .I3(
        ram[5828]), .S0(n27195), .S1(n26720), .ZN(n23588) );
  MUX41 U10458 ( .I0(ram[5724]), .I1(ram[5716]), .I2(ram[5708]), .I3(
        ram[5700]), .S0(n27195), .S1(n26720), .ZN(n23583) );
  MUX41 U10459 ( .I0(ram[4444]), .I1(ram[4436]), .I2(ram[4428]), .I3(
        ram[4420]), .S0(n27192), .S1(n26717), .ZN(n23533) );
  MUX41 U10460 ( .I0(ram[4572]), .I1(ram[4564]), .I2(ram[4556]), .I3(
        ram[4548]), .S0(n27192), .S1(n26717), .ZN(n23538) );
  MUX41 U10461 ( .I0(ram[4956]), .I1(ram[4948]), .I2(ram[4940]), .I3(
        ram[4932]), .S0(n27193), .S1(n26718), .ZN(n23553) );
  MUX41 U10462 ( .I0(ram[11612]), .I1(ram[11604]), .I2(ram[11596]), .I3(
        ram[11588]), .S0(n27209), .S1(n26734), .ZN(n23829) );
  MUX41 U10463 ( .I0(ram[11740]), .I1(ram[11732]), .I2(ram[11724]), .I3(
        ram[11716]), .S0(n27209), .S1(n26734), .ZN(n23834) );
  MUX41 U10464 ( .I0(ram[11484]), .I1(ram[11476]), .I2(ram[11468]), .I3(
        ram[11460]), .S0(n27209), .S1(n26734), .ZN(n23824) );
  MUX41 U10465 ( .I0(ram[11356]), .I1(ram[11348]), .I2(ram[11340]), .I3(
        ram[11332]), .S0(n27208), .S1(n26733), .ZN(n23819) );
  MUX41 U10466 ( .I0(ram[12124]), .I1(ram[12116]), .I2(ram[12108]), .I3(
        ram[12100]), .S0(n27210), .S1(n26735), .ZN(n23849) );
  MUX41 U10467 ( .I0(ram[12252]), .I1(ram[12244]), .I2(ram[12236]), .I3(
        ram[12228]), .S0(n27210), .S1(n26735), .ZN(n23854) );
  MUX41 U10468 ( .I0(ram[11996]), .I1(ram[11988]), .I2(ram[11980]), .I3(
        ram[11972]), .S0(n27210), .S1(n26735), .ZN(n23844) );
  MUX41 U10469 ( .I0(ram[11868]), .I1(ram[11860]), .I2(ram[11852]), .I3(
        ram[11844]), .S0(n27209), .S1(n26734), .ZN(n23839) );
  MUX41 U10470 ( .I0(ram[10588]), .I1(ram[10580]), .I2(ram[10572]), .I3(
        ram[10564]), .S0(n27206), .S1(n26731), .ZN(n23789) );
  MUX41 U10471 ( .I0(ram[10716]), .I1(ram[10708]), .I2(ram[10700]), .I3(
        ram[10692]), .S0(n27207), .S1(n26732), .ZN(n23794) );
  MUX41 U10472 ( .I0(ram[10460]), .I1(ram[10452]), .I2(ram[10444]), .I3(
        ram[10436]), .S0(n27206), .S1(n26731), .ZN(n23784) );
  MUX41 U10473 ( .I0(ram[10332]), .I1(ram[10324]), .I2(ram[10316]), .I3(
        ram[10308]), .S0(n27206), .S1(n26731), .ZN(n23779) );
  MUX41 U10474 ( .I0(ram[11100]), .I1(ram[11092]), .I2(ram[11084]), .I3(
        ram[11076]), .S0(n27208), .S1(n26733), .ZN(n23809) );
  MUX41 U10475 ( .I0(ram[11228]), .I1(ram[11220]), .I2(ram[11212]), .I3(
        ram[11204]), .S0(n27208), .S1(n26733), .ZN(n23814) );
  MUX41 U10476 ( .I0(ram[10972]), .I1(ram[10964]), .I2(ram[10956]), .I3(
        ram[10948]), .S0(n27207), .S1(n26732), .ZN(n23804) );
  MUX41 U10477 ( .I0(ram[9564]), .I1(ram[9556]), .I2(ram[9548]), .I3(
        ram[9540]), .S0(n27204), .S1(n26729), .ZN(n23744) );
  MUX41 U10478 ( .I0(ram[9692]), .I1(ram[9684]), .I2(ram[9676]), .I3(
        ram[9668]), .S0(n27204), .S1(n26729), .ZN(n23749) );
  MUX41 U10479 ( .I0(ram[9436]), .I1(ram[9428]), .I2(ram[9420]), .I3(
        ram[9412]), .S0(n27204), .S1(n26729), .ZN(n23739) );
  MUX41 U10480 ( .I0(ram[9308]), .I1(ram[9300]), .I2(ram[9292]), .I3(
        ram[9284]), .S0(n27203), .S1(n26728), .ZN(n23734) );
  MUX41 U10481 ( .I0(ram[10076]), .I1(ram[10068]), .I2(ram[10060]), .I3(
        ram[10052]), .S0(n27205), .S1(n26730), .ZN(n23764) );
  MUX41 U10482 ( .I0(ram[10204]), .I1(ram[10196]), .I2(ram[10188]), .I3(
        ram[10180]), .S0(n27205), .S1(n26730), .ZN(n23769) );
  MUX41 U10483 ( .I0(ram[9948]), .I1(ram[9940]), .I2(ram[9932]), .I3(
        ram[9924]), .S0(n27205), .S1(n26730), .ZN(n23759) );
  MUX41 U10484 ( .I0(ram[9820]), .I1(ram[9812]), .I2(ram[9804]), .I3(
        ram[9796]), .S0(n27205), .S1(n26730), .ZN(n23754) );
  MUX41 U10485 ( .I0(ram[8540]), .I1(ram[8532]), .I2(ram[8524]), .I3(
        ram[8516]), .S0(n27201), .S1(n26726), .ZN(n23704) );
  MUX41 U10486 ( .I0(ram[8668]), .I1(ram[8660]), .I2(ram[8652]), .I3(
        ram[8644]), .S0(n27202), .S1(n26727), .ZN(n23709) );
  MUX41 U10487 ( .I0(ram[8412]), .I1(ram[8404]), .I2(ram[8396]), .I3(
        ram[8388]), .S0(n27201), .S1(n26726), .ZN(n23699) );
  MUX41 U10488 ( .I0(ram[8284]), .I1(ram[8276]), .I2(ram[8268]), .I3(
        ram[8260]), .S0(n27201), .S1(n26726), .ZN(n23694) );
  MUX41 U10489 ( .I0(ram[9052]), .I1(ram[9044]), .I2(ram[9036]), .I3(
        ram[9028]), .S0(n27203), .S1(n26728), .ZN(n23724) );
  MUX41 U10490 ( .I0(ram[9180]), .I1(ram[9172]), .I2(ram[9164]), .I3(
        ram[9156]), .S0(n27203), .S1(n26728), .ZN(n23729) );
  MUX41 U10491 ( .I0(ram[15709]), .I1(ram[15701]), .I2(ram[15693]), .I3(
        ram[15685]), .S0(n27258), .S1(n26783), .ZN(n24684) );
  MUX41 U10492 ( .I0(ram[15837]), .I1(ram[15829]), .I2(ram[15821]), .I3(
        ram[15813]), .S0(n27258), .S1(n26783), .ZN(n24689) );
  MUX41 U10493 ( .I0(ram[15581]), .I1(ram[15573]), .I2(ram[15565]), .I3(
        ram[15557]), .S0(n27258), .S1(n26783), .ZN(n24679) );
  MUX41 U10494 ( .I0(ram[15453]), .I1(ram[15445]), .I2(ram[15437]), .I3(
        ram[15429]), .S0(n27257), .S1(n26782), .ZN(n24674) );
  MUX41 U10495 ( .I0(ram[16221]), .I1(ram[16213]), .I2(ram[16205]), .I3(
        ram[16197]), .S0(n27259), .S1(n26784), .ZN(n24704) );
  MUX41 U10496 ( .I0(ram[16349]), .I1(ram[16341]), .I2(ram[16333]), .I3(
        ram[16325]), .S0(n27260), .S1(n26785), .ZN(n24709) );
  MUX41 U10497 ( .I0(ram[16093]), .I1(ram[16085]), .I2(ram[16077]), .I3(
        ram[16069]), .S0(n27259), .S1(n26784), .ZN(n24699) );
  MUX41 U10498 ( .I0(ram[15965]), .I1(ram[15957]), .I2(ram[15949]), .I3(
        ram[15941]), .S0(n27259), .S1(n26784), .ZN(n24694) );
  MUX41 U10499 ( .I0(ram[15197]), .I1(ram[15189]), .I2(ram[15181]), .I3(
        ram[15173]), .S0(n27257), .S1(n26782), .ZN(n24664) );
  MUX41 U10500 ( .I0(ram[15325]), .I1(ram[15317]), .I2(ram[15309]), .I3(
        ram[15301]), .S0(n27257), .S1(n26782), .ZN(n24669) );
  MUX41 U10501 ( .I0(ram[15069]), .I1(ram[15061]), .I2(ram[15053]), .I3(
        ram[15045]), .S0(n27257), .S1(n26782), .ZN(n24659) );
  MUX41 U10502 ( .I0(ram[14941]), .I1(ram[14933]), .I2(ram[14925]), .I3(
        ram[14917]), .S0(n27256), .S1(n26781), .ZN(n24654) );
  MUX41 U10503 ( .I0(ram[14685]), .I1(ram[14677]), .I2(ram[14669]), .I3(
        ram[14661]), .S0(n27256), .S1(n26781), .ZN(n24644) );
  MUX41 U10504 ( .I0(ram[14813]), .I1(ram[14805]), .I2(ram[14797]), .I3(
        ram[14789]), .S0(n27256), .S1(n26781), .ZN(n24649) );
  MUX41 U10505 ( .I0(ram[14557]), .I1(ram[14549]), .I2(ram[14541]), .I3(
        ram[14533]), .S0(n27255), .S1(n26780), .ZN(n24639) );
  MUX41 U10506 ( .I0(ram[14429]), .I1(ram[14421]), .I2(ram[14413]), .I3(
        ram[14405]), .S0(n27255), .S1(n26780), .ZN(n24634) );
  MUX41 U10507 ( .I0(ram[13661]), .I1(ram[13653]), .I2(ram[13645]), .I3(
        ram[13637]), .S0(n27253), .S1(n26778), .ZN(n24599) );
  MUX41 U10508 ( .I0(ram[13789]), .I1(ram[13781]), .I2(ram[13773]), .I3(
        ram[13765]), .S0(n27253), .S1(n26778), .ZN(n24604) );
  MUX41 U10509 ( .I0(ram[13533]), .I1(ram[13525]), .I2(ram[13517]), .I3(
        ram[13509]), .S0(n27253), .S1(n26778), .ZN(n24594) );
  MUX41 U10510 ( .I0(ram[13405]), .I1(ram[13397]), .I2(ram[13389]), .I3(
        ram[13381]), .S0(n27253), .S1(n26778), .ZN(n24589) );
  MUX41 U10511 ( .I0(ram[14173]), .I1(ram[14165]), .I2(ram[14157]), .I3(
        ram[14149]), .S0(n27254), .S1(n26779), .ZN(n24619) );
  MUX41 U10512 ( .I0(ram[14301]), .I1(ram[14293]), .I2(ram[14285]), .I3(
        ram[14277]), .S0(n27255), .S1(n26780), .ZN(n24624) );
  MUX41 U10513 ( .I0(ram[14045]), .I1(ram[14037]), .I2(ram[14029]), .I3(
        ram[14021]), .S0(n27254), .S1(n26779), .ZN(n24614) );
  MUX41 U10514 ( .I0(ram[13917]), .I1(ram[13909]), .I2(ram[13901]), .I3(
        ram[13893]), .S0(n27254), .S1(n26779), .ZN(n24609) );
  MUX41 U10515 ( .I0(ram[13149]), .I1(ram[13141]), .I2(ram[13133]), .I3(
        ram[13125]), .S0(n27252), .S1(n26777), .ZN(n24579) );
  MUX41 U10516 ( .I0(ram[13277]), .I1(ram[13269]), .I2(ram[13261]), .I3(
        ram[13253]), .S0(n27252), .S1(n26777), .ZN(n24584) );
  MUX41 U10517 ( .I0(ram[13021]), .I1(ram[13013]), .I2(ram[13005]), .I3(
        ram[12997]), .S0(n27252), .S1(n26777), .ZN(n24574) );
  MUX41 U10518 ( .I0(ram[12893]), .I1(ram[12885]), .I2(ram[12877]), .I3(
        ram[12869]), .S0(n27251), .S1(n26776), .ZN(n24569) );
  MUX41 U10519 ( .I0(ram[12637]), .I1(ram[12629]), .I2(ram[12621]), .I3(
        ram[12613]), .S0(n27251), .S1(n26776), .ZN(n24559) );
  MUX41 U10520 ( .I0(ram[12765]), .I1(ram[12757]), .I2(ram[12749]), .I3(
        ram[12741]), .S0(n27251), .S1(n26776), .ZN(n24564) );
  MUX41 U10521 ( .I0(ram[12509]), .I1(ram[12501]), .I2(ram[12493]), .I3(
        ram[12485]), .S0(n27250), .S1(n26775), .ZN(n24554) );
  MUX41 U10522 ( .I0(ram[12381]), .I1(ram[12373]), .I2(ram[12365]), .I3(
        ram[12357]), .S0(n27250), .S1(n26775), .ZN(n24549) );
  MUX41 U10523 ( .I0(n24169), .I1(n24170), .I2(n24171), .I3(n24172), .S0(
        n26245), .S1(n26363), .ZN(n24168) );
  MUX41 U10524 ( .I0(ram[3389]), .I1(ram[3381]), .I2(ram[3373]), .I3(
        ram[3365]), .S0(n27228), .S1(n26753), .ZN(n24170) );
  MUX41 U10525 ( .I0(ram[3357]), .I1(ram[3349]), .I2(ram[3341]), .I3(
        ram[3333]), .S0(n27228), .S1(n26753), .ZN(n24172) );
  MUX41 U10526 ( .I0(ram[3453]), .I1(ram[3445]), .I2(ram[3437]), .I3(
        ram[3429]), .S0(n27229), .S1(n26754), .ZN(n24169) );
  MUX41 U10527 ( .I0(n24189), .I1(n24190), .I2(n24191), .I3(n24192), .S0(
        n26245), .S1(n26363), .ZN(n24188) );
  MUX41 U10528 ( .I0(ram[3901]), .I1(ram[3893]), .I2(ram[3885]), .I3(
        ram[3877]), .S0(n27230), .S1(n26755), .ZN(n24190) );
  MUX41 U10529 ( .I0(ram[3869]), .I1(ram[3861]), .I2(ram[3853]), .I3(
        ram[3845]), .S0(n27230), .S1(n26755), .ZN(n24192) );
  MUX41 U10530 ( .I0(ram[3965]), .I1(ram[3957]), .I2(ram[3949]), .I3(
        ram[3941]), .S0(n27230), .S1(n26755), .ZN(n24189) );
  MUX41 U10531 ( .I0(n24129), .I1(n24130), .I2(n24131), .I3(n24132), .S0(
        n26244), .S1(n26362), .ZN(n24128) );
  MUX41 U10532 ( .I0(ram[2333]), .I1(ram[2325]), .I2(ram[2317]), .I3(
        ram[2309]), .S0(n27226), .S1(n26751), .ZN(n24132) );
  MUX41 U10533 ( .I0(ram[2365]), .I1(ram[2357]), .I2(ram[2349]), .I3(
        ram[2341]), .S0(n27226), .S1(n26751), .ZN(n24130) );
  MUX41 U10534 ( .I0(ram[2429]), .I1(ram[2421]), .I2(ram[2413]), .I3(
        ram[2405]), .S0(n27226), .S1(n26751), .ZN(n24129) );
  MUX41 U10535 ( .I0(n24149), .I1(n24150), .I2(n24151), .I3(n24152), .S0(
        n26245), .S1(n26363), .ZN(n24148) );
  MUX41 U10536 ( .I0(ram[2845]), .I1(ram[2837]), .I2(ram[2829]), .I3(
        ram[2821]), .S0(n27227), .S1(n26752), .ZN(n24152) );
  MUX41 U10537 ( .I0(ram[2877]), .I1(ram[2869]), .I2(ram[2861]), .I3(
        ram[2853]), .S0(n27227), .S1(n26752), .ZN(n24150) );
  MUX41 U10538 ( .I0(ram[2941]), .I1(ram[2933]), .I2(ram[2925]), .I3(
        ram[2917]), .S0(n27227), .S1(n26752), .ZN(n24149) );
  MUX41 U10539 ( .I0(n24084), .I1(n24085), .I2(n24086), .I3(n24087), .S0(
        n26244), .S1(n26362), .ZN(n24083) );
  MUX41 U10540 ( .I0(ram[1341]), .I1(ram[1333]), .I2(ram[1325]), .I3(
        ram[1317]), .S0(n27224), .S1(n26749), .ZN(n24085) );
  MUX41 U10541 ( .I0(ram[1309]), .I1(ram[1301]), .I2(ram[1293]), .I3(
        ram[1285]), .S0(n27223), .S1(n26748), .ZN(n24087) );
  MUX41 U10542 ( .I0(ram[1405]), .I1(ram[1397]), .I2(ram[1389]), .I3(
        ram[1381]), .S0(n27224), .S1(n26749), .ZN(n24084) );
  MUX41 U10543 ( .I0(n24104), .I1(n24105), .I2(n24106), .I3(n24107), .S0(
        n26244), .S1(n26362), .ZN(n24103) );
  MUX41 U10544 ( .I0(ram[1821]), .I1(ram[1813]), .I2(ram[1805]), .I3(
        ram[1797]), .S0(n27225), .S1(n26750), .ZN(n24107) );
  MUX41 U10545 ( .I0(ram[1853]), .I1(ram[1845]), .I2(ram[1837]), .I3(
        ram[1829]), .S0(n27225), .S1(n26750), .ZN(n24105) );
  MUX41 U10546 ( .I0(ram[1917]), .I1(ram[1909]), .I2(ram[1901]), .I3(
        ram[1893]), .S0(n27225), .S1(n26750), .ZN(n24104) );
  MUX41 U10547 ( .I0(n24044), .I1(n24045), .I2(n24046), .I3(n24047), .S0(
        n26243), .S1(n26361), .ZN(n24043) );
  MUX41 U10548 ( .I0(ram[285]), .I1(ram[277]), .I2(ram[269]), .I3(
        ram[261]), .S0(n27221), .S1(n26746), .ZN(n24047) );
  MUX41 U10549 ( .I0(ram[317]), .I1(ram[309]), .I2(ram[301]), .I3(
        ram[293]), .S0(n27221), .S1(n26746), .ZN(n24045) );
  MUX41 U10550 ( .I0(ram[381]), .I1(ram[373]), .I2(ram[365]), .I3(
        ram[357]), .S0(n27221), .S1(n26746), .ZN(n24044) );
  MUX41 U10551 ( .I0(n24064), .I1(n24065), .I2(n24066), .I3(n24067), .S0(
        n26243), .S1(n26361), .ZN(n24063) );
  MUX41 U10552 ( .I0(ram[797]), .I1(ram[789]), .I2(ram[781]), .I3(
        ram[773]), .S0(n27222), .S1(n26747), .ZN(n24067) );
  MUX41 U10553 ( .I0(ram[829]), .I1(ram[821]), .I2(ram[813]), .I3(
        ram[805]), .S0(n27222), .S1(n26747), .ZN(n24065) );
  MUX41 U10554 ( .I0(ram[893]), .I1(ram[885]), .I2(ram[877]), .I3(
        ram[869]), .S0(n27222), .S1(n26747), .ZN(n24064) );
  MUX41 U10555 ( .I0(ram[7517]), .I1(ram[7509]), .I2(ram[7501]), .I3(
        ram[7493]), .S0(n27238), .S1(n26763), .ZN(n24342) );
  MUX41 U10556 ( .I0(ram[7645]), .I1(ram[7637]), .I2(ram[7629]), .I3(
        ram[7621]), .S0(n27239), .S1(n26764), .ZN(n24347) );
  MUX41 U10557 ( .I0(ram[7389]), .I1(ram[7381]), .I2(ram[7373]), .I3(
        ram[7365]), .S0(n27238), .S1(n26763), .ZN(n24337) );
  MUX41 U10558 ( .I0(ram[7261]), .I1(ram[7253]), .I2(ram[7245]), .I3(
        ram[7237]), .S0(n27238), .S1(n26763), .ZN(n24332) );
  MUX41 U10559 ( .I0(ram[8029]), .I1(ram[8021]), .I2(ram[8013]), .I3(
        ram[8005]), .S0(n27240), .S1(n26765), .ZN(n24362) );
  MUX41 U10560 ( .I0(ram[8157]), .I1(ram[8149]), .I2(ram[8141]), .I3(
        ram[8133]), .S0(n27240), .S1(n26765), .ZN(n24367) );
  MUX41 U10561 ( .I0(ram[7901]), .I1(ram[7893]), .I2(ram[7885]), .I3(
        ram[7877]), .S0(n27239), .S1(n26764), .ZN(n24357) );
  MUX41 U10562 ( .I0(ram[7773]), .I1(ram[7765]), .I2(ram[7757]), .I3(
        ram[7749]), .S0(n27239), .S1(n26764), .ZN(n24352) );
  MUX41 U10563 ( .I0(ram[6493]), .I1(ram[6485]), .I2(ram[6477]), .I3(
        ram[6469]), .S0(n27236), .S1(n26761), .ZN(n24302) );
  MUX41 U10564 ( .I0(ram[6621]), .I1(ram[6613]), .I2(ram[6605]), .I3(
        ram[6597]), .S0(n27236), .S1(n26761), .ZN(n24307) );
  MUX41 U10565 ( .I0(ram[6365]), .I1(ram[6357]), .I2(ram[6349]), .I3(
        ram[6341]), .S0(n27236), .S1(n26761), .ZN(n24297) );
  MUX41 U10566 ( .I0(ram[6237]), .I1(ram[6229]), .I2(ram[6221]), .I3(
        ram[6213]), .S0(n27235), .S1(n26760), .ZN(n24292) );
  MUX41 U10567 ( .I0(ram[7005]), .I1(ram[6997]), .I2(ram[6989]), .I3(
        ram[6981]), .S0(n27237), .S1(n26762), .ZN(n24322) );
  MUX41 U10568 ( .I0(ram[7133]), .I1(ram[7125]), .I2(ram[7117]), .I3(
        ram[7109]), .S0(n27237), .S1(n26762), .ZN(n24327) );
  MUX41 U10569 ( .I0(ram[6877]), .I1(ram[6869]), .I2(ram[6861]), .I3(
        ram[6853]), .S0(n27237), .S1(n26762), .ZN(n24317) );
  MUX41 U10570 ( .I0(ram[6749]), .I1(ram[6741]), .I2(ram[6733]), .I3(
        ram[6725]), .S0(n27237), .S1(n26762), .ZN(n24312) );
  MUX41 U10571 ( .I0(ram[5469]), .I1(ram[5461]), .I2(ram[5453]), .I3(
        ram[5445]), .S0(n27233), .S1(n26758), .ZN(n24257) );
  MUX41 U10572 ( .I0(ram[5597]), .I1(ram[5589]), .I2(ram[5581]), .I3(
        ram[5573]), .S0(n27234), .S1(n26759), .ZN(n24262) );
  MUX41 U10573 ( .I0(ram[5341]), .I1(ram[5333]), .I2(ram[5325]), .I3(
        ram[5317]), .S0(n27233), .S1(n26758), .ZN(n24252) );
  MUX41 U10574 ( .I0(ram[5213]), .I1(ram[5205]), .I2(ram[5197]), .I3(
        ram[5189]), .S0(n27233), .S1(n26758), .ZN(n24247) );
  MUX41 U10575 ( .I0(ram[5981]), .I1(ram[5973]), .I2(ram[5965]), .I3(
        ram[5957]), .S0(n27235), .S1(n26760), .ZN(n24277) );
  MUX41 U10576 ( .I0(ram[6109]), .I1(ram[6101]), .I2(ram[6093]), .I3(
        ram[6085]), .S0(n27235), .S1(n26760), .ZN(n24282) );
  MUX41 U10577 ( .I0(ram[5853]), .I1(ram[5845]), .I2(ram[5837]), .I3(
        ram[5829]), .S0(n27234), .S1(n26759), .ZN(n24272) );
  MUX41 U10578 ( .I0(ram[5725]), .I1(ram[5717]), .I2(ram[5709]), .I3(
        ram[5701]), .S0(n27234), .S1(n26759), .ZN(n24267) );
  MUX41 U10579 ( .I0(ram[4445]), .I1(ram[4437]), .I2(ram[4429]), .I3(
        ram[4421]), .S0(n27231), .S1(n26756), .ZN(n24217) );
  MUX41 U10580 ( .I0(ram[4573]), .I1(ram[4565]), .I2(ram[4557]), .I3(
        ram[4549]), .S0(n27231), .S1(n26756), .ZN(n24222) );
  MUX41 U10581 ( .I0(ram[4957]), .I1(ram[4949]), .I2(ram[4941]), .I3(
        ram[4933]), .S0(n27232), .S1(n26757), .ZN(n24237) );
  MUX41 U10582 ( .I0(ram[11613]), .I1(ram[11605]), .I2(ram[11597]), .I3(
        ram[11589]), .S0(n27248), .S1(n26773), .ZN(n24513) );
  MUX41 U10583 ( .I0(ram[11741]), .I1(ram[11733]), .I2(ram[11725]), .I3(
        ram[11717]), .S0(n27249), .S1(n26774), .ZN(n24518) );
  MUX41 U10584 ( .I0(ram[11485]), .I1(ram[11477]), .I2(ram[11469]), .I3(
        ram[11461]), .S0(n27248), .S1(n26773), .ZN(n24508) );
  MUX41 U10585 ( .I0(ram[11357]), .I1(ram[11349]), .I2(ram[11341]), .I3(
        ram[11333]), .S0(n27248), .S1(n26773), .ZN(n24503) );
  MUX41 U10586 ( .I0(ram[12125]), .I1(ram[12117]), .I2(ram[12109]), .I3(
        ram[12101]), .S0(n27249), .S1(n26774), .ZN(n24533) );
  MUX41 U10587 ( .I0(ram[12253]), .I1(ram[12245]), .I2(ram[12237]), .I3(
        ram[12229]), .S0(n27250), .S1(n26775), .ZN(n24538) );
  MUX41 U10588 ( .I0(ram[11997]), .I1(ram[11989]), .I2(ram[11981]), .I3(
        ram[11973]), .S0(n27249), .S1(n26774), .ZN(n24528) );
  MUX41 U10589 ( .I0(ram[11869]), .I1(ram[11861]), .I2(ram[11853]), .I3(
        ram[11845]), .S0(n27249), .S1(n26774), .ZN(n24523) );
  MUX41 U10590 ( .I0(ram[10589]), .I1(ram[10581]), .I2(ram[10573]), .I3(
        ram[10565]), .S0(n27246), .S1(n26771), .ZN(n24473) );
  MUX41 U10591 ( .I0(ram[10717]), .I1(ram[10709]), .I2(ram[10701]), .I3(
        ram[10693]), .S0(n27246), .S1(n26771), .ZN(n24478) );
  MUX41 U10592 ( .I0(ram[10461]), .I1(ram[10453]), .I2(ram[10445]), .I3(
        ram[10437]), .S0(n27245), .S1(n26770), .ZN(n24468) );
  MUX41 U10593 ( .I0(ram[10333]), .I1(ram[10325]), .I2(ram[10317]), .I3(
        ram[10309]), .S0(n27245), .S1(n26770), .ZN(n24463) );
  MUX41 U10594 ( .I0(ram[11101]), .I1(ram[11093]), .I2(ram[11085]), .I3(
        ram[11077]), .S0(n27247), .S1(n26772), .ZN(n24493) );
  MUX41 U10595 ( .I0(ram[11229]), .I1(ram[11221]), .I2(ram[11213]), .I3(
        ram[11205]), .S0(n27247), .S1(n26772), .ZN(n24498) );
  MUX41 U10596 ( .I0(ram[10973]), .I1(ram[10965]), .I2(ram[10957]), .I3(
        ram[10949]), .S0(n27247), .S1(n26772), .ZN(n24488) );
  MUX41 U10597 ( .I0(ram[9565]), .I1(ram[9557]), .I2(ram[9549]), .I3(
        ram[9541]), .S0(n27243), .S1(n26768), .ZN(n24428) );
  MUX41 U10598 ( .I0(ram[9693]), .I1(ram[9685]), .I2(ram[9677]), .I3(
        ram[9669]), .S0(n27244), .S1(n26769), .ZN(n24433) );
  MUX41 U10599 ( .I0(ram[9437]), .I1(ram[9429]), .I2(ram[9421]), .I3(
        ram[9413]), .S0(n27243), .S1(n26768), .ZN(n24423) );
  MUX41 U10600 ( .I0(ram[9309]), .I1(ram[9301]), .I2(ram[9293]), .I3(
        ram[9285]), .S0(n27243), .S1(n26768), .ZN(n24418) );
  MUX41 U10601 ( .I0(ram[10077]), .I1(ram[10069]), .I2(ram[10061]), .I3(
        ram[10053]), .S0(n27245), .S1(n26770), .ZN(n24448) );
  MUX41 U10602 ( .I0(ram[10205]), .I1(ram[10197]), .I2(ram[10189]), .I3(
        ram[10181]), .S0(n27245), .S1(n26770), .ZN(n24453) );
  MUX41 U10603 ( .I0(ram[9949]), .I1(ram[9941]), .I2(ram[9933]), .I3(
        ram[9925]), .S0(n27244), .S1(n26769), .ZN(n24443) );
  MUX41 U10604 ( .I0(ram[9821]), .I1(ram[9813]), .I2(ram[9805]), .I3(
        ram[9797]), .S0(n27244), .S1(n26769), .ZN(n24438) );
  MUX41 U10605 ( .I0(ram[8541]), .I1(ram[8533]), .I2(ram[8525]), .I3(
        ram[8517]), .S0(n27241), .S1(n26766), .ZN(n24388) );
  MUX41 U10606 ( .I0(ram[8669]), .I1(ram[8661]), .I2(ram[8653]), .I3(
        ram[8645]), .S0(n27241), .S1(n26766), .ZN(n24393) );
  MUX41 U10607 ( .I0(ram[8413]), .I1(ram[8405]), .I2(ram[8397]), .I3(
        ram[8389]), .S0(n27241), .S1(n26766), .ZN(n24383) );
  MUX41 U10608 ( .I0(ram[8285]), .I1(ram[8277]), .I2(ram[8269]), .I3(
        ram[8261]), .S0(n27240), .S1(n26765), .ZN(n24378) );
  MUX41 U10609 ( .I0(ram[9053]), .I1(ram[9045]), .I2(ram[9037]), .I3(
        ram[9029]), .S0(n27242), .S1(n26767), .ZN(n24408) );
  MUX41 U10610 ( .I0(ram[9181]), .I1(ram[9173]), .I2(ram[9165]), .I3(
        ram[9157]), .S0(n27242), .S1(n26767), .ZN(n24413) );
  MUX41 U10611 ( .I0(ram[15710]), .I1(ram[15702]), .I2(ram[15694]), .I3(
        ram[15686]), .S0(n27297), .S1(n26822), .ZN(n25368) );
  MUX41 U10612 ( .I0(ram[15838]), .I1(ram[15830]), .I2(ram[15822]), .I3(
        ram[15814]), .S0(n27298), .S1(n26823), .ZN(n25373) );
  MUX41 U10613 ( .I0(ram[15582]), .I1(ram[15574]), .I2(ram[15566]), .I3(
        ram[15558]), .S0(n27297), .S1(n26822), .ZN(n25363) );
  MUX41 U10614 ( .I0(ram[15454]), .I1(ram[15446]), .I2(ram[15438]), .I3(
        ram[15430]), .S0(n27297), .S1(n26822), .ZN(n25358) );
  MUX41 U10615 ( .I0(ram[16222]), .I1(ram[16214]), .I2(ram[16206]), .I3(
        ram[16198]), .S0(n27299), .S1(n26824), .ZN(n25388) );
  MUX41 U10616 ( .I0(ram[16350]), .I1(ram[16342]), .I2(ram[16334]), .I3(
        ram[16326]), .S0(n27299), .S1(n26824), .ZN(n25393) );
  MUX41 U10617 ( .I0(ram[16094]), .I1(ram[16086]), .I2(ram[16078]), .I3(
        ram[16070]), .S0(n27298), .S1(n26823), .ZN(n25383) );
  MUX41 U10618 ( .I0(ram[15966]), .I1(ram[15958]), .I2(ram[15950]), .I3(
        ram[15942]), .S0(n27298), .S1(n26823), .ZN(n25378) );
  MUX41 U10619 ( .I0(ram[15198]), .I1(ram[15190]), .I2(ram[15182]), .I3(
        ram[15174]), .S0(n27296), .S1(n26821), .ZN(n25348) );
  MUX41 U10620 ( .I0(ram[15326]), .I1(ram[15318]), .I2(ram[15310]), .I3(
        ram[15302]), .S0(n27297), .S1(n26822), .ZN(n25353) );
  MUX41 U10621 ( .I0(ram[15070]), .I1(ram[15062]), .I2(ram[15054]), .I3(
        ram[15046]), .S0(n27296), .S1(n26821), .ZN(n25343) );
  MUX41 U10622 ( .I0(ram[14942]), .I1(ram[14934]), .I2(ram[14926]), .I3(
        ram[14918]), .S0(n27296), .S1(n26821), .ZN(n25338) );
  MUX41 U10623 ( .I0(ram[14686]), .I1(ram[14678]), .I2(ram[14670]), .I3(
        ram[14662]), .S0(n27295), .S1(n26820), .ZN(n25328) );
  MUX41 U10624 ( .I0(ram[14814]), .I1(ram[14806]), .I2(ram[14798]), .I3(
        ram[14790]), .S0(n27295), .S1(n26820), .ZN(n25333) );
  MUX41 U10625 ( .I0(ram[14558]), .I1(ram[14550]), .I2(ram[14542]), .I3(
        ram[14534]), .S0(n27295), .S1(n26820), .ZN(n25323) );
  MUX41 U10626 ( .I0(ram[14430]), .I1(ram[14422]), .I2(ram[14414]), .I3(
        ram[14406]), .S0(n27294), .S1(n26819), .ZN(n25318) );
  MUX41 U10627 ( .I0(ram[13662]), .I1(ram[13654]), .I2(ram[13646]), .I3(
        ram[13638]), .S0(n27293), .S1(n26818), .ZN(n25283) );
  MUX41 U10628 ( .I0(ram[13790]), .I1(ram[13782]), .I2(ram[13774]), .I3(
        ram[13766]), .S0(n27293), .S1(n26818), .ZN(n25288) );
  MUX41 U10629 ( .I0(ram[13534]), .I1(ram[13526]), .I2(ram[13518]), .I3(
        ram[13510]), .S0(n27292), .S1(n26817), .ZN(n25278) );
  MUX41 U10630 ( .I0(ram[13406]), .I1(ram[13398]), .I2(ram[13390]), .I3(
        ram[13382]), .S0(n27292), .S1(n26817), .ZN(n25273) );
  MUX41 U10631 ( .I0(ram[14174]), .I1(ram[14166]), .I2(ram[14158]), .I3(
        ram[14150]), .S0(n27294), .S1(n26819), .ZN(n25303) );
  MUX41 U10632 ( .I0(ram[14302]), .I1(ram[14294]), .I2(ram[14286]), .I3(
        ram[14278]), .S0(n27294), .S1(n26819), .ZN(n25308) );
  MUX41 U10633 ( .I0(ram[14046]), .I1(ram[14038]), .I2(ram[14030]), .I3(
        ram[14022]), .S0(n27293), .S1(n26818), .ZN(n25298) );
  MUX41 U10634 ( .I0(ram[13918]), .I1(ram[13910]), .I2(ram[13902]), .I3(
        ram[13894]), .S0(n27293), .S1(n26818), .ZN(n25293) );
  MUX41 U10635 ( .I0(ram[13150]), .I1(ram[13142]), .I2(ram[13134]), .I3(
        ram[13126]), .S0(n27291), .S1(n26816), .ZN(n25263) );
  MUX41 U10636 ( .I0(ram[13278]), .I1(ram[13270]), .I2(ram[13262]), .I3(
        ram[13254]), .S0(n27292), .S1(n26817), .ZN(n25268) );
  MUX41 U10637 ( .I0(ram[13022]), .I1(ram[13014]), .I2(ram[13006]), .I3(
        ram[12998]), .S0(n27291), .S1(n26816), .ZN(n25258) );
  MUX41 U10638 ( .I0(ram[12894]), .I1(ram[12886]), .I2(ram[12878]), .I3(
        ram[12870]), .S0(n27291), .S1(n26816), .ZN(n25253) );
  MUX41 U10639 ( .I0(ram[12638]), .I1(ram[12630]), .I2(ram[12622]), .I3(
        ram[12614]), .S0(n27290), .S1(n26815), .ZN(n25243) );
  MUX41 U10640 ( .I0(ram[12766]), .I1(ram[12758]), .I2(ram[12750]), .I3(
        ram[12742]), .S0(n27290), .S1(n26815), .ZN(n25248) );
  MUX41 U10641 ( .I0(ram[12510]), .I1(ram[12502]), .I2(ram[12494]), .I3(
        ram[12486]), .S0(n27290), .S1(n26815), .ZN(n25238) );
  MUX41 U10642 ( .I0(ram[12382]), .I1(ram[12374]), .I2(ram[12366]), .I3(
        ram[12358]), .S0(n27289), .S1(n26814), .ZN(n25233) );
  MUX41 U10643 ( .I0(n24853), .I1(n24854), .I2(n24855), .I3(n24856), .S0(
        n26255), .S1(n26373), .ZN(n24852) );
  MUX41 U10644 ( .I0(ram[3390]), .I1(ram[3382]), .I2(ram[3374]), .I3(
        ram[3366]), .S0(n27268), .S1(n26793), .ZN(n24854) );
  MUX41 U10645 ( .I0(ram[3358]), .I1(ram[3350]), .I2(ram[3342]), .I3(
        ram[3334]), .S0(n27268), .S1(n26793), .ZN(n24856) );
  MUX41 U10646 ( .I0(ram[3454]), .I1(ram[3446]), .I2(ram[3438]), .I3(
        ram[3430]), .S0(n27268), .S1(n26793), .ZN(n24853) );
  MUX41 U10647 ( .I0(n24873), .I1(n24874), .I2(n24875), .I3(n24876), .S0(
        n26255), .S1(n26373), .ZN(n24872) );
  MUX41 U10648 ( .I0(ram[3902]), .I1(ram[3894]), .I2(ram[3886]), .I3(
        ram[3878]), .S0(n27269), .S1(n26794), .ZN(n24874) );
  MUX41 U10649 ( .I0(ram[3870]), .I1(ram[3862]), .I2(ram[3854]), .I3(
        ram[3846]), .S0(n27269), .S1(n26794), .ZN(n24876) );
  MUX41 U10650 ( .I0(ram[3966]), .I1(ram[3958]), .I2(ram[3950]), .I3(
        ram[3942]), .S0(n27269), .S1(n26794), .ZN(n24873) );
  MUX41 U10651 ( .I0(n24813), .I1(n24814), .I2(n24815), .I3(n24816), .S0(
        n26254), .S1(n26372), .ZN(n24812) );
  MUX41 U10652 ( .I0(ram[2334]), .I1(ram[2326]), .I2(ram[2318]), .I3(
        ram[2310]), .S0(n27265), .S1(n26790), .ZN(n24816) );
  MUX41 U10653 ( .I0(ram[2366]), .I1(ram[2358]), .I2(ram[2350]), .I3(
        ram[2342]), .S0(n27265), .S1(n26790), .ZN(n24814) );
  MUX41 U10654 ( .I0(ram[2430]), .I1(ram[2422]), .I2(ram[2414]), .I3(
        ram[2406]), .S0(n27266), .S1(n26791), .ZN(n24813) );
  MUX41 U10655 ( .I0(n24833), .I1(n24834), .I2(n24835), .I3(n24836), .S0(
        n26255), .S1(n26373), .ZN(n24832) );
  MUX41 U10656 ( .I0(ram[2846]), .I1(ram[2838]), .I2(ram[2830]), .I3(
        ram[2822]), .S0(n27267), .S1(n26792), .ZN(n24836) );
  MUX41 U10657 ( .I0(ram[2878]), .I1(ram[2870]), .I2(ram[2862]), .I3(
        ram[2854]), .S0(n27267), .S1(n26792), .ZN(n24834) );
  MUX41 U10658 ( .I0(ram[2942]), .I1(ram[2934]), .I2(ram[2926]), .I3(
        ram[2918]), .S0(n27267), .S1(n26792), .ZN(n24833) );
  MUX41 U10659 ( .I0(n24768), .I1(n24769), .I2(n24770), .I3(n24771), .S0(
        n26254), .S1(n26372), .ZN(n24767) );
  MUX41 U10660 ( .I0(ram[1342]), .I1(ram[1334]), .I2(ram[1326]), .I3(
        ram[1318]), .S0(n27263), .S1(n26788), .ZN(n24769) );
  MUX41 U10661 ( .I0(ram[1310]), .I1(ram[1302]), .I2(ram[1294]), .I3(
        ram[1286]), .S0(n27263), .S1(n26788), .ZN(n24771) );
  MUX41 U10662 ( .I0(ram[1406]), .I1(ram[1398]), .I2(ram[1390]), .I3(
        ram[1382]), .S0(n27263), .S1(n26788), .ZN(n24768) );
  MUX41 U10663 ( .I0(n24788), .I1(n24789), .I2(n24790), .I3(n24791), .S0(
        n26254), .S1(n26372), .ZN(n24787) );
  MUX41 U10664 ( .I0(ram[1822]), .I1(ram[1814]), .I2(ram[1806]), .I3(
        ram[1798]), .S0(n27264), .S1(n26789), .ZN(n24791) );
  MUX41 U10665 ( .I0(ram[1854]), .I1(ram[1846]), .I2(ram[1838]), .I3(
        ram[1830]), .S0(n27264), .S1(n26789), .ZN(n24789) );
  MUX41 U10666 ( .I0(ram[1918]), .I1(ram[1910]), .I2(ram[1902]), .I3(
        ram[1894]), .S0(n27264), .S1(n26789), .ZN(n24788) );
  MUX41 U10667 ( .I0(n24728), .I1(n24729), .I2(n24730), .I3(n24731), .S0(
        n26253), .S1(n26371), .ZN(n24727) );
  MUX41 U10668 ( .I0(ram[286]), .I1(ram[278]), .I2(ram[270]), .I3(
        ram[262]), .S0(n27260), .S1(n26785), .ZN(n24731) );
  MUX41 U10669 ( .I0(ram[318]), .I1(ram[310]), .I2(ram[302]), .I3(
        ram[294]), .S0(n27260), .S1(n26785), .ZN(n24729) );
  MUX41 U10670 ( .I0(ram[382]), .I1(ram[374]), .I2(ram[366]), .I3(
        ram[358]), .S0(n27261), .S1(n26786), .ZN(n24728) );
  MUX41 U10671 ( .I0(n24748), .I1(n24749), .I2(n24750), .I3(n24751), .S0(
        n26253), .S1(n26371), .ZN(n24747) );
  MUX41 U10672 ( .I0(ram[798]), .I1(ram[790]), .I2(ram[782]), .I3(
        ram[774]), .S0(n27262), .S1(n26787), .ZN(n24751) );
  MUX41 U10673 ( .I0(ram[830]), .I1(ram[822]), .I2(ram[814]), .I3(
        ram[806]), .S0(n27262), .S1(n26787), .ZN(n24749) );
  MUX41 U10674 ( .I0(ram[894]), .I1(ram[886]), .I2(ram[878]), .I3(
        ram[870]), .S0(n27262), .S1(n26787), .ZN(n24748) );
  MUX41 U10675 ( .I0(ram[7518]), .I1(ram[7510]), .I2(ram[7502]), .I3(
        ram[7494]), .S0(n27278), .S1(n26803), .ZN(n25026) );
  MUX41 U10676 ( .I0(ram[7646]), .I1(ram[7638]), .I2(ram[7630]), .I3(
        ram[7622]), .S0(n27278), .S1(n26803), .ZN(n25031) );
  MUX41 U10677 ( .I0(ram[7390]), .I1(ram[7382]), .I2(ram[7374]), .I3(
        ram[7366]), .S0(n27277), .S1(n26802), .ZN(n25021) );
  MUX41 U10678 ( .I0(ram[7262]), .I1(ram[7254]), .I2(ram[7246]), .I3(
        ram[7238]), .S0(n27277), .S1(n26802), .ZN(n25016) );
  MUX41 U10679 ( .I0(ram[8030]), .I1(ram[8022]), .I2(ram[8014]), .I3(
        ram[8006]), .S0(n27279), .S1(n26804), .ZN(n25046) );
  MUX41 U10680 ( .I0(ram[8158]), .I1(ram[8150]), .I2(ram[8142]), .I3(
        ram[8134]), .S0(n27279), .S1(n26804), .ZN(n25051) );
  MUX41 U10681 ( .I0(ram[7902]), .I1(ram[7894]), .I2(ram[7886]), .I3(
        ram[7878]), .S0(n27279), .S1(n26804), .ZN(n25041) );
  MUX41 U10682 ( .I0(ram[7774]), .I1(ram[7766]), .I2(ram[7758]), .I3(
        ram[7750]), .S0(n27278), .S1(n26803), .ZN(n25036) );
  MUX41 U10683 ( .I0(ram[6494]), .I1(ram[6486]), .I2(ram[6478]), .I3(
        ram[6470]), .S0(n27275), .S1(n26800), .ZN(n24986) );
  MUX41 U10684 ( .I0(ram[6622]), .I1(ram[6614]), .I2(ram[6606]), .I3(
        ram[6598]), .S0(n27276), .S1(n26801), .ZN(n24991) );
  MUX41 U10685 ( .I0(ram[6366]), .I1(ram[6358]), .I2(ram[6350]), .I3(
        ram[6342]), .S0(n27275), .S1(n26800), .ZN(n24981) );
  MUX41 U10686 ( .I0(ram[6238]), .I1(ram[6230]), .I2(ram[6222]), .I3(
        ram[6214]), .S0(n27275), .S1(n26800), .ZN(n24976) );
  MUX41 U10687 ( .I0(ram[7006]), .I1(ram[6998]), .I2(ram[6990]), .I3(
        ram[6982]), .S0(n27277), .S1(n26802), .ZN(n25006) );
  MUX41 U10688 ( .I0(ram[7134]), .I1(ram[7126]), .I2(ram[7118]), .I3(
        ram[7110]), .S0(n27277), .S1(n26802), .ZN(n25011) );
  MUX41 U10689 ( .I0(ram[6878]), .I1(ram[6870]), .I2(ram[6862]), .I3(
        ram[6854]), .S0(n27276), .S1(n26801), .ZN(n25001) );
  MUX41 U10690 ( .I0(ram[6750]), .I1(ram[6742]), .I2(ram[6734]), .I3(
        ram[6726]), .S0(n27276), .S1(n26801), .ZN(n24996) );
  MUX41 U10691 ( .I0(ram[5470]), .I1(ram[5462]), .I2(ram[5454]), .I3(
        ram[5446]), .S0(n27273), .S1(n26798), .ZN(n24941) );
  MUX41 U10692 ( .I0(ram[5598]), .I1(ram[5590]), .I2(ram[5582]), .I3(
        ram[5574]), .S0(n27273), .S1(n26798), .ZN(n24946) );
  MUX41 U10693 ( .I0(ram[5342]), .I1(ram[5334]), .I2(ram[5326]), .I3(
        ram[5318]), .S0(n27273), .S1(n26798), .ZN(n24936) );
  MUX41 U10694 ( .I0(ram[5214]), .I1(ram[5206]), .I2(ram[5198]), .I3(
        ram[5190]), .S0(n27272), .S1(n26797), .ZN(n24931) );
  MUX41 U10695 ( .I0(ram[5982]), .I1(ram[5974]), .I2(ram[5966]), .I3(
        ram[5958]), .S0(n27274), .S1(n26799), .ZN(n24961) );
  MUX41 U10696 ( .I0(ram[6110]), .I1(ram[6102]), .I2(ram[6094]), .I3(
        ram[6086]), .S0(n27274), .S1(n26799), .ZN(n24966) );
  MUX41 U10697 ( .I0(ram[5854]), .I1(ram[5846]), .I2(ram[5838]), .I3(
        ram[5830]), .S0(n27274), .S1(n26799), .ZN(n24956) );
  MUX41 U10698 ( .I0(ram[5726]), .I1(ram[5718]), .I2(ram[5710]), .I3(
        ram[5702]), .S0(n27273), .S1(n26798), .ZN(n24951) );
  MUX41 U10699 ( .I0(ram[4446]), .I1(ram[4438]), .I2(ram[4430]), .I3(
        ram[4422]), .S0(n27270), .S1(n26795), .ZN(n24901) );
  MUX41 U10700 ( .I0(ram[4574]), .I1(ram[4566]), .I2(ram[4558]), .I3(
        ram[4550]), .S0(n27271), .S1(n26796), .ZN(n24906) );
  MUX41 U10701 ( .I0(ram[4958]), .I1(ram[4950]), .I2(ram[4942]), .I3(
        ram[4934]), .S0(n27272), .S1(n26797), .ZN(n24921) );
  MUX41 U10702 ( .I0(ram[11614]), .I1(ram[11606]), .I2(ram[11598]), .I3(
        ram[11590]), .S0(n27288), .S1(n26813), .ZN(n25197) );
  MUX41 U10703 ( .I0(ram[11742]), .I1(ram[11734]), .I2(ram[11726]), .I3(
        ram[11718]), .S0(n27288), .S1(n26813), .ZN(n25202) );
  MUX41 U10704 ( .I0(ram[11486]), .I1(ram[11478]), .I2(ram[11470]), .I3(
        ram[11462]), .S0(n27287), .S1(n26812), .ZN(n25192) );
  MUX41 U10705 ( .I0(ram[11358]), .I1(ram[11350]), .I2(ram[11342]), .I3(
        ram[11334]), .S0(n27287), .S1(n26812), .ZN(n25187) );
  MUX41 U10706 ( .I0(ram[12126]), .I1(ram[12118]), .I2(ram[12110]), .I3(
        ram[12102]), .S0(n27289), .S1(n26814), .ZN(n25217) );
  MUX41 U10707 ( .I0(ram[12254]), .I1(ram[12246]), .I2(ram[12238]), .I3(
        ram[12230]), .S0(n27289), .S1(n26814), .ZN(n25222) );
  MUX41 U10708 ( .I0(ram[11998]), .I1(ram[11990]), .I2(ram[11982]), .I3(
        ram[11974]), .S0(n27289), .S1(n26814), .ZN(n25212) );
  MUX41 U10709 ( .I0(ram[11870]), .I1(ram[11862]), .I2(ram[11854]), .I3(
        ram[11846]), .S0(n27288), .S1(n26813), .ZN(n25207) );
  MUX41 U10710 ( .I0(ram[10590]), .I1(ram[10582]), .I2(ram[10574]), .I3(
        ram[10566]), .S0(n27285), .S1(n26810), .ZN(n25157) );
  MUX41 U10711 ( .I0(ram[10718]), .I1(ram[10710]), .I2(ram[10702]), .I3(
        ram[10694]), .S0(n27285), .S1(n26810), .ZN(n25162) );
  MUX41 U10712 ( .I0(ram[10462]), .I1(ram[10454]), .I2(ram[10446]), .I3(
        ram[10438]), .S0(n27285), .S1(n26810), .ZN(n25152) );
  MUX41 U10713 ( .I0(ram[10334]), .I1(ram[10326]), .I2(ram[10318]), .I3(
        ram[10310]), .S0(n27285), .S1(n26810), .ZN(n25147) );
  MUX41 U10714 ( .I0(ram[11102]), .I1(ram[11094]), .I2(ram[11086]), .I3(
        ram[11078]), .S0(n27286), .S1(n26811), .ZN(n25177) );
  MUX41 U10715 ( .I0(ram[11230]), .I1(ram[11222]), .I2(ram[11214]), .I3(
        ram[11206]), .S0(n27287), .S1(n26812), .ZN(n25182) );
  MUX41 U10716 ( .I0(ram[10974]), .I1(ram[10966]), .I2(ram[10958]), .I3(
        ram[10950]), .S0(n27286), .S1(n26811), .ZN(n25172) );
  MUX41 U10717 ( .I0(ram[9566]), .I1(ram[9558]), .I2(ram[9550]), .I3(
        ram[9542]), .S0(n27283), .S1(n26808), .ZN(n25112) );
  MUX41 U10718 ( .I0(ram[9694]), .I1(ram[9686]), .I2(ram[9678]), .I3(
        ram[9670]), .S0(n27283), .S1(n26808), .ZN(n25117) );
  MUX41 U10719 ( .I0(ram[9438]), .I1(ram[9430]), .I2(ram[9422]), .I3(
        ram[9414]), .S0(n27282), .S1(n26807), .ZN(n25107) );
  MUX41 U10720 ( .I0(ram[9310]), .I1(ram[9302]), .I2(ram[9294]), .I3(
        ram[9286]), .S0(n27282), .S1(n26807), .ZN(n25102) );
  MUX41 U10721 ( .I0(ram[10078]), .I1(ram[10070]), .I2(ram[10062]), .I3(
        ram[10054]), .S0(n27284), .S1(n26809), .ZN(n25132) );
  MUX41 U10722 ( .I0(ram[10206]), .I1(ram[10198]), .I2(ram[10190]), .I3(
        ram[10182]), .S0(n27284), .S1(n26809), .ZN(n25137) );
  MUX41 U10723 ( .I0(ram[9950]), .I1(ram[9942]), .I2(ram[9934]), .I3(
        ram[9926]), .S0(n27284), .S1(n26809), .ZN(n25127) );
  MUX41 U10724 ( .I0(ram[9822]), .I1(ram[9814]), .I2(ram[9806]), .I3(
        ram[9798]), .S0(n27283), .S1(n26808), .ZN(n25122) );
  MUX41 U10725 ( .I0(ram[8542]), .I1(ram[8534]), .I2(ram[8526]), .I3(
        ram[8518]), .S0(n27280), .S1(n26805), .ZN(n25072) );
  MUX41 U10726 ( .I0(ram[8670]), .I1(ram[8662]), .I2(ram[8654]), .I3(
        ram[8646]), .S0(n27281), .S1(n26806), .ZN(n25077) );
  MUX41 U10727 ( .I0(ram[8414]), .I1(ram[8406]), .I2(ram[8398]), .I3(
        ram[8390]), .S0(n27280), .S1(n26805), .ZN(n25067) );
  MUX41 U10728 ( .I0(ram[8286]), .I1(ram[8278]), .I2(ram[8270]), .I3(
        ram[8262]), .S0(n27280), .S1(n26805), .ZN(n25062) );
  MUX41 U10729 ( .I0(ram[9054]), .I1(ram[9046]), .I2(ram[9038]), .I3(
        ram[9030]), .S0(n27281), .S1(n26806), .ZN(n25092) );
  MUX41 U10730 ( .I0(ram[9182]), .I1(ram[9174]), .I2(ram[9166]), .I3(
        ram[9158]), .S0(n27282), .S1(n26807), .ZN(n25097) );
  MUX41 U10731 ( .I0(ram[15711]), .I1(ram[15703]), .I2(ram[15695]), .I3(
        ram[15687]), .S0(n27337), .S1(n26862), .ZN(n26052) );
  MUX41 U10732 ( .I0(ram[15839]), .I1(ram[15831]), .I2(ram[15823]), .I3(
        ram[15815]), .S0(n27337), .S1(n26862), .ZN(n26057) );
  MUX41 U10733 ( .I0(ram[15583]), .I1(ram[15575]), .I2(ram[15567]), .I3(
        ram[15559]), .S0(n27337), .S1(n26862), .ZN(n26047) );
  MUX41 U10734 ( .I0(ram[15455]), .I1(ram[15447]), .I2(ram[15439]), .I3(
        ram[15431]), .S0(n27336), .S1(n26861), .ZN(n26042) );
  MUX41 U10735 ( .I0(ram[16223]), .I1(ram[16215]), .I2(ram[16207]), .I3(
        ram[16199]), .S0(n27338), .S1(n26863), .ZN(n26072) );
  MUX41 U10736 ( .I0(ram[16351]), .I1(ram[16343]), .I2(ram[16335]), .I3(
        ram[16327]), .S0(n27338), .S1(n26863), .ZN(n26077) );
  MUX41 U10737 ( .I0(ram[15967]), .I1(ram[15959]), .I2(ram[15951]), .I3(
        ram[15943]), .S0(n27337), .S1(n26862), .ZN(n26062) );
  MUX41 U10738 ( .I0(ram[16095]), .I1(ram[16087]), .I2(ram[16079]), .I3(
        ram[16071]), .S0(n27338), .S1(n26863), .ZN(n26067) );
  MUX41 U10739 ( .I0(ram[15199]), .I1(ram[15191]), .I2(ram[15183]), .I3(
        ram[15175]), .S0(n27336), .S1(n26861), .ZN(n26032) );
  MUX41 U10740 ( .I0(ram[15327]), .I1(ram[15319]), .I2(ram[15311]), .I3(
        ram[15303]), .S0(n27336), .S1(n26861), .ZN(n26037) );
  MUX41 U10741 ( .I0(ram[15071]), .I1(ram[15063]), .I2(ram[15055]), .I3(
        ram[15047]), .S0(n27335), .S1(n26860), .ZN(n26027) );
  MUX41 U10742 ( .I0(ram[14943]), .I1(ram[14935]), .I2(ram[14927]), .I3(
        ram[14919]), .S0(n27335), .S1(n26860), .ZN(n26022) );
  MUX41 U10743 ( .I0(ram[14687]), .I1(ram[14679]), .I2(ram[14671]), .I3(
        ram[14663]), .S0(n27334), .S1(n26859), .ZN(n26012) );
  MUX41 U10744 ( .I0(ram[14815]), .I1(ram[14807]), .I2(ram[14799]), .I3(
        ram[14791]), .S0(n27335), .S1(n26860), .ZN(n26017) );
  MUX41 U10745 ( .I0(ram[14559]), .I1(ram[14551]), .I2(ram[14543]), .I3(
        ram[14535]), .S0(n27334), .S1(n26859), .ZN(n26007) );
  MUX41 U10746 ( .I0(ram[14431]), .I1(ram[14423]), .I2(ram[14415]), .I3(
        ram[14407]), .S0(n27334), .S1(n26859), .ZN(n26002) );
  MUX41 U10747 ( .I0(ram[13663]), .I1(ram[13655]), .I2(ram[13647]), .I3(
        ram[13639]), .S0(n27332), .S1(n26857), .ZN(n25967) );
  MUX41 U10748 ( .I0(ram[13791]), .I1(ram[13783]), .I2(ram[13775]), .I3(
        ram[13767]), .S0(n27332), .S1(n26857), .ZN(n25972) );
  MUX41 U10749 ( .I0(ram[13535]), .I1(ram[13527]), .I2(ram[13519]), .I3(
        ram[13511]), .S0(n27332), .S1(n26857), .ZN(n25962) );
  MUX41 U10750 ( .I0(ram[13407]), .I1(ram[13399]), .I2(ram[13391]), .I3(
        ram[13383]), .S0(n27331), .S1(n26856), .ZN(n25957) );
  MUX41 U10751 ( .I0(ram[14175]), .I1(ram[14167]), .I2(ram[14159]), .I3(
        ram[14151]), .S0(n27333), .S1(n26858), .ZN(n25987) );
  MUX41 U10752 ( .I0(ram[14303]), .I1(ram[14295]), .I2(ram[14287]), .I3(
        ram[14279]), .S0(n27333), .S1(n26858), .ZN(n25992) );
  MUX41 U10753 ( .I0(ram[14047]), .I1(ram[14039]), .I2(ram[14031]), .I3(
        ram[14023]), .S0(n27333), .S1(n26858), .ZN(n25982) );
  MUX41 U10754 ( .I0(ram[13919]), .I1(ram[13911]), .I2(ram[13903]), .I3(
        ram[13895]), .S0(n27333), .S1(n26858), .ZN(n25977) );
  MUX41 U10755 ( .I0(ram[13151]), .I1(ram[13143]), .I2(ram[13135]), .I3(
        ram[13127]), .S0(n27331), .S1(n26856), .ZN(n25947) );
  MUX41 U10756 ( .I0(ram[13279]), .I1(ram[13271]), .I2(ram[13263]), .I3(
        ram[13255]), .S0(n27331), .S1(n26856), .ZN(n25952) );
  MUX41 U10757 ( .I0(ram[13023]), .I1(ram[13015]), .I2(ram[13007]), .I3(
        ram[12999]), .S0(n27330), .S1(n26855), .ZN(n25942) );
  MUX41 U10758 ( .I0(ram[12895]), .I1(ram[12887]), .I2(ram[12879]), .I3(
        ram[12871]), .S0(n27330), .S1(n26855), .ZN(n25937) );
  MUX41 U10759 ( .I0(ram[12639]), .I1(ram[12631]), .I2(ram[12623]), .I3(
        ram[12615]), .S0(n27329), .S1(n26854), .ZN(n25927) );
  MUX41 U10760 ( .I0(ram[12767]), .I1(ram[12759]), .I2(ram[12751]), .I3(
        ram[12743]), .S0(n27330), .S1(n26855), .ZN(n25932) );
  MUX41 U10761 ( .I0(ram[12511]), .I1(ram[12503]), .I2(ram[12495]), .I3(
        ram[12487]), .S0(n27329), .S1(n26854), .ZN(n25922) );
  MUX41 U10762 ( .I0(ram[12383]), .I1(ram[12375]), .I2(ram[12367]), .I3(
        ram[12359]), .S0(n27329), .S1(n26854), .ZN(n25917) );
  MUX41 U10763 ( .I0(n25537), .I1(n25538), .I2(n25539), .I3(n25540), .S0(
        n26265), .S1(n26383), .ZN(n25536) );
  MUX41 U10764 ( .I0(ram[3391]), .I1(ram[3383]), .I2(ram[3375]), .I3(
        ram[3367]), .S0(n27307), .S1(n26832), .ZN(n25538) );
  MUX41 U10765 ( .I0(ram[3359]), .I1(ram[3351]), .I2(ram[3343]), .I3(
        ram[3335]), .S0(n27307), .S1(n26832), .ZN(n25540) );
  MUX41 U10766 ( .I0(ram[3455]), .I1(ram[3447]), .I2(ram[3439]), .I3(
        ram[3431]), .S0(n27307), .S1(n26832), .ZN(n25537) );
  MUX41 U10767 ( .I0(n25557), .I1(n25558), .I2(n25559), .I3(n25560), .S0(
        n26265), .S1(n26383), .ZN(n25556) );
  MUX41 U10768 ( .I0(ram[3903]), .I1(ram[3895]), .I2(ram[3887]), .I3(
        ram[3879]), .S0(n27308), .S1(n26833), .ZN(n25558) );
  MUX41 U10769 ( .I0(ram[3871]), .I1(ram[3863]), .I2(ram[3855]), .I3(
        ram[3847]), .S0(n27308), .S1(n26833), .ZN(n25560) );
  MUX41 U10770 ( .I0(ram[3967]), .I1(ram[3959]), .I2(ram[3951]), .I3(
        ram[3943]), .S0(n27309), .S1(n26834), .ZN(n25557) );
  MUX41 U10771 ( .I0(n25497), .I1(n25498), .I2(n25499), .I3(n25500), .S0(
        n26264), .S1(n26382), .ZN(n25496) );
  MUX41 U10772 ( .I0(ram[2335]), .I1(ram[2327]), .I2(ram[2319]), .I3(
        ram[2311]), .S0(n27305), .S1(n26830), .ZN(n25500) );
  MUX41 U10773 ( .I0(ram[2367]), .I1(ram[2359]), .I2(ram[2351]), .I3(
        ram[2343]), .S0(n27305), .S1(n26830), .ZN(n25498) );
  MUX41 U10774 ( .I0(ram[2431]), .I1(ram[2423]), .I2(ram[2415]), .I3(
        ram[2407]), .S0(n27305), .S1(n26830), .ZN(n25497) );
  MUX41 U10775 ( .I0(n25517), .I1(n25518), .I2(n25519), .I3(n25520), .S0(
        n26264), .S1(n26382), .ZN(n25516) );
  MUX41 U10776 ( .I0(ram[2847]), .I1(ram[2839]), .I2(ram[2831]), .I3(
        ram[2823]), .S0(n27306), .S1(n26831), .ZN(n25520) );
  MUX41 U10777 ( .I0(ram[2879]), .I1(ram[2871]), .I2(ram[2863]), .I3(
        ram[2855]), .S0(n27306), .S1(n26831), .ZN(n25518) );
  MUX41 U10778 ( .I0(ram[2943]), .I1(ram[2935]), .I2(ram[2927]), .I3(
        ram[2919]), .S0(n27306), .S1(n26831), .ZN(n25517) );
  MUX41 U10779 ( .I0(n25452), .I1(n25453), .I2(n25454), .I3(n25455), .S0(
        n26263), .S1(n26381), .ZN(n25451) );
  MUX41 U10780 ( .I0(ram[1343]), .I1(ram[1335]), .I2(ram[1327]), .I3(
        ram[1319]), .S0(n27302), .S1(n26827), .ZN(n25453) );
  MUX41 U10781 ( .I0(ram[1311]), .I1(ram[1303]), .I2(ram[1295]), .I3(
        ram[1287]), .S0(n27302), .S1(n26827), .ZN(n25455) );
  MUX41 U10782 ( .I0(ram[1407]), .I1(ram[1399]), .I2(ram[1391]), .I3(
        ram[1383]), .S0(n27302), .S1(n26827), .ZN(n25452) );
  MUX41 U10783 ( .I0(n25472), .I1(n25473), .I2(n25474), .I3(n25475), .S0(
        n26264), .S1(n26382), .ZN(n25471) );
  MUX41 U10784 ( .I0(ram[1823]), .I1(ram[1815]), .I2(ram[1807]), .I3(
        ram[1799]), .S0(n27303), .S1(n26828), .ZN(n25475) );
  MUX41 U10785 ( .I0(ram[1855]), .I1(ram[1847]), .I2(ram[1839]), .I3(
        ram[1831]), .S0(n27304), .S1(n26829), .ZN(n25473) );
  MUX41 U10786 ( .I0(ram[1919]), .I1(ram[1911]), .I2(ram[1903]), .I3(
        ram[1895]), .S0(n27304), .S1(n26829), .ZN(n25472) );
  MUX41 U10787 ( .I0(n25412), .I1(n25413), .I2(n25414), .I3(n25415), .S0(
        n26263), .S1(n26381), .ZN(n25411) );
  MUX41 U10788 ( .I0(ram[287]), .I1(ram[279]), .I2(ram[271]), .I3(
        ram[263]), .S0(n27300), .S1(n26825), .ZN(n25415) );
  MUX41 U10789 ( .I0(ram[319]), .I1(ram[311]), .I2(ram[303]), .I3(
        ram[295]), .S0(n27300), .S1(n26825), .ZN(n25413) );
  MUX41 U10790 ( .I0(ram[383]), .I1(ram[375]), .I2(ram[367]), .I3(
        ram[359]), .S0(n27300), .S1(n26825), .ZN(n25412) );
  MUX41 U10791 ( .I0(n25432), .I1(n25433), .I2(n25434), .I3(n25435), .S0(
        n26263), .S1(n26381), .ZN(n25431) );
  MUX41 U10792 ( .I0(ram[799]), .I1(ram[791]), .I2(ram[783]), .I3(
        ram[775]), .S0(n27301), .S1(n26826), .ZN(n25435) );
  MUX41 U10793 ( .I0(ram[831]), .I1(ram[823]), .I2(ram[815]), .I3(
        ram[807]), .S0(n27301), .S1(n26826), .ZN(n25433) );
  MUX41 U10794 ( .I0(ram[895]), .I1(ram[887]), .I2(ram[879]), .I3(
        ram[871]), .S0(n27301), .S1(n26826), .ZN(n25432) );
  MUX41 U10795 ( .I0(ram[7519]), .I1(ram[7511]), .I2(ram[7503]), .I3(
        ram[7495]), .S0(n27317), .S1(n26842), .ZN(n25710) );
  MUX41 U10796 ( .I0(ram[7647]), .I1(ram[7639]), .I2(ram[7631]), .I3(
        ram[7623]), .S0(n27317), .S1(n26842), .ZN(n25715) );
  MUX41 U10797 ( .I0(ram[7391]), .I1(ram[7383]), .I2(ram[7375]), .I3(
        ram[7367]), .S0(n27317), .S1(n26842), .ZN(n25705) );
  MUX41 U10798 ( .I0(ram[7263]), .I1(ram[7255]), .I2(ram[7247]), .I3(
        ram[7239]), .S0(n27317), .S1(n26842), .ZN(n25700) );
  MUX41 U10799 ( .I0(ram[8031]), .I1(ram[8023]), .I2(ram[8015]), .I3(
        ram[8007]), .S0(n27318), .S1(n26843), .ZN(n25730) );
  MUX41 U10800 ( .I0(ram[8159]), .I1(ram[8151]), .I2(ram[8143]), .I3(
        ram[8135]), .S0(n27319), .S1(n26844), .ZN(n25735) );
  MUX41 U10801 ( .I0(ram[7903]), .I1(ram[7895]), .I2(ram[7887]), .I3(
        ram[7879]), .S0(n27318), .S1(n26843), .ZN(n25725) );
  MUX41 U10802 ( .I0(ram[7775]), .I1(ram[7767]), .I2(ram[7759]), .I3(
        ram[7751]), .S0(n27318), .S1(n26843), .ZN(n25720) );
  MUX41 U10803 ( .I0(ram[6495]), .I1(ram[6487]), .I2(ram[6479]), .I3(
        ram[6471]), .S0(n27315), .S1(n26840), .ZN(n25670) );
  MUX41 U10804 ( .I0(ram[6623]), .I1(ram[6615]), .I2(ram[6607]), .I3(
        ram[6599]), .S0(n27315), .S1(n26840), .ZN(n25675) );
  MUX41 U10805 ( .I0(ram[6367]), .I1(ram[6359]), .I2(ram[6351]), .I3(
        ram[6343]), .S0(n27314), .S1(n26839), .ZN(n25665) );
  MUX41 U10806 ( .I0(ram[6239]), .I1(ram[6231]), .I2(ram[6223]), .I3(
        ram[6215]), .S0(n27314), .S1(n26839), .ZN(n25660) );
  MUX41 U10807 ( .I0(ram[7007]), .I1(ram[6999]), .I2(ram[6991]), .I3(
        ram[6983]), .S0(n27316), .S1(n26841), .ZN(n25690) );
  MUX41 U10808 ( .I0(ram[7135]), .I1(ram[7127]), .I2(ram[7119]), .I3(
        ram[7111]), .S0(n27316), .S1(n26841), .ZN(n25695) );
  MUX41 U10809 ( .I0(ram[6879]), .I1(ram[6871]), .I2(ram[6863]), .I3(
        ram[6855]), .S0(n27316), .S1(n26841), .ZN(n25685) );
  MUX41 U10810 ( .I0(ram[6751]), .I1(ram[6743]), .I2(ram[6735]), .I3(
        ram[6727]), .S0(n27315), .S1(n26840), .ZN(n25680) );
  MUX41 U10811 ( .I0(ram[5471]), .I1(ram[5463]), .I2(ram[5455]), .I3(
        ram[5447]), .S0(n27312), .S1(n26837), .ZN(n25625) );
  MUX41 U10812 ( .I0(ram[5599]), .I1(ram[5591]), .I2(ram[5583]), .I3(
        ram[5575]), .S0(n27313), .S1(n26838), .ZN(n25630) );
  MUX41 U10813 ( .I0(ram[5343]), .I1(ram[5335]), .I2(ram[5327]), .I3(
        ram[5319]), .S0(n27312), .S1(n26837), .ZN(n25620) );
  MUX41 U10814 ( .I0(ram[5215]), .I1(ram[5207]), .I2(ram[5199]), .I3(
        ram[5191]), .S0(n27312), .S1(n26837), .ZN(n25615) );
  MUX41 U10815 ( .I0(ram[5983]), .I1(ram[5975]), .I2(ram[5967]), .I3(
        ram[5959]), .S0(n27313), .S1(n26838), .ZN(n25645) );
  MUX41 U10816 ( .I0(ram[6111]), .I1(ram[6103]), .I2(ram[6095]), .I3(
        ram[6087]), .S0(n27314), .S1(n26839), .ZN(n25650) );
  MUX41 U10817 ( .I0(ram[5855]), .I1(ram[5847]), .I2(ram[5839]), .I3(
        ram[5831]), .S0(n27313), .S1(n26838), .ZN(n25640) );
  MUX41 U10818 ( .I0(ram[5727]), .I1(ram[5719]), .I2(ram[5711]), .I3(
        ram[5703]), .S0(n27313), .S1(n26838), .ZN(n25635) );
  MUX41 U10819 ( .I0(ram[4447]), .I1(ram[4439]), .I2(ram[4431]), .I3(
        ram[4423]), .S0(n27310), .S1(n26835), .ZN(n25585) );
  MUX41 U10820 ( .I0(ram[4575]), .I1(ram[4567]), .I2(ram[4559]), .I3(
        ram[4551]), .S0(n27310), .S1(n26835), .ZN(n25590) );
  MUX41 U10821 ( .I0(ram[4959]), .I1(ram[4951]), .I2(ram[4943]), .I3(
        ram[4935]), .S0(n27311), .S1(n26836), .ZN(n25605) );
  MUX41 U10822 ( .I0(ram[11615]), .I1(ram[11607]), .I2(ram[11599]), .I3(
        ram[11591]), .S0(n27327), .S1(n26852), .ZN(n25881) );
  MUX41 U10823 ( .I0(ram[11743]), .I1(ram[11735]), .I2(ram[11727]), .I3(
        ram[11719]), .S0(n27327), .S1(n26852), .ZN(n25886) );
  MUX41 U10824 ( .I0(ram[11487]), .I1(ram[11479]), .I2(ram[11471]), .I3(
        ram[11463]), .S0(n27327), .S1(n26852), .ZN(n25876) );
  MUX41 U10825 ( .I0(ram[11359]), .I1(ram[11351]), .I2(ram[11343]), .I3(
        ram[11335]), .S0(n27326), .S1(n26851), .ZN(n25871) );
  MUX41 U10826 ( .I0(ram[12127]), .I1(ram[12119]), .I2(ram[12111]), .I3(
        ram[12103]), .S0(n27328), .S1(n26853), .ZN(n25901) );
  MUX41 U10827 ( .I0(ram[12255]), .I1(ram[12247]), .I2(ram[12239]), .I3(
        ram[12231]), .S0(n27329), .S1(n26854), .ZN(n25906) );
  MUX41 U10828 ( .I0(ram[11999]), .I1(ram[11991]), .I2(ram[11983]), .I3(
        ram[11975]), .S0(n27328), .S1(n26853), .ZN(n25896) );
  MUX41 U10829 ( .I0(ram[11871]), .I1(ram[11863]), .I2(ram[11855]), .I3(
        ram[11847]), .S0(n27328), .S1(n26853), .ZN(n25891) );
  MUX41 U10830 ( .I0(ram[10591]), .I1(ram[10583]), .I2(ram[10575]), .I3(
        ram[10567]), .S0(n27325), .S1(n26850), .ZN(n25841) );
  MUX41 U10831 ( .I0(ram[10719]), .I1(ram[10711]), .I2(ram[10703]), .I3(
        ram[10695]), .S0(n27325), .S1(n26850), .ZN(n25846) );
  MUX41 U10832 ( .I0(ram[10463]), .I1(ram[10455]), .I2(ram[10447]), .I3(
        ram[10439]), .S0(n27324), .S1(n26849), .ZN(n25836) );
  MUX41 U10833 ( .I0(ram[10335]), .I1(ram[10327]), .I2(ram[10319]), .I3(
        ram[10311]), .S0(n27324), .S1(n26849), .ZN(n25831) );
  MUX41 U10834 ( .I0(ram[11103]), .I1(ram[11095]), .I2(ram[11087]), .I3(
        ram[11079]), .S0(n27326), .S1(n26851), .ZN(n25861) );
  MUX41 U10835 ( .I0(ram[11231]), .I1(ram[11223]), .I2(ram[11215]), .I3(
        ram[11207]), .S0(n27326), .S1(n26851), .ZN(n25866) );
  MUX41 U10836 ( .I0(ram[10975]), .I1(ram[10967]), .I2(ram[10959]), .I3(
        ram[10951]), .S0(n27325), .S1(n26850), .ZN(n25856) );
  MUX41 U10837 ( .I0(ram[9567]), .I1(ram[9559]), .I2(ram[9551]), .I3(
        ram[9543]), .S0(n27322), .S1(n26847), .ZN(n25796) );
  MUX41 U10838 ( .I0(ram[9695]), .I1(ram[9687]), .I2(ram[9679]), .I3(
        ram[9671]), .S0(n27322), .S1(n26847), .ZN(n25801) );
  MUX41 U10839 ( .I0(ram[9439]), .I1(ram[9431]), .I2(ram[9423]), .I3(
        ram[9415]), .S0(n27322), .S1(n26847), .ZN(n25791) );
  MUX41 U10840 ( .I0(ram[9311]), .I1(ram[9303]), .I2(ram[9295]), .I3(
        ram[9287]), .S0(n27321), .S1(n26846), .ZN(n25786) );
  MUX41 U10841 ( .I0(ram[10079]), .I1(ram[10071]), .I2(ram[10063]), .I3(
        ram[10055]), .S0(n27323), .S1(n26848), .ZN(n25816) );
  MUX41 U10842 ( .I0(ram[10207]), .I1(ram[10199]), .I2(ram[10191]), .I3(
        ram[10183]), .S0(n27324), .S1(n26849), .ZN(n25821) );
  MUX41 U10843 ( .I0(ram[9951]), .I1(ram[9943]), .I2(ram[9935]), .I3(
        ram[9927]), .S0(n27323), .S1(n26848), .ZN(n25811) );
  MUX41 U10844 ( .I0(ram[9823]), .I1(ram[9815]), .I2(ram[9807]), .I3(
        ram[9799]), .S0(n27323), .S1(n26848), .ZN(n25806) );
  MUX41 U10845 ( .I0(ram[8543]), .I1(ram[8535]), .I2(ram[8527]), .I3(
        ram[8519]), .S0(n27320), .S1(n26845), .ZN(n25756) );
  MUX41 U10846 ( .I0(ram[8671]), .I1(ram[8663]), .I2(ram[8655]), .I3(
        ram[8647]), .S0(n27320), .S1(n26845), .ZN(n25761) );
  MUX41 U10847 ( .I0(ram[8415]), .I1(ram[8407]), .I2(ram[8399]), .I3(
        ram[8391]), .S0(n27319), .S1(n26844), .ZN(n25751) );
  MUX41 U10848 ( .I0(ram[8287]), .I1(ram[8279]), .I2(ram[8271]), .I3(
        ram[8263]), .S0(n27319), .S1(n26844), .ZN(n25746) );
  MUX41 U10849 ( .I0(ram[9055]), .I1(ram[9047]), .I2(ram[9039]), .I3(
        ram[9031]), .S0(n27321), .S1(n26846), .ZN(n25776) );
  MUX41 U10850 ( .I0(ram[9183]), .I1(ram[9175]), .I2(ram[9167]), .I3(
        ram[9159]), .S0(n27321), .S1(n26846), .ZN(n25781) );
  MUX41 U10851 ( .I0(n21262), .I1(n21263), .I2(n21264), .I3(n21265), .S0(
        n26203), .S1(n26321), .ZN(n21261) );
  MUX41 U10852 ( .I0(ram[15640]), .I1(ram[15632]), .I2(ram[15624]), .I3(
        ram[15616]), .S0(n27061), .S1(n26586), .ZN(n21265) );
  MUX41 U10853 ( .I0(ram[15672]), .I1(ram[15664]), .I2(ram[15656]), .I3(
        ram[15648]), .S0(n27061), .S1(n26586), .ZN(n21263) );
  MUX41 U10854 ( .I0(ram[15736]), .I1(ram[15728]), .I2(ram[15720]), .I3(
        ram[15712]), .S0(n27061), .S1(n26586), .ZN(n21262) );
  MUX41 U10855 ( .I0(n21282), .I1(n21283), .I2(n21284), .I3(n21285), .S0(
        n26203), .S1(n26321), .ZN(n21281) );
  MUX41 U10856 ( .I0(ram[16152]), .I1(ram[16144]), .I2(ram[16136]), .I3(
        ram[16128]), .S0(n27062), .S1(n26587), .ZN(n21285) );
  MUX41 U10857 ( .I0(ram[16184]), .I1(ram[16176]), .I2(ram[16168]), .I3(
        ram[16160]), .S0(n27062), .S1(n26587), .ZN(n21283) );
  MUX41 U10858 ( .I0(ram[16248]), .I1(ram[16240]), .I2(ram[16232]), .I3(
        ram[16224]), .S0(n27062), .S1(n26587), .ZN(n21282) );
  MUX41 U10859 ( .I0(n21242), .I1(n21243), .I2(n21244), .I3(n21245), .S0(
        n26203), .S1(n26321), .ZN(n21241) );
  MUX41 U10860 ( .I0(ram[15128]), .I1(ram[15120]), .I2(ram[15112]), .I3(
        ram[15104]), .S0(n27060), .S1(n26585), .ZN(n21245) );
  MUX41 U10861 ( .I0(ram[15160]), .I1(ram[15152]), .I2(ram[15144]), .I3(
        ram[15136]), .S0(n27060), .S1(n26585), .ZN(n21243) );
  MUX41 U10862 ( .I0(ram[15224]), .I1(ram[15216]), .I2(ram[15208]), .I3(
        ram[15200]), .S0(n27060), .S1(n26585), .ZN(n21242) );
  MUX41 U10863 ( .I0(n21222), .I1(n21223), .I2(n21224), .I3(n21225), .S0(
        n26203), .S1(n26321), .ZN(n21221) );
  MUX41 U10864 ( .I0(ram[14616]), .I1(ram[14608]), .I2(ram[14600]), .I3(
        ram[14592]), .S0(n27059), .S1(n26584), .ZN(n21225) );
  MUX41 U10865 ( .I0(ram[14648]), .I1(ram[14640]), .I2(ram[14632]), .I3(
        ram[14624]), .S0(n27059), .S1(n26584), .ZN(n21223) );
  MUX41 U10866 ( .I0(ram[14712]), .I1(ram[14704]), .I2(ram[14696]), .I3(
        ram[14688]), .S0(n27059), .S1(n26584), .ZN(n21222) );
  MUX41 U10867 ( .I0(n21177), .I1(n21178), .I2(n21179), .I3(n21180), .S0(
        n26202), .S1(n26320), .ZN(n21176) );
  MUX41 U10868 ( .I0(ram[13592]), .I1(ram[13584]), .I2(ram[13576]), .I3(
        ram[13568]), .S0(n27056), .S1(n26581), .ZN(n21180) );
  MUX41 U10869 ( .I0(ram[13624]), .I1(ram[13616]), .I2(ram[13608]), .I3(
        ram[13600]), .S0(n27056), .S1(n26581), .ZN(n21178) );
  MUX41 U10870 ( .I0(ram[13688]), .I1(ram[13680]), .I2(ram[13672]), .I3(
        ram[13664]), .S0(n27056), .S1(n26581), .ZN(n21177) );
  MUX41 U10871 ( .I0(n21197), .I1(n21198), .I2(n21199), .I3(n21200), .S0(
        n26202), .S1(n26320), .ZN(n21196) );
  MUX41 U10872 ( .I0(ram[14104]), .I1(ram[14096]), .I2(ram[14088]), .I3(
        ram[14080]), .S0(n27057), .S1(n26582), .ZN(n21200) );
  MUX41 U10873 ( .I0(ram[14136]), .I1(ram[14128]), .I2(ram[14120]), .I3(
        ram[14112]), .S0(n27057), .S1(n26582), .ZN(n21198) );
  MUX41 U10874 ( .I0(ram[14200]), .I1(ram[14192]), .I2(ram[14184]), .I3(
        ram[14176]), .S0(n27058), .S1(n26583), .ZN(n21197) );
  MUX41 U10875 ( .I0(n21157), .I1(n21158), .I2(n21159), .I3(n21160), .S0(
        n26202), .S1(n26320), .ZN(n21156) );
  MUX41 U10876 ( .I0(ram[13080]), .I1(ram[13072]), .I2(ram[13064]), .I3(
        ram[13056]), .S0(n27055), .S1(n26580), .ZN(n21160) );
  MUX41 U10877 ( .I0(ram[13112]), .I1(ram[13104]), .I2(ram[13096]), .I3(
        ram[13088]), .S0(n27055), .S1(n26580), .ZN(n21158) );
  MUX41 U10878 ( .I0(ram[13176]), .I1(ram[13168]), .I2(ram[13160]), .I3(
        ram[13152]), .S0(n27055), .S1(n26580), .ZN(n21157) );
  MUX41 U10879 ( .I0(n21137), .I1(n21138), .I2(n21139), .I3(n21140), .S0(
        n26201), .S1(n26319), .ZN(n21136) );
  MUX41 U10880 ( .I0(ram[12568]), .I1(ram[12560]), .I2(ram[12552]), .I3(
        ram[12544]), .S0(n27054), .S1(n26579), .ZN(n21140) );
  MUX41 U10881 ( .I0(ram[12600]), .I1(ram[12592]), .I2(ram[12584]), .I3(
        ram[12576]), .S0(n27054), .S1(n26579), .ZN(n21138) );
  MUX41 U10882 ( .I0(ram[12664]), .I1(ram[12656]), .I2(ram[12648]), .I3(
        ram[12640]), .S0(n27054), .S1(n26579), .ZN(n21137) );
  MUX41 U10883 ( .I0(n20920), .I1(n20921), .I2(n20922), .I3(n20923), .S0(
        n26198), .S1(n26316), .ZN(n20919) );
  MUX41 U10884 ( .I0(ram[7480]), .I1(ram[7472]), .I2(ram[7464]), .I3(
        ram[7456]), .S0(n27041), .S1(n26566), .ZN(n20921) );
  MUX41 U10885 ( .I0(ram[7448]), .I1(ram[7440]), .I2(ram[7432]), .I3(
        ram[7424]), .S0(n27041), .S1(n26566), .ZN(n20923) );
  MUX41 U10886 ( .I0(ram[7544]), .I1(ram[7536]), .I2(ram[7528]), .I3(
        ram[7520]), .S0(n27042), .S1(n26567), .ZN(n20920) );
  MUX41 U10887 ( .I0(n20940), .I1(n20941), .I2(n20942), .I3(n20943), .S0(
        n26199), .S1(n26317), .ZN(n20939) );
  MUX41 U10888 ( .I0(ram[7960]), .I1(ram[7952]), .I2(ram[7944]), .I3(
        ram[7936]), .S0(n27043), .S1(n26568), .ZN(n20943) );
  MUX41 U10889 ( .I0(ram[7992]), .I1(ram[7984]), .I2(ram[7976]), .I3(
        ram[7968]), .S0(n27043), .S1(n26568), .ZN(n20941) );
  MUX41 U10890 ( .I0(ram[8056]), .I1(ram[8048]), .I2(ram[8040]), .I3(
        ram[8032]), .S0(n27043), .S1(n26568), .ZN(n20940) );
  MUX41 U10891 ( .I0(n20880), .I1(n20881), .I2(n20882), .I3(n20883), .S0(
        n26198), .S1(n26316), .ZN(n20879) );
  MUX41 U10892 ( .I0(ram[6424]), .I1(ram[6416]), .I2(ram[6408]), .I3(
        ram[6400]), .S0(n27039), .S1(n26564), .ZN(n20883) );
  MUX41 U10893 ( .I0(ram[6456]), .I1(ram[6448]), .I2(ram[6440]), .I3(
        ram[6432]), .S0(n27039), .S1(n26564), .ZN(n20881) );
  MUX41 U10894 ( .I0(ram[6520]), .I1(ram[6512]), .I2(ram[6504]), .I3(
        ram[6496]), .S0(n27039), .S1(n26564), .ZN(n20880) );
  MUX41 U10895 ( .I0(n20900), .I1(n20901), .I2(n20902), .I3(n20903), .S0(
        n26198), .S1(n26316), .ZN(n20899) );
  MUX41 U10896 ( .I0(ram[6936]), .I1(ram[6928]), .I2(ram[6920]), .I3(
        ram[6912]), .S0(n27040), .S1(n26565), .ZN(n20903) );
  MUX41 U10897 ( .I0(ram[6968]), .I1(ram[6960]), .I2(ram[6952]), .I3(
        ram[6944]), .S0(n27040), .S1(n26565), .ZN(n20901) );
  MUX41 U10898 ( .I0(ram[7032]), .I1(ram[7024]), .I2(ram[7016]), .I3(
        ram[7008]), .S0(n27040), .S1(n26565), .ZN(n20900) );
  MUX41 U10899 ( .I0(n20835), .I1(n20836), .I2(n20837), .I3(n20838), .S0(
        n26197), .S1(n26315), .ZN(n20834) );
  MUX41 U10900 ( .I0(ram[5432]), .I1(ram[5424]), .I2(ram[5416]), .I3(
        ram[5408]), .S0(n27036), .S1(n26561), .ZN(n20836) );
  MUX41 U10901 ( .I0(ram[5400]), .I1(ram[5392]), .I2(ram[5384]), .I3(
        ram[5376]), .S0(n27036), .S1(n26561), .ZN(n20838) );
  MUX41 U10902 ( .I0(ram[5496]), .I1(ram[5488]), .I2(ram[5480]), .I3(
        ram[5472]), .S0(n27037), .S1(n26562), .ZN(n20835) );
  MUX41 U10903 ( .I0(n20855), .I1(n20856), .I2(n20857), .I3(n20858), .S0(
        n26197), .S1(n26315), .ZN(n20854) );
  MUX41 U10904 ( .I0(ram[5944]), .I1(ram[5936]), .I2(ram[5928]), .I3(
        ram[5920]), .S0(n27038), .S1(n26563), .ZN(n20856) );
  MUX41 U10905 ( .I0(ram[5912]), .I1(ram[5904]), .I2(ram[5896]), .I3(
        ram[5888]), .S0(n27038), .S1(n26563), .ZN(n20858) );
  MUX41 U10906 ( .I0(ram[6008]), .I1(ram[6000]), .I2(ram[5992]), .I3(
        ram[5984]), .S0(n27038), .S1(n26563), .ZN(n20855) );
  MUX41 U10907 ( .I0(n20795), .I1(n20796), .I2(n20797), .I3(n20798), .S0(
        n26196), .S1(n26314), .ZN(n20794) );
  MUX41 U10908 ( .I0(ram[4408]), .I1(ram[4400]), .I2(ram[4392]), .I3(
        ram[4384]), .S0(n27034), .S1(n26559), .ZN(n20796) );
  MUX41 U10909 ( .I0(ram[4376]), .I1(ram[4368]), .I2(ram[4360]), .I3(
        ram[4352]), .S0(n27034), .S1(n26559), .ZN(n20798) );
  MUX41 U10910 ( .I0(ram[4472]), .I1(ram[4464]), .I2(ram[4456]), .I3(
        ram[4448]), .S0(n27034), .S1(n26559), .ZN(n20795) );
  MUX41 U10911 ( .I0(n20815), .I1(n20816), .I2(n20817), .I3(n20818), .S0(
        n26197), .S1(n26315), .ZN(n20814) );
  MUX41 U10912 ( .I0(ram[4888]), .I1(ram[4880]), .I2(ram[4872]), .I3(
        ram[4864]), .S0(n27035), .S1(n26560), .ZN(n20818) );
  MUX41 U10913 ( .I0(ram[4920]), .I1(ram[4912]), .I2(ram[4904]), .I3(
        ram[4896]), .S0(n27035), .S1(n26560), .ZN(n20816) );
  MUX41 U10914 ( .I0(ram[4984]), .I1(ram[4976]), .I2(ram[4968]), .I3(
        ram[4960]), .S0(n27035), .S1(n26560), .ZN(n20815) );
  MUX41 U10915 ( .I0(n21091), .I1(n21092), .I2(n21093), .I3(n21094), .S0(
        n26201), .S1(n26319), .ZN(n21090) );
  MUX41 U10916 ( .I0(ram[11576]), .I1(ram[11568]), .I2(ram[11560]), .I3(
        ram[11552]), .S0(n27051), .S1(n26576), .ZN(n21092) );
  MUX41 U10917 ( .I0(ram[11544]), .I1(ram[11536]), .I2(ram[11528]), .I3(
        ram[11520]), .S0(n27051), .S1(n26576), .ZN(n21094) );
  MUX41 U10918 ( .I0(ram[11640]), .I1(ram[11632]), .I2(ram[11624]), .I3(
        ram[11616]), .S0(n27051), .S1(n26576), .ZN(n21091) );
  MUX41 U10919 ( .I0(n21111), .I1(n21112), .I2(n21113), .I3(n21114), .S0(
        n26201), .S1(n26319), .ZN(n21110) );
  MUX41 U10920 ( .I0(ram[12088]), .I1(ram[12080]), .I2(ram[12072]), .I3(
        ram[12064]), .S0(n27052), .S1(n26577), .ZN(n21112) );
  MUX41 U10921 ( .I0(ram[12056]), .I1(ram[12048]), .I2(ram[12040]), .I3(
        ram[12032]), .S0(n27052), .S1(n26577), .ZN(n21114) );
  MUX41 U10922 ( .I0(ram[12152]), .I1(ram[12144]), .I2(ram[12136]), .I3(
        ram[12128]), .S0(n27053), .S1(n26578), .ZN(n21111) );
  MUX41 U10923 ( .I0(n21051), .I1(n21052), .I2(n21053), .I3(n21054), .S0(
        n26200), .S1(n26318), .ZN(n21050) );
  MUX41 U10924 ( .I0(ram[10552]), .I1(ram[10544]), .I2(ram[10536]), .I3(
        ram[10528]), .S0(n27049), .S1(n26574), .ZN(n21052) );
  MUX41 U10925 ( .I0(ram[10520]), .I1(ram[10512]), .I2(ram[10504]), .I3(
        ram[10496]), .S0(n27049), .S1(n26574), .ZN(n21054) );
  MUX41 U10926 ( .I0(ram[10616]), .I1(ram[10608]), .I2(ram[10600]), .I3(
        ram[10592]), .S0(n27049), .S1(n26574), .ZN(n21051) );
  MUX41 U10927 ( .I0(n21071), .I1(n21072), .I2(n21073), .I3(n21074), .S0(
        n26200), .S1(n26318), .ZN(n21070) );
  MUX41 U10928 ( .I0(ram[11032]), .I1(ram[11024]), .I2(ram[11016]), .I3(
        ram[11008]), .S0(n27050), .S1(n26575), .ZN(n21074) );
  MUX41 U10929 ( .I0(ram[11064]), .I1(ram[11056]), .I2(ram[11048]), .I3(
        ram[11040]), .S0(n27050), .S1(n26575), .ZN(n21072) );
  MUX41 U10930 ( .I0(ram[11128]), .I1(ram[11120]), .I2(ram[11112]), .I3(
        ram[11104]), .S0(n27050), .S1(n26575), .ZN(n21071) );
  MUX41 U10931 ( .I0(n21006), .I1(n21007), .I2(n21008), .I3(n21009), .S0(
        n26199), .S1(n26317), .ZN(n21005) );
  MUX41 U10932 ( .I0(ram[9528]), .I1(ram[9520]), .I2(ram[9512]), .I3(
        ram[9504]), .S0(n27046), .S1(n26571), .ZN(n21007) );
  MUX41 U10933 ( .I0(ram[9496]), .I1(ram[9488]), .I2(ram[9480]), .I3(
        ram[9472]), .S0(n27046), .S1(n26571), .ZN(n21009) );
  MUX41 U10934 ( .I0(ram[9592]), .I1(ram[9584]), .I2(ram[9576]), .I3(
        ram[9568]), .S0(n27046), .S1(n26571), .ZN(n21006) );
  MUX41 U10935 ( .I0(n21026), .I1(n21027), .I2(n21028), .I3(n21029), .S0(
        n26200), .S1(n26318), .ZN(n21025) );
  MUX41 U10936 ( .I0(ram[10040]), .I1(ram[10032]), .I2(ram[10024]), .I3(
        ram[10016]), .S0(n27048), .S1(n26573), .ZN(n21027) );
  MUX41 U10937 ( .I0(ram[10008]), .I1(ram[10000]), .I2(ram[9992]), .I3(
        ram[9984]), .S0(n27047), .S1(n26572), .ZN(n21029) );
  MUX41 U10938 ( .I0(ram[10104]), .I1(ram[10096]), .I2(ram[10088]), .I3(
        ram[10080]), .S0(n27048), .S1(n26573), .ZN(n21026) );
  MUX41 U10939 ( .I0(n20966), .I1(n20967), .I2(n20968), .I3(n20969), .S0(
        n26199), .S1(n26317), .ZN(n20965) );
  MUX41 U10940 ( .I0(ram[8504]), .I1(ram[8496]), .I2(ram[8488]), .I3(
        ram[8480]), .S0(n27044), .S1(n26569), .ZN(n20967) );
  MUX41 U10941 ( .I0(ram[8472]), .I1(ram[8464]), .I2(ram[8456]), .I3(
        ram[8448]), .S0(n27044), .S1(n26569), .ZN(n20969) );
  MUX41 U10942 ( .I0(ram[8568]), .I1(ram[8560]), .I2(ram[8552]), .I3(
        ram[8544]), .S0(n27044), .S1(n26569), .ZN(n20966) );
  MUX41 U10943 ( .I0(n20986), .I1(n20987), .I2(n20988), .I3(n20989), .S0(
        n26199), .S1(n26317), .ZN(n20985) );
  MUX41 U10944 ( .I0(ram[8984]), .I1(ram[8976]), .I2(ram[8968]), .I3(
        ram[8960]), .S0(n27045), .S1(n26570), .ZN(n20989) );
  MUX41 U10945 ( .I0(ram[9016]), .I1(ram[9008]), .I2(ram[9000]), .I3(
        ram[8992]), .S0(n27045), .S1(n26570), .ZN(n20987) );
  MUX41 U10946 ( .I0(ram[9080]), .I1(ram[9072]), .I2(ram[9064]), .I3(
        ram[9056]), .S0(n27045), .S1(n26570), .ZN(n20986) );
  MUX41 U10947 ( .I0(n21946), .I1(n21947), .I2(n21948), .I3(n21949), .S0(
        n26213), .S1(n26331), .ZN(n21945) );
  MUX41 U10948 ( .I0(ram[15641]), .I1(ram[15633]), .I2(ram[15625]), .I3(
        ram[15617]), .S0(n27100), .S1(n26625), .ZN(n21949) );
  MUX41 U10949 ( .I0(ram[15673]), .I1(ram[15665]), .I2(ram[15657]), .I3(
        ram[15649]), .S0(n27100), .S1(n26625), .ZN(n21947) );
  MUX41 U10950 ( .I0(ram[15737]), .I1(ram[15729]), .I2(ram[15721]), .I3(
        ram[15713]), .S0(n27101), .S1(n26626), .ZN(n21946) );
  MUX41 U10951 ( .I0(n21966), .I1(n21967), .I2(n21968), .I3(n21969), .S0(
        n26213), .S1(n26331), .ZN(n21965) );
  MUX41 U10952 ( .I0(ram[16153]), .I1(ram[16145]), .I2(ram[16137]), .I3(
        ram[16129]), .S0(n27102), .S1(n26627), .ZN(n21969) );
  MUX41 U10953 ( .I0(ram[16185]), .I1(ram[16177]), .I2(ram[16169]), .I3(
        ram[16161]), .S0(n27102), .S1(n26627), .ZN(n21967) );
  MUX41 U10954 ( .I0(ram[16249]), .I1(ram[16241]), .I2(ram[16233]), .I3(
        ram[16225]), .S0(n27102), .S1(n26627), .ZN(n21966) );
  MUX41 U10955 ( .I0(n21926), .I1(n21927), .I2(n21928), .I3(n21929), .S0(
        n26213), .S1(n26331), .ZN(n21925) );
  MUX41 U10956 ( .I0(ram[15129]), .I1(ram[15121]), .I2(ram[15113]), .I3(
        ram[15105]), .S0(n27099), .S1(n26624), .ZN(n21929) );
  MUX41 U10957 ( .I0(ram[15161]), .I1(ram[15153]), .I2(ram[15145]), .I3(
        ram[15137]), .S0(n27099), .S1(n26624), .ZN(n21927) );
  MUX41 U10958 ( .I0(ram[15225]), .I1(ram[15217]), .I2(ram[15209]), .I3(
        ram[15201]), .S0(n27099), .S1(n26624), .ZN(n21926) );
  MUX41 U10959 ( .I0(n21906), .I1(n21907), .I2(n21908), .I3(n21909), .S0(
        n26212), .S1(n26330), .ZN(n21905) );
  MUX41 U10960 ( .I0(ram[14617]), .I1(ram[14609]), .I2(ram[14601]), .I3(
        ram[14593]), .S0(n27098), .S1(n26623), .ZN(n21909) );
  MUX41 U10961 ( .I0(ram[14649]), .I1(ram[14641]), .I2(ram[14633]), .I3(
        ram[14625]), .S0(n27098), .S1(n26623), .ZN(n21907) );
  MUX41 U10962 ( .I0(ram[14713]), .I1(ram[14705]), .I2(ram[14697]), .I3(
        ram[14689]), .S0(n27098), .S1(n26623), .ZN(n21906) );
  MUX41 U10963 ( .I0(n21861), .I1(n21862), .I2(n21863), .I3(n21864), .S0(
        n26212), .S1(n26330), .ZN(n21860) );
  MUX41 U10964 ( .I0(ram[13593]), .I1(ram[13585]), .I2(ram[13577]), .I3(
        ram[13569]), .S0(n27095), .S1(n26620), .ZN(n21864) );
  MUX41 U10965 ( .I0(ram[13625]), .I1(ram[13617]), .I2(ram[13609]), .I3(
        ram[13601]), .S0(n27096), .S1(n26621), .ZN(n21862) );
  MUX41 U10966 ( .I0(ram[13689]), .I1(ram[13681]), .I2(ram[13673]), .I3(
        ram[13665]), .S0(n27096), .S1(n26621), .ZN(n21861) );
  MUX41 U10967 ( .I0(n21881), .I1(n21882), .I2(n21883), .I3(n21884), .S0(
        n26212), .S1(n26330), .ZN(n21880) );
  MUX41 U10968 ( .I0(ram[14105]), .I1(ram[14097]), .I2(ram[14089]), .I3(
        ram[14081]), .S0(n27097), .S1(n26622), .ZN(n21884) );
  MUX41 U10969 ( .I0(ram[14137]), .I1(ram[14129]), .I2(ram[14121]), .I3(
        ram[14113]), .S0(n27097), .S1(n26622), .ZN(n21882) );
  MUX41 U10970 ( .I0(ram[14201]), .I1(ram[14193]), .I2(ram[14185]), .I3(
        ram[14177]), .S0(n27097), .S1(n26622), .ZN(n21881) );
  MUX41 U10971 ( .I0(n21841), .I1(n21842), .I2(n21843), .I3(n21844), .S0(
        n26211), .S1(n26329), .ZN(n21840) );
  MUX41 U10972 ( .I0(ram[13081]), .I1(ram[13073]), .I2(ram[13065]), .I3(
        ram[13057]), .S0(n27094), .S1(n26619), .ZN(n21844) );
  MUX41 U10973 ( .I0(ram[13113]), .I1(ram[13105]), .I2(ram[13097]), .I3(
        ram[13089]), .S0(n27094), .S1(n26619), .ZN(n21842) );
  MUX41 U10974 ( .I0(ram[13177]), .I1(ram[13169]), .I2(ram[13161]), .I3(
        ram[13153]), .S0(n27094), .S1(n26619), .ZN(n21841) );
  MUX41 U10975 ( .I0(n21821), .I1(n21822), .I2(n21823), .I3(n21824), .S0(
        n26211), .S1(n26329), .ZN(n21820) );
  MUX41 U10976 ( .I0(ram[12569]), .I1(ram[12561]), .I2(ram[12553]), .I3(
        ram[12545]), .S0(n27093), .S1(n26618), .ZN(n21824) );
  MUX41 U10977 ( .I0(ram[12601]), .I1(ram[12593]), .I2(ram[12585]), .I3(
        ram[12577]), .S0(n27093), .S1(n26618), .ZN(n21822) );
  MUX41 U10978 ( .I0(ram[12665]), .I1(ram[12657]), .I2(ram[12649]), .I3(
        ram[12641]), .S0(n27093), .S1(n26618), .ZN(n21821) );
  MUX41 U10979 ( .I0(n21604), .I1(n21605), .I2(n21606), .I3(n21607), .S0(
        n26208), .S1(n26326), .ZN(n21603) );
  MUX41 U10980 ( .I0(ram[7481]), .I1(ram[7473]), .I2(ram[7465]), .I3(
        ram[7457]), .S0(n27081), .S1(n26606), .ZN(n21605) );
  MUX41 U10981 ( .I0(ram[7449]), .I1(ram[7441]), .I2(ram[7433]), .I3(
        ram[7425]), .S0(n27081), .S1(n26606), .ZN(n21607) );
  MUX41 U10982 ( .I0(ram[7545]), .I1(ram[7537]), .I2(ram[7529]), .I3(
        ram[7521]), .S0(n27081), .S1(n26606), .ZN(n21604) );
  MUX41 U10983 ( .I0(n21624), .I1(n21625), .I2(n21626), .I3(n21627), .S0(
        n26208), .S1(n26326), .ZN(n21623) );
  MUX41 U10984 ( .I0(ram[7961]), .I1(ram[7953]), .I2(ram[7945]), .I3(
        ram[7937]), .S0(n27082), .S1(n26607), .ZN(n21627) );
  MUX41 U10985 ( .I0(ram[7993]), .I1(ram[7985]), .I2(ram[7977]), .I3(
        ram[7969]), .S0(n27082), .S1(n26607), .ZN(n21625) );
  MUX41 U10986 ( .I0(ram[8057]), .I1(ram[8049]), .I2(ram[8041]), .I3(
        ram[8033]), .S0(n27082), .S1(n26607), .ZN(n21624) );
  MUX41 U10987 ( .I0(n21564), .I1(n21565), .I2(n21566), .I3(n21567), .S0(
        n26207), .S1(n26325), .ZN(n21563) );
  MUX41 U10988 ( .I0(ram[6425]), .I1(ram[6417]), .I2(ram[6409]), .I3(
        ram[6401]), .S0(n27078), .S1(n26603), .ZN(n21567) );
  MUX41 U10989 ( .I0(ram[6457]), .I1(ram[6449]), .I2(ram[6441]), .I3(
        ram[6433]), .S0(n27078), .S1(n26603), .ZN(n21565) );
  MUX41 U10990 ( .I0(ram[6521]), .I1(ram[6513]), .I2(ram[6505]), .I3(
        ram[6497]), .S0(n27078), .S1(n26603), .ZN(n21564) );
  MUX41 U10991 ( .I0(n21584), .I1(n21585), .I2(n21586), .I3(n21587), .S0(
        n26208), .S1(n26326), .ZN(n21583) );
  MUX41 U10992 ( .I0(ram[6937]), .I1(ram[6929]), .I2(ram[6921]), .I3(
        ram[6913]), .S0(n27079), .S1(n26604), .ZN(n21587) );
  MUX41 U10993 ( .I0(ram[6969]), .I1(ram[6961]), .I2(ram[6953]), .I3(
        ram[6945]), .S0(n27080), .S1(n26605), .ZN(n21585) );
  MUX41 U10994 ( .I0(ram[7033]), .I1(ram[7025]), .I2(ram[7017]), .I3(
        ram[7009]), .S0(n27080), .S1(n26605), .ZN(n21584) );
  MUX41 U10995 ( .I0(n21519), .I1(n21520), .I2(n21521), .I3(n21522), .S0(
        n26207), .S1(n26325), .ZN(n21518) );
  MUX41 U10996 ( .I0(ram[5433]), .I1(ram[5425]), .I2(ram[5417]), .I3(
        ram[5409]), .S0(n27076), .S1(n26601), .ZN(n21520) );
  MUX41 U10997 ( .I0(ram[5401]), .I1(ram[5393]), .I2(ram[5385]), .I3(
        ram[5377]), .S0(n27076), .S1(n26601), .ZN(n21522) );
  MUX41 U10998 ( .I0(ram[5497]), .I1(ram[5489]), .I2(ram[5481]), .I3(
        ram[5473]), .S0(n27076), .S1(n26601), .ZN(n21519) );
  MUX41 U10999 ( .I0(n21539), .I1(n21540), .I2(n21541), .I3(n21542), .S0(
        n26207), .S1(n26325), .ZN(n21538) );
  MUX41 U11000 ( .I0(ram[5945]), .I1(ram[5937]), .I2(ram[5929]), .I3(
        ram[5921]), .S0(n27077), .S1(n26602), .ZN(n21540) );
  MUX41 U11001 ( .I0(ram[5913]), .I1(ram[5905]), .I2(ram[5897]), .I3(
        ram[5889]), .S0(n27077), .S1(n26602), .ZN(n21542) );
  MUX41 U11002 ( .I0(ram[6009]), .I1(ram[6001]), .I2(ram[5993]), .I3(
        ram[5985]), .S0(n27077), .S1(n26602), .ZN(n21539) );
  MUX41 U11003 ( .I0(n21479), .I1(n21480), .I2(n21481), .I3(n21482), .S0(
        n26206), .S1(n26324), .ZN(n21478) );
  MUX41 U11004 ( .I0(ram[4409]), .I1(ram[4401]), .I2(ram[4393]), .I3(
        ram[4385]), .S0(n27073), .S1(n26598), .ZN(n21480) );
  MUX41 U11005 ( .I0(ram[4377]), .I1(ram[4369]), .I2(ram[4361]), .I3(
        ram[4353]), .S0(n27073), .S1(n26598), .ZN(n21482) );
  MUX41 U11006 ( .I0(ram[4473]), .I1(ram[4465]), .I2(ram[4457]), .I3(
        ram[4449]), .S0(n27074), .S1(n26599), .ZN(n21479) );
  MUX41 U11007 ( .I0(n21499), .I1(n21500), .I2(n21501), .I3(n21502), .S0(
        n26207), .S1(n26325), .ZN(n21498) );
  MUX41 U11008 ( .I0(ram[4889]), .I1(ram[4881]), .I2(ram[4873]), .I3(
        ram[4865]), .S0(n27075), .S1(n26600), .ZN(n21502) );
  MUX41 U11009 ( .I0(ram[4921]), .I1(ram[4913]), .I2(ram[4905]), .I3(
        ram[4897]), .S0(n27075), .S1(n26600), .ZN(n21500) );
  MUX41 U11010 ( .I0(ram[4985]), .I1(ram[4977]), .I2(ram[4969]), .I3(
        ram[4961]), .S0(n27075), .S1(n26600), .ZN(n21499) );
  MUX41 U11011 ( .I0(n21775), .I1(n21776), .I2(n21777), .I3(n21778), .S0(
        n26211), .S1(n26329), .ZN(n21774) );
  MUX41 U11012 ( .I0(ram[11577]), .I1(ram[11569]), .I2(ram[11561]), .I3(
        ram[11553]), .S0(n27091), .S1(n26616), .ZN(n21776) );
  MUX41 U11013 ( .I0(ram[11545]), .I1(ram[11537]), .I2(ram[11529]), .I3(
        ram[11521]), .S0(n27091), .S1(n26616), .ZN(n21778) );
  MUX41 U11014 ( .I0(ram[11641]), .I1(ram[11633]), .I2(ram[11625]), .I3(
        ram[11617]), .S0(n27091), .S1(n26616), .ZN(n21775) );
  MUX41 U11015 ( .I0(n21795), .I1(n21796), .I2(n21797), .I3(n21798), .S0(
        n26211), .S1(n26329), .ZN(n21794) );
  MUX41 U11016 ( .I0(ram[12089]), .I1(ram[12081]), .I2(ram[12073]), .I3(
        ram[12065]), .S0(n27092), .S1(n26617), .ZN(n21796) );
  MUX41 U11017 ( .I0(ram[12057]), .I1(ram[12049]), .I2(ram[12041]), .I3(
        ram[12033]), .S0(n27092), .S1(n26617), .ZN(n21798) );
  MUX41 U11018 ( .I0(ram[12153]), .I1(ram[12145]), .I2(ram[12137]), .I3(
        ram[12129]), .S0(n27092), .S1(n26617), .ZN(n21795) );
  MUX41 U11019 ( .I0(n21735), .I1(n21736), .I2(n21737), .I3(n21738), .S0(
        n26210), .S1(n26328), .ZN(n21734) );
  MUX41 U11020 ( .I0(ram[10553]), .I1(ram[10545]), .I2(ram[10537]), .I3(
        ram[10529]), .S0(n27088), .S1(n26613), .ZN(n21736) );
  MUX41 U11021 ( .I0(ram[10521]), .I1(ram[10513]), .I2(ram[10505]), .I3(
        ram[10497]), .S0(n27088), .S1(n26613), .ZN(n21738) );
  MUX41 U11022 ( .I0(ram[10617]), .I1(ram[10609]), .I2(ram[10601]), .I3(
        ram[10593]), .S0(n27088), .S1(n26613), .ZN(n21735) );
  MUX41 U11023 ( .I0(n21755), .I1(n21756), .I2(n21757), .I3(n21758), .S0(
        n26210), .S1(n26328), .ZN(n21754) );
  MUX41 U11024 ( .I0(ram[11033]), .I1(ram[11025]), .I2(ram[11017]), .I3(
        ram[11009]), .S0(n27089), .S1(n26614), .ZN(n21758) );
  MUX41 U11025 ( .I0(ram[11065]), .I1(ram[11057]), .I2(ram[11049]), .I3(
        ram[11041]), .S0(n27089), .S1(n26614), .ZN(n21756) );
  MUX41 U11026 ( .I0(ram[11129]), .I1(ram[11121]), .I2(ram[11113]), .I3(
        ram[11105]), .S0(n27090), .S1(n26615), .ZN(n21755) );
  MUX41 U11027 ( .I0(n21690), .I1(n21691), .I2(n21692), .I3(n21693), .S0(
        n26209), .S1(n26327), .ZN(n21689) );
  MUX41 U11028 ( .I0(ram[9529]), .I1(ram[9521]), .I2(ram[9513]), .I3(
        ram[9505]), .S0(n27086), .S1(n26611), .ZN(n21691) );
  MUX41 U11029 ( .I0(ram[9497]), .I1(ram[9489]), .I2(ram[9481]), .I3(
        ram[9473]), .S0(n27086), .S1(n26611), .ZN(n21693) );
  MUX41 U11030 ( .I0(ram[9593]), .I1(ram[9585]), .I2(ram[9577]), .I3(
        ram[9569]), .S0(n27086), .S1(n26611), .ZN(n21690) );
  MUX41 U11031 ( .I0(n21710), .I1(n21711), .I2(n21712), .I3(n21713), .S0(
        n26210), .S1(n26328), .ZN(n21709) );
  MUX41 U11032 ( .I0(ram[10041]), .I1(ram[10033]), .I2(ram[10025]), .I3(
        ram[10017]), .S0(n27087), .S1(n26612), .ZN(n21711) );
  MUX41 U11033 ( .I0(ram[10009]), .I1(ram[10001]), .I2(ram[9993]), .I3(
        ram[9985]), .S0(n27087), .S1(n26612), .ZN(n21713) );
  MUX41 U11034 ( .I0(ram[10105]), .I1(ram[10097]), .I2(ram[10089]), .I3(
        ram[10081]), .S0(n27087), .S1(n26612), .ZN(n21710) );
  MUX41 U11035 ( .I0(n21650), .I1(n21651), .I2(n21652), .I3(n21653), .S0(
        n26209), .S1(n26327), .ZN(n21649) );
  MUX41 U11036 ( .I0(ram[8505]), .I1(ram[8497]), .I2(ram[8489]), .I3(
        ram[8481]), .S0(n27083), .S1(n26608), .ZN(n21651) );
  MUX41 U11037 ( .I0(ram[8473]), .I1(ram[8465]), .I2(ram[8457]), .I3(
        ram[8449]), .S0(n27083), .S1(n26608), .ZN(n21653) );
  MUX41 U11038 ( .I0(ram[8569]), .I1(ram[8561]), .I2(ram[8553]), .I3(
        ram[8545]), .S0(n27083), .S1(n26608), .ZN(n21650) );
  MUX41 U11039 ( .I0(n21670), .I1(n21671), .I2(n21672), .I3(n21673), .S0(
        n26209), .S1(n26327), .ZN(n21669) );
  MUX41 U11040 ( .I0(ram[8985]), .I1(ram[8977]), .I2(ram[8969]), .I3(
        ram[8961]), .S0(n27084), .S1(n26609), .ZN(n21673) );
  MUX41 U11041 ( .I0(ram[9017]), .I1(ram[9009]), .I2(ram[9001]), .I3(
        ram[8993]), .S0(n27084), .S1(n26609), .ZN(n21671) );
  MUX41 U11042 ( .I0(ram[9081]), .I1(ram[9073]), .I2(ram[9065]), .I3(
        ram[9057]), .S0(n27085), .S1(n26610), .ZN(n21670) );
  MUX41 U11043 ( .I0(n22630), .I1(n22631), .I2(n22632), .I3(n22633), .S0(
        n26223), .S1(n26341), .ZN(n22629) );
  MUX41 U11044 ( .I0(ram[15642]), .I1(ram[15634]), .I2(ram[15626]), .I3(
        ram[15618]), .S0(n27140), .S1(n26665), .ZN(n22633) );
  MUX41 U11045 ( .I0(ram[15674]), .I1(ram[15666]), .I2(ram[15658]), .I3(
        ram[15650]), .S0(n27140), .S1(n26665), .ZN(n22631) );
  MUX41 U11046 ( .I0(ram[15738]), .I1(ram[15730]), .I2(ram[15722]), .I3(
        ram[15714]), .S0(n27140), .S1(n26665), .ZN(n22630) );
  MUX41 U11047 ( .I0(n22650), .I1(n22651), .I2(n22652), .I3(n22653), .S0(
        n26223), .S1(n26341), .ZN(n22649) );
  MUX41 U11048 ( .I0(ram[16154]), .I1(ram[16146]), .I2(ram[16138]), .I3(
        ram[16130]), .S0(n27141), .S1(n26666), .ZN(n22653) );
  MUX41 U11049 ( .I0(ram[16186]), .I1(ram[16178]), .I2(ram[16170]), .I3(
        ram[16162]), .S0(n27141), .S1(n26666), .ZN(n22651) );
  MUX41 U11050 ( .I0(ram[16250]), .I1(ram[16242]), .I2(ram[16234]), .I3(
        ram[16226]), .S0(n27141), .S1(n26666), .ZN(n22650) );
  MUX41 U11051 ( .I0(n22610), .I1(n22611), .I2(n22612), .I3(n22613), .S0(
        n26223), .S1(n26341), .ZN(n22609) );
  MUX41 U11052 ( .I0(ram[15130]), .I1(ram[15122]), .I2(ram[15114]), .I3(
        ram[15106]), .S0(n27139), .S1(n26664), .ZN(n22613) );
  MUX41 U11053 ( .I0(ram[15162]), .I1(ram[15154]), .I2(ram[15146]), .I3(
        ram[15138]), .S0(n27139), .S1(n26664), .ZN(n22611) );
  MUX41 U11054 ( .I0(ram[15226]), .I1(ram[15218]), .I2(ram[15210]), .I3(
        ram[15202]), .S0(n27139), .S1(n26664), .ZN(n22610) );
  MUX41 U11055 ( .I0(n22590), .I1(n22591), .I2(n22592), .I3(n22593), .S0(
        n26222), .S1(n26340), .ZN(n22589) );
  MUX41 U11056 ( .I0(ram[14618]), .I1(ram[14610]), .I2(ram[14602]), .I3(
        ram[14594]), .S0(n27137), .S1(n26662), .ZN(n22593) );
  MUX41 U11057 ( .I0(ram[14650]), .I1(ram[14642]), .I2(ram[14634]), .I3(
        ram[14626]), .S0(n27137), .S1(n26662), .ZN(n22591) );
  MUX41 U11058 ( .I0(ram[14714]), .I1(ram[14706]), .I2(ram[14698]), .I3(
        ram[14690]), .S0(n27138), .S1(n26663), .ZN(n22590) );
  MUX41 U11059 ( .I0(n22545), .I1(n22546), .I2(n22547), .I3(n22548), .S0(
        n26222), .S1(n26340), .ZN(n22544) );
  MUX41 U11060 ( .I0(ram[13594]), .I1(ram[13586]), .I2(ram[13578]), .I3(
        ram[13570]), .S0(n27135), .S1(n26660), .ZN(n22548) );
  MUX41 U11061 ( .I0(ram[13626]), .I1(ram[13618]), .I2(ram[13610]), .I3(
        ram[13602]), .S0(n27135), .S1(n26660), .ZN(n22546) );
  MUX41 U11062 ( .I0(ram[13690]), .I1(ram[13682]), .I2(ram[13674]), .I3(
        ram[13666]), .S0(n27135), .S1(n26660), .ZN(n22545) );
  MUX41 U11063 ( .I0(n22565), .I1(n22566), .I2(n22567), .I3(n22568), .S0(
        n26222), .S1(n26340), .ZN(n22564) );
  MUX41 U11064 ( .I0(ram[14106]), .I1(ram[14098]), .I2(ram[14090]), .I3(
        ram[14082]), .S0(n27136), .S1(n26661), .ZN(n22568) );
  MUX41 U11065 ( .I0(ram[14138]), .I1(ram[14130]), .I2(ram[14122]), .I3(
        ram[14114]), .S0(n27136), .S1(n26661), .ZN(n22566) );
  MUX41 U11066 ( .I0(ram[14202]), .I1(ram[14194]), .I2(ram[14186]), .I3(
        ram[14178]), .S0(n27136), .S1(n26661), .ZN(n22565) );
  MUX41 U11067 ( .I0(n22525), .I1(n22526), .I2(n22527), .I3(n22528), .S0(
        n26221), .S1(n26339), .ZN(n22524) );
  MUX41 U11068 ( .I0(ram[13082]), .I1(ram[13074]), .I2(ram[13066]), .I3(
        ram[13058]), .S0(n27134), .S1(n26659), .ZN(n22528) );
  MUX41 U11069 ( .I0(ram[13114]), .I1(ram[13106]), .I2(ram[13098]), .I3(
        ram[13090]), .S0(n27134), .S1(n26659), .ZN(n22526) );
  MUX41 U11070 ( .I0(ram[13178]), .I1(ram[13170]), .I2(ram[13162]), .I3(
        ram[13154]), .S0(n27134), .S1(n26659), .ZN(n22525) );
  MUX41 U11071 ( .I0(n22505), .I1(n22506), .I2(n22507), .I3(n22508), .S0(
        n26221), .S1(n26339), .ZN(n22504) );
  MUX41 U11072 ( .I0(ram[12570]), .I1(ram[12562]), .I2(ram[12554]), .I3(
        ram[12546]), .S0(n27132), .S1(n26657), .ZN(n22508) );
  MUX41 U11073 ( .I0(ram[12602]), .I1(ram[12594]), .I2(ram[12586]), .I3(
        ram[12578]), .S0(n27132), .S1(n26657), .ZN(n22506) );
  MUX41 U11074 ( .I0(ram[12666]), .I1(ram[12658]), .I2(ram[12650]), .I3(
        ram[12642]), .S0(n27133), .S1(n26658), .ZN(n22505) );
  MUX41 U11075 ( .I0(n22288), .I1(n22289), .I2(n22290), .I3(n22291), .S0(
        n26218), .S1(n26336), .ZN(n22287) );
  MUX41 U11076 ( .I0(ram[7482]), .I1(ram[7474]), .I2(ram[7466]), .I3(
        ram[7458]), .S0(n27120), .S1(n26645), .ZN(n22289) );
  MUX41 U11077 ( .I0(ram[7450]), .I1(ram[7442]), .I2(ram[7434]), .I3(
        ram[7426]), .S0(n27120), .S1(n26645), .ZN(n22291) );
  MUX41 U11078 ( .I0(ram[7546]), .I1(ram[7538]), .I2(ram[7530]), .I3(
        ram[7522]), .S0(n27120), .S1(n26645), .ZN(n22288) );
  MUX41 U11079 ( .I0(n22308), .I1(n22309), .I2(n22310), .I3(n22311), .S0(
        n26218), .S1(n26336), .ZN(n22307) );
  MUX41 U11080 ( .I0(ram[7962]), .I1(ram[7954]), .I2(ram[7946]), .I3(
        ram[7938]), .S0(n27121), .S1(n26646), .ZN(n22311) );
  MUX41 U11081 ( .I0(ram[7994]), .I1(ram[7986]), .I2(ram[7978]), .I3(
        ram[7970]), .S0(n27121), .S1(n26646), .ZN(n22309) );
  MUX41 U11082 ( .I0(ram[8058]), .I1(ram[8050]), .I2(ram[8042]), .I3(
        ram[8034]), .S0(n27122), .S1(n26647), .ZN(n22308) );
  MUX41 U11083 ( .I0(n22248), .I1(n22249), .I2(n22250), .I3(n22251), .S0(
        n26217), .S1(n26335), .ZN(n22247) );
  MUX41 U11084 ( .I0(ram[6426]), .I1(ram[6418]), .I2(ram[6410]), .I3(
        ram[6402]), .S0(n27118), .S1(n26643), .ZN(n22251) );
  MUX41 U11085 ( .I0(ram[6458]), .I1(ram[6450]), .I2(ram[6442]), .I3(
        ram[6434]), .S0(n27118), .S1(n26643), .ZN(n22249) );
  MUX41 U11086 ( .I0(ram[6522]), .I1(ram[6514]), .I2(ram[6506]), .I3(
        ram[6498]), .S0(n27118), .S1(n26643), .ZN(n22248) );
  MUX41 U11087 ( .I0(n22268), .I1(n22269), .I2(n22270), .I3(n22271), .S0(
        n26218), .S1(n26336), .ZN(n22267) );
  MUX41 U11088 ( .I0(ram[6938]), .I1(ram[6930]), .I2(ram[6922]), .I3(
        ram[6914]), .S0(n27119), .S1(n26644), .ZN(n22271) );
  MUX41 U11089 ( .I0(ram[6970]), .I1(ram[6962]), .I2(ram[6954]), .I3(
        ram[6946]), .S0(n27119), .S1(n26644), .ZN(n22269) );
  MUX41 U11090 ( .I0(ram[7034]), .I1(ram[7026]), .I2(ram[7018]), .I3(
        ram[7010]), .S0(n27119), .S1(n26644), .ZN(n22268) );
  MUX41 U11091 ( .I0(n22203), .I1(n22204), .I2(n22205), .I3(n22206), .S0(
        n26217), .S1(n26335), .ZN(n22202) );
  MUX41 U11092 ( .I0(ram[5434]), .I1(ram[5426]), .I2(ram[5418]), .I3(
        ram[5410]), .S0(n27115), .S1(n26640), .ZN(n22204) );
  MUX41 U11093 ( .I0(ram[5402]), .I1(ram[5394]), .I2(ram[5386]), .I3(
        ram[5378]), .S0(n27115), .S1(n26640), .ZN(n22206) );
  MUX41 U11094 ( .I0(ram[5498]), .I1(ram[5490]), .I2(ram[5482]), .I3(
        ram[5474]), .S0(n27115), .S1(n26640), .ZN(n22203) );
  MUX41 U11095 ( .I0(n22223), .I1(n22224), .I2(n22225), .I3(n22226), .S0(
        n26217), .S1(n26335), .ZN(n22222) );
  MUX41 U11096 ( .I0(ram[5946]), .I1(ram[5938]), .I2(ram[5930]), .I3(
        ram[5922]), .S0(n27116), .S1(n26641), .ZN(n22224) );
  MUX41 U11097 ( .I0(ram[5914]), .I1(ram[5906]), .I2(ram[5898]), .I3(
        ram[5890]), .S0(n27116), .S1(n26641), .ZN(n22226) );
  MUX41 U11098 ( .I0(ram[6010]), .I1(ram[6002]), .I2(ram[5994]), .I3(
        ram[5986]), .S0(n27117), .S1(n26642), .ZN(n22223) );
  MUX41 U11099 ( .I0(n22163), .I1(n22164), .I2(n22165), .I3(n22166), .S0(
        n26216), .S1(n26334), .ZN(n22162) );
  MUX41 U11100 ( .I0(ram[4410]), .I1(ram[4402]), .I2(ram[4394]), .I3(
        ram[4386]), .S0(n27113), .S1(n26638), .ZN(n22164) );
  MUX41 U11101 ( .I0(ram[4378]), .I1(ram[4370]), .I2(ram[4362]), .I3(
        ram[4354]), .S0(n27113), .S1(n26638), .ZN(n22166) );
  MUX41 U11102 ( .I0(ram[4474]), .I1(ram[4466]), .I2(ram[4458]), .I3(
        ram[4450]), .S0(n27113), .S1(n26638), .ZN(n22163) );
  MUX41 U11103 ( .I0(n22183), .I1(n22184), .I2(n22185), .I3(n22186), .S0(
        n26216), .S1(n26334), .ZN(n22182) );
  MUX41 U11104 ( .I0(ram[4890]), .I1(ram[4882]), .I2(ram[4874]), .I3(
        ram[4866]), .S0(n27114), .S1(n26639), .ZN(n22186) );
  MUX41 U11105 ( .I0(ram[4922]), .I1(ram[4914]), .I2(ram[4906]), .I3(
        ram[4898]), .S0(n27114), .S1(n26639), .ZN(n22184) );
  MUX41 U11106 ( .I0(ram[4986]), .I1(ram[4978]), .I2(ram[4970]), .I3(
        ram[4962]), .S0(n27114), .S1(n26639), .ZN(n22183) );
  MUX41 U11107 ( .I0(n22459), .I1(n22460), .I2(n22461), .I3(n22462), .S0(
        n26220), .S1(n26338), .ZN(n22458) );
  MUX41 U11108 ( .I0(ram[11578]), .I1(ram[11570]), .I2(ram[11562]), .I3(
        ram[11554]), .S0(n27130), .S1(n26655), .ZN(n22460) );
  MUX41 U11109 ( .I0(ram[11546]), .I1(ram[11538]), .I2(ram[11530]), .I3(
        ram[11522]), .S0(n27130), .S1(n26655), .ZN(n22462) );
  MUX41 U11110 ( .I0(ram[11642]), .I1(ram[11634]), .I2(ram[11626]), .I3(
        ram[11618]), .S0(n27130), .S1(n26655), .ZN(n22459) );
  MUX41 U11111 ( .I0(n22479), .I1(n22480), .I2(n22481), .I3(n22482), .S0(
        n26221), .S1(n26339), .ZN(n22478) );
  MUX41 U11112 ( .I0(ram[12090]), .I1(ram[12082]), .I2(ram[12074]), .I3(
        ram[12066]), .S0(n27131), .S1(n26656), .ZN(n22480) );
  MUX41 U11113 ( .I0(ram[12058]), .I1(ram[12050]), .I2(ram[12042]), .I3(
        ram[12034]), .S0(n27131), .S1(n26656), .ZN(n22482) );
  MUX41 U11114 ( .I0(ram[12154]), .I1(ram[12146]), .I2(ram[12138]), .I3(
        ram[12130]), .S0(n27131), .S1(n26656), .ZN(n22479) );
  MUX41 U11115 ( .I0(n22419), .I1(n22420), .I2(n22421), .I3(n22422), .S0(
        n26220), .S1(n26338), .ZN(n22418) );
  MUX41 U11116 ( .I0(ram[10554]), .I1(ram[10546]), .I2(ram[10538]), .I3(
        ram[10530]), .S0(n27128), .S1(n26653), .ZN(n22420) );
  MUX41 U11117 ( .I0(ram[10522]), .I1(ram[10514]), .I2(ram[10506]), .I3(
        ram[10498]), .S0(n27127), .S1(n26652), .ZN(n22422) );
  MUX41 U11118 ( .I0(ram[10618]), .I1(ram[10610]), .I2(ram[10602]), .I3(
        ram[10594]), .S0(n27128), .S1(n26653), .ZN(n22419) );
  MUX41 U11119 ( .I0(n22439), .I1(n22440), .I2(n22441), .I3(n22442), .S0(
        n26220), .S1(n26338), .ZN(n22438) );
  MUX41 U11120 ( .I0(ram[11034]), .I1(ram[11026]), .I2(ram[11018]), .I3(
        ram[11010]), .S0(n27129), .S1(n26654), .ZN(n22442) );
  MUX41 U11121 ( .I0(ram[11066]), .I1(ram[11058]), .I2(ram[11050]), .I3(
        ram[11042]), .S0(n27129), .S1(n26654), .ZN(n22440) );
  MUX41 U11122 ( .I0(ram[11130]), .I1(ram[11122]), .I2(ram[11114]), .I3(
        ram[11106]), .S0(n27129), .S1(n26654), .ZN(n22439) );
  MUX41 U11123 ( .I0(n22374), .I1(n22375), .I2(n22376), .I3(n22377), .S0(
        n26219), .S1(n26337), .ZN(n22373) );
  MUX41 U11124 ( .I0(ram[9530]), .I1(ram[9522]), .I2(ram[9514]), .I3(
        ram[9506]), .S0(n27125), .S1(n26650), .ZN(n22375) );
  MUX41 U11125 ( .I0(ram[9498]), .I1(ram[9490]), .I2(ram[9482]), .I3(
        ram[9474]), .S0(n27125), .S1(n26650), .ZN(n22377) );
  MUX41 U11126 ( .I0(ram[9594]), .I1(ram[9586]), .I2(ram[9578]), .I3(
        ram[9570]), .S0(n27125), .S1(n26650), .ZN(n22374) );
  MUX41 U11127 ( .I0(n22394), .I1(n22395), .I2(n22396), .I3(n22397), .S0(
        n26219), .S1(n26337), .ZN(n22393) );
  MUX41 U11128 ( .I0(ram[10042]), .I1(ram[10034]), .I2(ram[10026]), .I3(
        ram[10018]), .S0(n27126), .S1(n26651), .ZN(n22395) );
  MUX41 U11129 ( .I0(ram[10010]), .I1(ram[10002]), .I2(ram[9994]), .I3(
        ram[9986]), .S0(n27126), .S1(n26651), .ZN(n22397) );
  MUX41 U11130 ( .I0(ram[10106]), .I1(ram[10098]), .I2(ram[10090]), .I3(
        ram[10082]), .S0(n27126), .S1(n26651), .ZN(n22394) );
  MUX41 U11131 ( .I0(n22334), .I1(n22335), .I2(n22336), .I3(n22337), .S0(
        n26219), .S1(n26337), .ZN(n22333) );
  MUX41 U11132 ( .I0(ram[8506]), .I1(ram[8498]), .I2(ram[8490]), .I3(
        ram[8482]), .S0(n27123), .S1(n26648), .ZN(n22335) );
  MUX41 U11133 ( .I0(ram[8474]), .I1(ram[8466]), .I2(ram[8458]), .I3(
        ram[8450]), .S0(n27123), .S1(n26648), .ZN(n22337) );
  MUX41 U11134 ( .I0(ram[8570]), .I1(ram[8562]), .I2(ram[8554]), .I3(
        ram[8546]), .S0(n27123), .S1(n26648), .ZN(n22334) );
  MUX41 U11135 ( .I0(n22354), .I1(n22355), .I2(n22356), .I3(n22357), .S0(
        n26219), .S1(n26337), .ZN(n22353) );
  MUX41 U11136 ( .I0(ram[8986]), .I1(ram[8978]), .I2(ram[8970]), .I3(
        ram[8962]), .S0(n27124), .S1(n26649), .ZN(n22357) );
  MUX41 U11137 ( .I0(ram[9018]), .I1(ram[9010]), .I2(ram[9002]), .I3(
        ram[8994]), .S0(n27124), .S1(n26649), .ZN(n22355) );
  MUX41 U11138 ( .I0(ram[9082]), .I1(ram[9074]), .I2(ram[9066]), .I3(
        ram[9058]), .S0(n27124), .S1(n26649), .ZN(n22354) );
  MUX41 U11139 ( .I0(n23314), .I1(n23315), .I2(n23316), .I3(n23317), .S0(
        n26233), .S1(n26351), .ZN(n23313) );
  MUX41 U11140 ( .I0(ram[15643]), .I1(ram[15635]), .I2(ram[15627]), .I3(
        ram[15619]), .S0(n27179), .S1(n26704), .ZN(n23317) );
  MUX41 U11141 ( .I0(ram[15675]), .I1(ram[15667]), .I2(ram[15659]), .I3(
        ram[15651]), .S0(n27179), .S1(n26704), .ZN(n23315) );
  MUX41 U11142 ( .I0(ram[15739]), .I1(ram[15731]), .I2(ram[15723]), .I3(
        ram[15715]), .S0(n27179), .S1(n26704), .ZN(n23314) );
  MUX41 U11143 ( .I0(n23334), .I1(n23335), .I2(n23336), .I3(n23337), .S0(
        n26233), .S1(n26351), .ZN(n23333) );
  MUX41 U11144 ( .I0(ram[16155]), .I1(ram[16147]), .I2(ram[16139]), .I3(
        ram[16131]), .S0(n27180), .S1(n26705), .ZN(n23337) );
  MUX41 U11145 ( .I0(ram[16187]), .I1(ram[16179]), .I2(ram[16171]), .I3(
        ram[16163]), .S0(n27180), .S1(n26705), .ZN(n23335) );
  MUX41 U11146 ( .I0(ram[16251]), .I1(ram[16243]), .I2(ram[16235]), .I3(
        ram[16227]), .S0(n27181), .S1(n26706), .ZN(n23334) );
  MUX41 U11147 ( .I0(n23294), .I1(n23295), .I2(n23296), .I3(n23297), .S0(
        n26232), .S1(n26350), .ZN(n23293) );
  MUX41 U11148 ( .I0(ram[15131]), .I1(ram[15123]), .I2(ram[15115]), .I3(
        ram[15107]), .S0(n27178), .S1(n26703), .ZN(n23297) );
  MUX41 U11149 ( .I0(ram[15163]), .I1(ram[15155]), .I2(ram[15147]), .I3(
        ram[15139]), .S0(n27178), .S1(n26703), .ZN(n23295) );
  MUX41 U11150 ( .I0(ram[15227]), .I1(ram[15219]), .I2(ram[15211]), .I3(
        ram[15203]), .S0(n27178), .S1(n26703), .ZN(n23294) );
  MUX41 U11151 ( .I0(n23274), .I1(n23275), .I2(n23276), .I3(n23277), .S0(
        n26232), .S1(n26350), .ZN(n23273) );
  MUX41 U11152 ( .I0(ram[14619]), .I1(ram[14611]), .I2(ram[14603]), .I3(
        ram[14595]), .S0(n27177), .S1(n26702), .ZN(n23277) );
  MUX41 U11153 ( .I0(ram[14651]), .I1(ram[14643]), .I2(ram[14635]), .I3(
        ram[14627]), .S0(n27177), .S1(n26702), .ZN(n23275) );
  MUX41 U11154 ( .I0(ram[14715]), .I1(ram[14707]), .I2(ram[14699]), .I3(
        ram[14691]), .S0(n27177), .S1(n26702), .ZN(n23274) );
  MUX41 U11155 ( .I0(n23229), .I1(n23230), .I2(n23231), .I3(n23232), .S0(
        n26231), .S1(n26349), .ZN(n23228) );
  MUX41 U11156 ( .I0(ram[13595]), .I1(ram[13587]), .I2(ram[13579]), .I3(
        ram[13571]), .S0(n27174), .S1(n26699), .ZN(n23232) );
  MUX41 U11157 ( .I0(ram[13627]), .I1(ram[13619]), .I2(ram[13611]), .I3(
        ram[13603]), .S0(n27174), .S1(n26699), .ZN(n23230) );
  MUX41 U11158 ( .I0(ram[13691]), .I1(ram[13683]), .I2(ram[13675]), .I3(
        ram[13667]), .S0(n27174), .S1(n26699), .ZN(n23229) );
  MUX41 U11159 ( .I0(n23249), .I1(n23250), .I2(n23251), .I3(n23252), .S0(
        n26232), .S1(n26350), .ZN(n23248) );
  MUX41 U11160 ( .I0(ram[14107]), .I1(ram[14099]), .I2(ram[14091]), .I3(
        ram[14083]), .S0(n27175), .S1(n26700), .ZN(n23252) );
  MUX41 U11161 ( .I0(ram[14139]), .I1(ram[14131]), .I2(ram[14123]), .I3(
        ram[14115]), .S0(n27176), .S1(n26701), .ZN(n23250) );
  MUX41 U11162 ( .I0(ram[14203]), .I1(ram[14195]), .I2(ram[14187]), .I3(
        ram[14179]), .S0(n27176), .S1(n26701), .ZN(n23249) );
  MUX41 U11163 ( .I0(n23209), .I1(n23210), .I2(n23211), .I3(n23212), .S0(
        n26231), .S1(n26349), .ZN(n23208) );
  MUX41 U11164 ( .I0(ram[13083]), .I1(ram[13075]), .I2(ram[13067]), .I3(
        ram[13059]), .S0(n27173), .S1(n26698), .ZN(n23212) );
  MUX41 U11165 ( .I0(ram[13115]), .I1(ram[13107]), .I2(ram[13099]), .I3(
        ram[13091]), .S0(n27173), .S1(n26698), .ZN(n23210) );
  MUX41 U11166 ( .I0(ram[13179]), .I1(ram[13171]), .I2(ram[13163]), .I3(
        ram[13155]), .S0(n27173), .S1(n26698), .ZN(n23209) );
  MUX41 U11167 ( .I0(n23189), .I1(n23190), .I2(n23191), .I3(n23192), .S0(
        n26231), .S1(n26349), .ZN(n23188) );
  MUX41 U11168 ( .I0(ram[12571]), .I1(ram[12563]), .I2(ram[12555]), .I3(
        ram[12547]), .S0(n27172), .S1(n26697), .ZN(n23192) );
  MUX41 U11169 ( .I0(ram[12603]), .I1(ram[12595]), .I2(ram[12587]), .I3(
        ram[12579]), .S0(n27172), .S1(n26697), .ZN(n23190) );
  MUX41 U11170 ( .I0(ram[12667]), .I1(ram[12659]), .I2(ram[12651]), .I3(
        ram[12643]), .S0(n27172), .S1(n26697), .ZN(n23189) );
  MUX41 U11171 ( .I0(n22972), .I1(n22973), .I2(n22974), .I3(n22975), .S0(
        n26228), .S1(n26346), .ZN(n22971) );
  MUX41 U11172 ( .I0(ram[7483]), .I1(ram[7475]), .I2(ram[7467]), .I3(
        ram[7459]), .S0(n27160), .S1(n26685), .ZN(n22973) );
  MUX41 U11173 ( .I0(ram[7451]), .I1(ram[7443]), .I2(ram[7435]), .I3(
        ram[7427]), .S0(n27159), .S1(n26684), .ZN(n22975) );
  MUX41 U11174 ( .I0(ram[7547]), .I1(ram[7539]), .I2(ram[7531]), .I3(
        ram[7523]), .S0(n27160), .S1(n26685), .ZN(n22972) );
  MUX41 U11175 ( .I0(n22992), .I1(n22993), .I2(n22994), .I3(n22995), .S0(
        n26228), .S1(n26346), .ZN(n22991) );
  MUX41 U11176 ( .I0(ram[7963]), .I1(ram[7955]), .I2(ram[7947]), .I3(
        ram[7939]), .S0(n27161), .S1(n26686), .ZN(n22995) );
  MUX41 U11177 ( .I0(ram[7995]), .I1(ram[7987]), .I2(ram[7979]), .I3(
        ram[7971]), .S0(n27161), .S1(n26686), .ZN(n22993) );
  MUX41 U11178 ( .I0(ram[8059]), .I1(ram[8051]), .I2(ram[8043]), .I3(
        ram[8035]), .S0(n27161), .S1(n26686), .ZN(n22992) );
  MUX41 U11179 ( .I0(n22932), .I1(n22933), .I2(n22934), .I3(n22935), .S0(
        n26227), .S1(n26345), .ZN(n22931) );
  MUX41 U11180 ( .I0(ram[6427]), .I1(ram[6419]), .I2(ram[6411]), .I3(
        ram[6403]), .S0(n27157), .S1(n26682), .ZN(n22935) );
  MUX41 U11181 ( .I0(ram[6459]), .I1(ram[6451]), .I2(ram[6443]), .I3(
        ram[6435]), .S0(n27157), .S1(n26682), .ZN(n22933) );
  MUX41 U11182 ( .I0(ram[6523]), .I1(ram[6515]), .I2(ram[6507]), .I3(
        ram[6499]), .S0(n27157), .S1(n26682), .ZN(n22932) );
  MUX41 U11183 ( .I0(n22952), .I1(n22953), .I2(n22954), .I3(n22955), .S0(
        n26227), .S1(n26345), .ZN(n22951) );
  MUX41 U11184 ( .I0(ram[6939]), .I1(ram[6931]), .I2(ram[6923]), .I3(
        ram[6915]), .S0(n27158), .S1(n26683), .ZN(n22955) );
  MUX41 U11185 ( .I0(ram[6971]), .I1(ram[6963]), .I2(ram[6955]), .I3(
        ram[6947]), .S0(n27158), .S1(n26683), .ZN(n22953) );
  MUX41 U11186 ( .I0(ram[7035]), .I1(ram[7027]), .I2(ram[7019]), .I3(
        ram[7011]), .S0(n27158), .S1(n26683), .ZN(n22952) );
  MUX41 U11187 ( .I0(n22887), .I1(n22888), .I2(n22889), .I3(n22890), .S0(
        n26227), .S1(n26345), .ZN(n22886) );
  MUX41 U11188 ( .I0(ram[5435]), .I1(ram[5427]), .I2(ram[5419]), .I3(
        ram[5411]), .S0(n27155), .S1(n26680), .ZN(n22888) );
  MUX41 U11189 ( .I0(ram[5403]), .I1(ram[5395]), .I2(ram[5387]), .I3(
        ram[5379]), .S0(n27155), .S1(n26680), .ZN(n22890) );
  MUX41 U11190 ( .I0(ram[5499]), .I1(ram[5491]), .I2(ram[5483]), .I3(
        ram[5475]), .S0(n27155), .S1(n26680), .ZN(n22887) );
  MUX41 U11191 ( .I0(n22907), .I1(n22908), .I2(n22909), .I3(n22910), .S0(
        n26227), .S1(n26345), .ZN(n22906) );
  MUX41 U11192 ( .I0(ram[5947]), .I1(ram[5939]), .I2(ram[5931]), .I3(
        ram[5923]), .S0(n27156), .S1(n26681), .ZN(n22908) );
  MUX41 U11193 ( .I0(ram[5915]), .I1(ram[5907]), .I2(ram[5899]), .I3(
        ram[5891]), .S0(n27156), .S1(n26681), .ZN(n22910) );
  MUX41 U11194 ( .I0(ram[6011]), .I1(ram[6003]), .I2(ram[5995]), .I3(
        ram[5987]), .S0(n27156), .S1(n26681), .ZN(n22907) );
  MUX41 U11195 ( .I0(n22847), .I1(n22848), .I2(n22849), .I3(n22850), .S0(
        n26226), .S1(n26344), .ZN(n22846) );
  MUX41 U11196 ( .I0(ram[4411]), .I1(ram[4403]), .I2(ram[4395]), .I3(
        ram[4387]), .S0(n27152), .S1(n26677), .ZN(n22848) );
  MUX41 U11197 ( .I0(ram[4379]), .I1(ram[4371]), .I2(ram[4363]), .I3(
        ram[4355]), .S0(n27152), .S1(n26677), .ZN(n22850) );
  MUX41 U11198 ( .I0(ram[4475]), .I1(ram[4467]), .I2(ram[4459]), .I3(
        ram[4451]), .S0(n27152), .S1(n26677), .ZN(n22847) );
  MUX41 U11199 ( .I0(n22867), .I1(n22868), .I2(n22869), .I3(n22870), .S0(
        n26226), .S1(n26344), .ZN(n22866) );
  MUX41 U11200 ( .I0(ram[4891]), .I1(ram[4883]), .I2(ram[4875]), .I3(
        ram[4867]), .S0(n27153), .S1(n26678), .ZN(n22870) );
  MUX41 U11201 ( .I0(ram[4923]), .I1(ram[4915]), .I2(ram[4907]), .I3(
        ram[4899]), .S0(n27153), .S1(n26678), .ZN(n22868) );
  MUX41 U11202 ( .I0(ram[4987]), .I1(ram[4979]), .I2(ram[4971]), .I3(
        ram[4963]), .S0(n27154), .S1(n26679), .ZN(n22867) );
  MUX41 U11203 ( .I0(n23143), .I1(n23144), .I2(n23145), .I3(n23146), .S0(
        n26230), .S1(n26348), .ZN(n23142) );
  MUX41 U11204 ( .I0(ram[11579]), .I1(ram[11571]), .I2(ram[11563]), .I3(
        ram[11555]), .S0(n27169), .S1(n26694), .ZN(n23144) );
  MUX41 U11205 ( .I0(ram[11547]), .I1(ram[11539]), .I2(ram[11531]), .I3(
        ram[11523]), .S0(n27169), .S1(n26694), .ZN(n23146) );
  MUX41 U11206 ( .I0(ram[11643]), .I1(ram[11635]), .I2(ram[11627]), .I3(
        ram[11619]), .S0(n27170), .S1(n26695), .ZN(n23143) );
  MUX41 U11207 ( .I0(n23163), .I1(n23164), .I2(n23165), .I3(n23166), .S0(
        n26231), .S1(n26349), .ZN(n23162) );
  MUX41 U11208 ( .I0(ram[12091]), .I1(ram[12083]), .I2(ram[12075]), .I3(
        ram[12067]), .S0(n27171), .S1(n26696), .ZN(n23164) );
  MUX41 U11209 ( .I0(ram[12059]), .I1(ram[12051]), .I2(ram[12043]), .I3(
        ram[12035]), .S0(n27171), .S1(n26696), .ZN(n23166) );
  MUX41 U11210 ( .I0(ram[12155]), .I1(ram[12147]), .I2(ram[12139]), .I3(
        ram[12131]), .S0(n27171), .S1(n26696), .ZN(n23163) );
  MUX41 U11211 ( .I0(n23103), .I1(n23104), .I2(n23105), .I3(n23106), .S0(
        n26230), .S1(n26348), .ZN(n23102) );
  MUX41 U11212 ( .I0(ram[10555]), .I1(ram[10547]), .I2(ram[10539]), .I3(
        ram[10531]), .S0(n27167), .S1(n26692), .ZN(n23104) );
  MUX41 U11213 ( .I0(ram[10523]), .I1(ram[10515]), .I2(ram[10507]), .I3(
        ram[10499]), .S0(n27167), .S1(n26692), .ZN(n23106) );
  MUX41 U11214 ( .I0(ram[10619]), .I1(ram[10611]), .I2(ram[10603]), .I3(
        ram[10595]), .S0(n27167), .S1(n26692), .ZN(n23103) );
  MUX41 U11215 ( .I0(n23123), .I1(n23124), .I2(n23125), .I3(n23126), .S0(
        n26230), .S1(n26348), .ZN(n23122) );
  MUX41 U11216 ( .I0(ram[11035]), .I1(ram[11027]), .I2(ram[11019]), .I3(
        ram[11011]), .S0(n27168), .S1(n26693), .ZN(n23126) );
  MUX41 U11217 ( .I0(ram[11067]), .I1(ram[11059]), .I2(ram[11051]), .I3(
        ram[11043]), .S0(n27168), .S1(n26693), .ZN(n23124) );
  MUX41 U11218 ( .I0(ram[11131]), .I1(ram[11123]), .I2(ram[11115]), .I3(
        ram[11107]), .S0(n27168), .S1(n26693), .ZN(n23123) );
  MUX41 U11219 ( .I0(n23058), .I1(n23059), .I2(n23060), .I3(n23061), .S0(
        n26229), .S1(n26347), .ZN(n23057) );
  MUX41 U11220 ( .I0(ram[9531]), .I1(ram[9523]), .I2(ram[9515]), .I3(
        ram[9507]), .S0(n27164), .S1(n26689), .ZN(n23059) );
  MUX41 U11221 ( .I0(ram[9499]), .I1(ram[9491]), .I2(ram[9483]), .I3(
        ram[9475]), .S0(n27164), .S1(n26689), .ZN(n23061) );
  MUX41 U11222 ( .I0(ram[9595]), .I1(ram[9587]), .I2(ram[9579]), .I3(
        ram[9571]), .S0(n27165), .S1(n26690), .ZN(n23058) );
  MUX41 U11223 ( .I0(n23078), .I1(n23079), .I2(n23080), .I3(n23081), .S0(
        n26229), .S1(n26347), .ZN(n23077) );
  MUX41 U11224 ( .I0(ram[10043]), .I1(ram[10035]), .I2(ram[10027]), .I3(
        ram[10019]), .S0(n27166), .S1(n26691), .ZN(n23079) );
  MUX41 U11225 ( .I0(ram[10011]), .I1(ram[10003]), .I2(ram[9995]), .I3(
        ram[9987]), .S0(n27166), .S1(n26691), .ZN(n23081) );
  MUX41 U11226 ( .I0(ram[10107]), .I1(ram[10099]), .I2(ram[10091]), .I3(
        ram[10083]), .S0(n27166), .S1(n26691), .ZN(n23078) );
  MUX41 U11227 ( .I0(n23018), .I1(n23019), .I2(n23020), .I3(n23021), .S0(
        n26228), .S1(n26346), .ZN(n23017) );
  MUX41 U11228 ( .I0(ram[8507]), .I1(ram[8499]), .I2(ram[8491]), .I3(
        ram[8483]), .S0(n27162), .S1(n26687), .ZN(n23019) );
  MUX41 U11229 ( .I0(ram[8475]), .I1(ram[8467]), .I2(ram[8459]), .I3(
        ram[8451]), .S0(n27162), .S1(n26687), .ZN(n23021) );
  MUX41 U11230 ( .I0(ram[8571]), .I1(ram[8563]), .I2(ram[8555]), .I3(
        ram[8547]), .S0(n27162), .S1(n26687), .ZN(n23018) );
  MUX41 U11231 ( .I0(n23038), .I1(n23039), .I2(n23040), .I3(n23041), .S0(
        n26229), .S1(n26347), .ZN(n23037) );
  MUX41 U11232 ( .I0(ram[8987]), .I1(ram[8979]), .I2(ram[8971]), .I3(
        ram[8963]), .S0(n27163), .S1(n26688), .ZN(n23041) );
  MUX41 U11233 ( .I0(ram[9019]), .I1(ram[9011]), .I2(ram[9003]), .I3(
        ram[8995]), .S0(n27163), .S1(n26688), .ZN(n23039) );
  MUX41 U11234 ( .I0(ram[9083]), .I1(ram[9075]), .I2(ram[9067]), .I3(
        ram[9059]), .S0(n27163), .S1(n26688), .ZN(n23038) );
  MUX41 U11235 ( .I0(n23998), .I1(n23999), .I2(n24000), .I3(n24001), .S0(
        n26243), .S1(n26361), .ZN(n23997) );
  MUX41 U11236 ( .I0(ram[15644]), .I1(ram[15636]), .I2(ram[15628]), .I3(
        ram[15620]), .S0(n27219), .S1(n26744), .ZN(n24001) );
  MUX41 U11237 ( .I0(ram[15676]), .I1(ram[15668]), .I2(ram[15660]), .I3(
        ram[15652]), .S0(n27219), .S1(n26744), .ZN(n23999) );
  MUX41 U11238 ( .I0(ram[15740]), .I1(ram[15732]), .I2(ram[15724]), .I3(
        ram[15716]), .S0(n27219), .S1(n26744), .ZN(n23998) );
  MUX41 U11239 ( .I0(n24018), .I1(n24019), .I2(n24020), .I3(n24021), .S0(
        n26243), .S1(n26361), .ZN(n24017) );
  MUX41 U11240 ( .I0(ram[16156]), .I1(ram[16148]), .I2(ram[16140]), .I3(
        ram[16132]), .S0(n27220), .S1(n26745), .ZN(n24021) );
  MUX41 U11241 ( .I0(ram[16188]), .I1(ram[16180]), .I2(ram[16172]), .I3(
        ram[16164]), .S0(n27220), .S1(n26745), .ZN(n24019) );
  MUX41 U11242 ( .I0(ram[16252]), .I1(ram[16244]), .I2(ram[16236]), .I3(
        ram[16228]), .S0(n27220), .S1(n26745), .ZN(n24018) );
  MUX41 U11243 ( .I0(n23978), .I1(n23979), .I2(n23980), .I3(n23981), .S0(
        n26242), .S1(n26360), .ZN(n23977) );
  MUX41 U11244 ( .I0(ram[15132]), .I1(ram[15124]), .I2(ram[15116]), .I3(
        ram[15108]), .S0(n27217), .S1(n26742), .ZN(n23981) );
  MUX41 U11245 ( .I0(ram[15164]), .I1(ram[15156]), .I2(ram[15148]), .I3(
        ram[15140]), .S0(n27217), .S1(n26742), .ZN(n23979) );
  MUX41 U11246 ( .I0(ram[15228]), .I1(ram[15220]), .I2(ram[15212]), .I3(
        ram[15204]), .S0(n27218), .S1(n26743), .ZN(n23978) );
  MUX41 U11247 ( .I0(n23958), .I1(n23959), .I2(n23960), .I3(n23961), .S0(
        n26242), .S1(n26360), .ZN(n23957) );
  MUX41 U11248 ( .I0(ram[14620]), .I1(ram[14612]), .I2(ram[14604]), .I3(
        ram[14596]), .S0(n27216), .S1(n26741), .ZN(n23961) );
  MUX41 U11249 ( .I0(ram[14652]), .I1(ram[14644]), .I2(ram[14636]), .I3(
        ram[14628]), .S0(n27216), .S1(n26741), .ZN(n23959) );
  MUX41 U11250 ( .I0(ram[14716]), .I1(ram[14708]), .I2(ram[14700]), .I3(
        ram[14692]), .S0(n27216), .S1(n26741), .ZN(n23958) );
  MUX41 U11251 ( .I0(n23913), .I1(n23914), .I2(n23915), .I3(n23916), .S0(
        n26241), .S1(n26359), .ZN(n23912) );
  MUX41 U11252 ( .I0(ram[13596]), .I1(ram[13588]), .I2(ram[13580]), .I3(
        ram[13572]), .S0(n27214), .S1(n26739), .ZN(n23916) );
  MUX41 U11253 ( .I0(ram[13628]), .I1(ram[13620]), .I2(ram[13612]), .I3(
        ram[13604]), .S0(n27214), .S1(n26739), .ZN(n23914) );
  MUX41 U11254 ( .I0(ram[13692]), .I1(ram[13684]), .I2(ram[13676]), .I3(
        ram[13668]), .S0(n27214), .S1(n26739), .ZN(n23913) );
  MUX41 U11255 ( .I0(n23933), .I1(n23934), .I2(n23935), .I3(n23936), .S0(
        n26242), .S1(n26360), .ZN(n23932) );
  MUX41 U11256 ( .I0(ram[14108]), .I1(ram[14100]), .I2(ram[14092]), .I3(
        ram[14084]), .S0(n27215), .S1(n26740), .ZN(n23936) );
  MUX41 U11257 ( .I0(ram[14140]), .I1(ram[14132]), .I2(ram[14124]), .I3(
        ram[14116]), .S0(n27215), .S1(n26740), .ZN(n23934) );
  MUX41 U11258 ( .I0(ram[14204]), .I1(ram[14196]), .I2(ram[14188]), .I3(
        ram[14180]), .S0(n27215), .S1(n26740), .ZN(n23933) );
  MUX41 U11259 ( .I0(n23893), .I1(n23894), .I2(n23895), .I3(n23896), .S0(
        n26241), .S1(n26359), .ZN(n23892) );
  MUX41 U11260 ( .I0(ram[13084]), .I1(ram[13076]), .I2(ram[13068]), .I3(
        ram[13060]), .S0(n27212), .S1(n26737), .ZN(n23896) );
  MUX41 U11261 ( .I0(ram[13116]), .I1(ram[13108]), .I2(ram[13100]), .I3(
        ram[13092]), .S0(n27212), .S1(n26737), .ZN(n23894) );
  MUX41 U11262 ( .I0(ram[13180]), .I1(ram[13172]), .I2(ram[13164]), .I3(
        ram[13156]), .S0(n27213), .S1(n26738), .ZN(n23893) );
  MUX41 U11263 ( .I0(n23873), .I1(n23874), .I2(n23875), .I3(n23876), .S0(
        n26241), .S1(n26359), .ZN(n23872) );
  MUX41 U11264 ( .I0(ram[12572]), .I1(ram[12564]), .I2(ram[12556]), .I3(
        ram[12548]), .S0(n27211), .S1(n26736), .ZN(n23876) );
  MUX41 U11265 ( .I0(ram[12604]), .I1(ram[12596]), .I2(ram[12588]), .I3(
        ram[12580]), .S0(n27211), .S1(n26736), .ZN(n23874) );
  MUX41 U11266 ( .I0(ram[12668]), .I1(ram[12660]), .I2(ram[12652]), .I3(
        ram[12644]), .S0(n27211), .S1(n26736), .ZN(n23873) );
  MUX41 U11267 ( .I0(n23656), .I1(n23657), .I2(n23658), .I3(n23659), .S0(
        n26238), .S1(n26356), .ZN(n23655) );
  MUX41 U11268 ( .I0(ram[7484]), .I1(ram[7476]), .I2(ram[7468]), .I3(
        ram[7460]), .S0(n27199), .S1(n26724), .ZN(n23657) );
  MUX41 U11269 ( .I0(ram[7452]), .I1(ram[7444]), .I2(ram[7436]), .I3(
        ram[7428]), .S0(n27199), .S1(n26724), .ZN(n23659) );
  MUX41 U11270 ( .I0(ram[7548]), .I1(ram[7540]), .I2(ram[7532]), .I3(
        ram[7524]), .S0(n27199), .S1(n26724), .ZN(n23656) );
  MUX41 U11271 ( .I0(n23676), .I1(n23677), .I2(n23678), .I3(n23679), .S0(
        n26238), .S1(n26356), .ZN(n23675) );
  MUX41 U11272 ( .I0(ram[7964]), .I1(ram[7956]), .I2(ram[7948]), .I3(
        ram[7940]), .S0(n27200), .S1(n26725), .ZN(n23679) );
  MUX41 U11273 ( .I0(ram[7996]), .I1(ram[7988]), .I2(ram[7980]), .I3(
        ram[7972]), .S0(n27200), .S1(n26725), .ZN(n23677) );
  MUX41 U11274 ( .I0(ram[8060]), .I1(ram[8052]), .I2(ram[8044]), .I3(
        ram[8036]), .S0(n27200), .S1(n26725), .ZN(n23676) );
  MUX41 U11275 ( .I0(n23616), .I1(n23617), .I2(n23618), .I3(n23619), .S0(
        n26237), .S1(n26355), .ZN(n23615) );
  MUX41 U11276 ( .I0(ram[6428]), .I1(ram[6420]), .I2(ram[6412]), .I3(
        ram[6404]), .S0(n27196), .S1(n26721), .ZN(n23619) );
  MUX41 U11277 ( .I0(ram[6460]), .I1(ram[6452]), .I2(ram[6444]), .I3(
        ram[6436]), .S0(n27196), .S1(n26721), .ZN(n23617) );
  MUX41 U11278 ( .I0(ram[6524]), .I1(ram[6516]), .I2(ram[6508]), .I3(
        ram[6500]), .S0(n27197), .S1(n26722), .ZN(n23616) );
  MUX41 U11279 ( .I0(n23636), .I1(n23637), .I2(n23638), .I3(n23639), .S0(
        n26237), .S1(n26355), .ZN(n23635) );
  MUX41 U11280 ( .I0(ram[6940]), .I1(ram[6932]), .I2(ram[6924]), .I3(
        ram[6916]), .S0(n27198), .S1(n26723), .ZN(n23639) );
  MUX41 U11281 ( .I0(ram[6972]), .I1(ram[6964]), .I2(ram[6956]), .I3(
        ram[6948]), .S0(n27198), .S1(n26723), .ZN(n23637) );
  MUX41 U11282 ( .I0(ram[7036]), .I1(ram[7028]), .I2(ram[7020]), .I3(
        ram[7012]), .S0(n27198), .S1(n26723), .ZN(n23636) );
  MUX41 U11283 ( .I0(n23571), .I1(n23572), .I2(n23573), .I3(n23574), .S0(
        n26236), .S1(n26354), .ZN(n23570) );
  MUX41 U11284 ( .I0(ram[5436]), .I1(ram[5428]), .I2(ram[5420]), .I3(
        ram[5412]), .S0(n27194), .S1(n26719), .ZN(n23572) );
  MUX41 U11285 ( .I0(ram[5404]), .I1(ram[5396]), .I2(ram[5388]), .I3(
        ram[5380]), .S0(n27194), .S1(n26719), .ZN(n23574) );
  MUX41 U11286 ( .I0(ram[5500]), .I1(ram[5492]), .I2(ram[5484]), .I3(
        ram[5476]), .S0(n27194), .S1(n26719), .ZN(n23571) );
  MUX41 U11287 ( .I0(n23591), .I1(n23592), .I2(n23593), .I3(n23594), .S0(
        n26237), .S1(n26355), .ZN(n23590) );
  MUX41 U11288 ( .I0(ram[5948]), .I1(ram[5940]), .I2(ram[5932]), .I3(
        ram[5924]), .S0(n27195), .S1(n26720), .ZN(n23592) );
  MUX41 U11289 ( .I0(ram[5916]), .I1(ram[5908]), .I2(ram[5900]), .I3(
        ram[5892]), .S0(n27195), .S1(n26720), .ZN(n23594) );
  MUX41 U11290 ( .I0(ram[6012]), .I1(ram[6004]), .I2(ram[5996]), .I3(
        ram[5988]), .S0(n27195), .S1(n26720), .ZN(n23591) );
  MUX41 U11291 ( .I0(n23531), .I1(n23532), .I2(n23533), .I3(n23534), .S0(
        n26236), .S1(n26354), .ZN(n23530) );
  MUX41 U11292 ( .I0(ram[4412]), .I1(ram[4404]), .I2(ram[4396]), .I3(
        ram[4388]), .S0(n27192), .S1(n26717), .ZN(n23532) );
  MUX41 U11293 ( .I0(ram[4380]), .I1(ram[4372]), .I2(ram[4364]), .I3(
        ram[4356]), .S0(n27191), .S1(n26716), .ZN(n23534) );
  MUX41 U11294 ( .I0(ram[4476]), .I1(ram[4468]), .I2(ram[4460]), .I3(
        ram[4452]), .S0(n27192), .S1(n26717), .ZN(n23531) );
  MUX41 U11295 ( .I0(n23551), .I1(n23552), .I2(n23553), .I3(n23554), .S0(
        n26236), .S1(n26354), .ZN(n23550) );
  MUX41 U11296 ( .I0(ram[4892]), .I1(ram[4884]), .I2(ram[4876]), .I3(
        ram[4868]), .S0(n27193), .S1(n26718), .ZN(n23554) );
  MUX41 U11297 ( .I0(ram[4924]), .I1(ram[4916]), .I2(ram[4908]), .I3(
        ram[4900]), .S0(n27193), .S1(n26718), .ZN(n23552) );
  MUX41 U11298 ( .I0(ram[4988]), .I1(ram[4980]), .I2(ram[4972]), .I3(
        ram[4964]), .S0(n27193), .S1(n26718), .ZN(n23551) );
  MUX41 U11299 ( .I0(n23827), .I1(n23828), .I2(n23829), .I3(n23830), .S0(
        n26240), .S1(n26358), .ZN(n23826) );
  MUX41 U11300 ( .I0(ram[11580]), .I1(ram[11572]), .I2(ram[11564]), .I3(
        ram[11556]), .S0(n27209), .S1(n26734), .ZN(n23828) );
  MUX41 U11301 ( .I0(ram[11548]), .I1(ram[11540]), .I2(ram[11532]), .I3(
        ram[11524]), .S0(n27209), .S1(n26734), .ZN(n23830) );
  MUX41 U11302 ( .I0(ram[11644]), .I1(ram[11636]), .I2(ram[11628]), .I3(
        ram[11620]), .S0(n27209), .S1(n26734), .ZN(n23827) );
  MUX41 U11303 ( .I0(n23847), .I1(n23848), .I2(n23849), .I3(n23850), .S0(
        n26240), .S1(n26358), .ZN(n23846) );
  MUX41 U11304 ( .I0(ram[12092]), .I1(ram[12084]), .I2(ram[12076]), .I3(
        ram[12068]), .S0(n27210), .S1(n26735), .ZN(n23848) );
  MUX41 U11305 ( .I0(ram[12060]), .I1(ram[12052]), .I2(ram[12044]), .I3(
        ram[12036]), .S0(n27210), .S1(n26735), .ZN(n23850) );
  MUX41 U11306 ( .I0(ram[12156]), .I1(ram[12148]), .I2(ram[12140]), .I3(
        ram[12132]), .S0(n27210), .S1(n26735), .ZN(n23847) );
  MUX41 U11307 ( .I0(n23787), .I1(n23788), .I2(n23789), .I3(n23790), .S0(
        n26239), .S1(n26357), .ZN(n23786) );
  MUX41 U11308 ( .I0(ram[10556]), .I1(ram[10548]), .I2(ram[10540]), .I3(
        ram[10532]), .S0(n27206), .S1(n26731), .ZN(n23788) );
  MUX41 U11309 ( .I0(ram[10524]), .I1(ram[10516]), .I2(ram[10508]), .I3(
        ram[10500]), .S0(n27206), .S1(n26731), .ZN(n23790) );
  MUX41 U11310 ( .I0(ram[10620]), .I1(ram[10612]), .I2(ram[10604]), .I3(
        ram[10596]), .S0(n27206), .S1(n26731), .ZN(n23787) );
  MUX41 U11311 ( .I0(n23807), .I1(n23808), .I2(n23809), .I3(n23810), .S0(
        n26240), .S1(n26358), .ZN(n23806) );
  MUX41 U11312 ( .I0(ram[11036]), .I1(ram[11028]), .I2(ram[11020]), .I3(
        ram[11012]), .S0(n27207), .S1(n26732), .ZN(n23810) );
  MUX41 U11313 ( .I0(ram[11068]), .I1(ram[11060]), .I2(ram[11052]), .I3(
        ram[11044]), .S0(n27208), .S1(n26733), .ZN(n23808) );
  MUX41 U11314 ( .I0(ram[11132]), .I1(ram[11124]), .I2(ram[11116]), .I3(
        ram[11108]), .S0(n27208), .S1(n26733), .ZN(n23807) );
  MUX41 U11315 ( .I0(n23742), .I1(n23743), .I2(n23744), .I3(n23745), .S0(
        n26239), .S1(n26357), .ZN(n23741) );
  MUX41 U11316 ( .I0(ram[9532]), .I1(ram[9524]), .I2(ram[9516]), .I3(
        ram[9508]), .S0(n27204), .S1(n26729), .ZN(n23743) );
  MUX41 U11317 ( .I0(ram[9500]), .I1(ram[9492]), .I2(ram[9484]), .I3(
        ram[9476]), .S0(n27204), .S1(n26729), .ZN(n23745) );
  MUX41 U11318 ( .I0(ram[9596]), .I1(ram[9588]), .I2(ram[9580]), .I3(
        ram[9572]), .S0(n27204), .S1(n26729), .ZN(n23742) );
  MUX41 U11319 ( .I0(n23762), .I1(n23763), .I2(n23764), .I3(n23765), .S0(
        n26239), .S1(n26357), .ZN(n23761) );
  MUX41 U11320 ( .I0(ram[10044]), .I1(ram[10036]), .I2(ram[10028]), .I3(
        ram[10020]), .S0(n27205), .S1(n26730), .ZN(n23763) );
  MUX41 U11321 ( .I0(ram[10012]), .I1(ram[10004]), .I2(ram[9996]), .I3(
        ram[9988]), .S0(n27205), .S1(n26730), .ZN(n23765) );
  MUX41 U11322 ( .I0(ram[10108]), .I1(ram[10100]), .I2(ram[10092]), .I3(
        ram[10084]), .S0(n27205), .S1(n26730), .ZN(n23762) );
  MUX41 U11323 ( .I0(n23702), .I1(n23703), .I2(n23704), .I3(n23705), .S0(
        n26238), .S1(n26356), .ZN(n23701) );
  MUX41 U11324 ( .I0(ram[8508]), .I1(ram[8500]), .I2(ram[8492]), .I3(
        ram[8484]), .S0(n27201), .S1(n26726), .ZN(n23703) );
  MUX41 U11325 ( .I0(ram[8476]), .I1(ram[8468]), .I2(ram[8460]), .I3(
        ram[8452]), .S0(n27201), .S1(n26726), .ZN(n23705) );
  MUX41 U11326 ( .I0(ram[8572]), .I1(ram[8564]), .I2(ram[8556]), .I3(
        ram[8548]), .S0(n27202), .S1(n26727), .ZN(n23702) );
  MUX41 U11327 ( .I0(n23722), .I1(n23723), .I2(n23724), .I3(n23725), .S0(
        n26239), .S1(n26357), .ZN(n23721) );
  MUX41 U11328 ( .I0(ram[8988]), .I1(ram[8980]), .I2(ram[8972]), .I3(
        ram[8964]), .S0(n27203), .S1(n26728), .ZN(n23725) );
  MUX41 U11329 ( .I0(ram[9020]), .I1(ram[9012]), .I2(ram[9004]), .I3(
        ram[8996]), .S0(n27203), .S1(n26728), .ZN(n23723) );
  MUX41 U11330 ( .I0(ram[9084]), .I1(ram[9076]), .I2(ram[9068]), .I3(
        ram[9060]), .S0(n27203), .S1(n26728), .ZN(n23722) );
  MUX41 U11331 ( .I0(n24682), .I1(n24683), .I2(n24684), .I3(n24685), .S0(
        n26252), .S1(n26370), .ZN(n24681) );
  MUX41 U11332 ( .I0(ram[15645]), .I1(ram[15637]), .I2(ram[15629]), .I3(
        ram[15621]), .S0(n27258), .S1(n26783), .ZN(n24685) );
  MUX41 U11333 ( .I0(ram[15677]), .I1(ram[15669]), .I2(ram[15661]), .I3(
        ram[15653]), .S0(n27258), .S1(n26783), .ZN(n24683) );
  MUX41 U11334 ( .I0(ram[15741]), .I1(ram[15733]), .I2(ram[15725]), .I3(
        ram[15717]), .S0(n27258), .S1(n26783), .ZN(n24682) );
  MUX41 U11335 ( .I0(n24702), .I1(n24703), .I2(n24704), .I3(n24705), .S0(
        n26253), .S1(n26371), .ZN(n24701) );
  MUX41 U11336 ( .I0(ram[16157]), .I1(ram[16149]), .I2(ram[16141]), .I3(
        ram[16133]), .S0(n27259), .S1(n26784), .ZN(n24705) );
  MUX41 U11337 ( .I0(ram[16189]), .I1(ram[16181]), .I2(ram[16173]), .I3(
        ram[16165]), .S0(n27259), .S1(n26784), .ZN(n24703) );
  MUX41 U11338 ( .I0(ram[16253]), .I1(ram[16245]), .I2(ram[16237]), .I3(
        ram[16229]), .S0(n27259), .S1(n26784), .ZN(n24702) );
  MUX41 U11339 ( .I0(n24662), .I1(n24663), .I2(n24664), .I3(n24665), .S0(
        n26252), .S1(n26370), .ZN(n24661) );
  MUX41 U11340 ( .I0(ram[15133]), .I1(ram[15125]), .I2(ram[15117]), .I3(
        ram[15109]), .S0(n27257), .S1(n26782), .ZN(n24665) );
  MUX41 U11341 ( .I0(ram[15165]), .I1(ram[15157]), .I2(ram[15149]), .I3(
        ram[15141]), .S0(n27257), .S1(n26782), .ZN(n24663) );
  MUX41 U11342 ( .I0(ram[15229]), .I1(ram[15221]), .I2(ram[15213]), .I3(
        ram[15205]), .S0(n27257), .S1(n26782), .ZN(n24662) );
  MUX41 U11343 ( .I0(n24642), .I1(n24643), .I2(n24644), .I3(n24645), .S0(
        n26252), .S1(n26370), .ZN(n24641) );
  MUX41 U11344 ( .I0(ram[14621]), .I1(ram[14613]), .I2(ram[14605]), .I3(
        ram[14597]), .S0(n27255), .S1(n26780), .ZN(n24645) );
  MUX41 U11345 ( .I0(ram[14653]), .I1(ram[14645]), .I2(ram[14637]), .I3(
        ram[14629]), .S0(n27256), .S1(n26781), .ZN(n24643) );
  MUX41 U11346 ( .I0(ram[14717]), .I1(ram[14709]), .I2(ram[14701]), .I3(
        ram[14693]), .S0(n27256), .S1(n26781), .ZN(n24642) );
  MUX41 U11347 ( .I0(n24597), .I1(n24598), .I2(n24599), .I3(n24600), .S0(
        n26251), .S1(n26369), .ZN(n24596) );
  MUX41 U11348 ( .I0(ram[13597]), .I1(ram[13589]), .I2(ram[13581]), .I3(
        ram[13573]), .S0(n27253), .S1(n26778), .ZN(n24600) );
  MUX41 U11349 ( .I0(ram[13629]), .I1(ram[13621]), .I2(ram[13613]), .I3(
        ram[13605]), .S0(n27253), .S1(n26778), .ZN(n24598) );
  MUX41 U11350 ( .I0(ram[13693]), .I1(ram[13685]), .I2(ram[13677]), .I3(
        ram[13669]), .S0(n27253), .S1(n26778), .ZN(n24597) );
  MUX41 U11351 ( .I0(n24617), .I1(n24618), .I2(n24619), .I3(n24620), .S0(
        n26251), .S1(n26369), .ZN(n24616) );
  MUX41 U11352 ( .I0(ram[14109]), .I1(ram[14101]), .I2(ram[14093]), .I3(
        ram[14085]), .S0(n27254), .S1(n26779), .ZN(n24620) );
  MUX41 U11353 ( .I0(ram[14141]), .I1(ram[14133]), .I2(ram[14125]), .I3(
        ram[14117]), .S0(n27254), .S1(n26779), .ZN(n24618) );
  MUX41 U11354 ( .I0(ram[14205]), .I1(ram[14197]), .I2(ram[14189]), .I3(
        ram[14181]), .S0(n27254), .S1(n26779), .ZN(n24617) );
  MUX41 U11355 ( .I0(n24577), .I1(n24578), .I2(n24579), .I3(n24580), .S0(
        n26251), .S1(n26369), .ZN(n24576) );
  MUX41 U11356 ( .I0(ram[13085]), .I1(ram[13077]), .I2(ram[13069]), .I3(
        ram[13061]), .S0(n27252), .S1(n26777), .ZN(n24580) );
  MUX41 U11357 ( .I0(ram[13117]), .I1(ram[13109]), .I2(ram[13101]), .I3(
        ram[13093]), .S0(n27252), .S1(n26777), .ZN(n24578) );
  MUX41 U11358 ( .I0(ram[13181]), .I1(ram[13173]), .I2(ram[13165]), .I3(
        ram[13157]), .S0(n27252), .S1(n26777), .ZN(n24577) );
  MUX41 U11359 ( .I0(n24557), .I1(n24558), .I2(n24559), .I3(n24560), .S0(
        n26251), .S1(n26369), .ZN(n24556) );
  MUX41 U11360 ( .I0(ram[12573]), .I1(ram[12565]), .I2(ram[12557]), .I3(
        ram[12549]), .S0(n27251), .S1(n26776), .ZN(n24560) );
  MUX41 U11361 ( .I0(ram[12605]), .I1(ram[12597]), .I2(ram[12589]), .I3(
        ram[12581]), .S0(n27251), .S1(n26776), .ZN(n24558) );
  MUX41 U11362 ( .I0(ram[12669]), .I1(ram[12661]), .I2(ram[12653]), .I3(
        ram[12645]), .S0(n27251), .S1(n26776), .ZN(n24557) );
  MUX41 U11363 ( .I0(n24340), .I1(n24341), .I2(n24342), .I3(n24343), .S0(
        n26247), .S1(n26365), .ZN(n24339) );
  MUX41 U11364 ( .I0(ram[7485]), .I1(ram[7477]), .I2(ram[7469]), .I3(
        ram[7461]), .S0(n27238), .S1(n26763), .ZN(n24341) );
  MUX41 U11365 ( .I0(ram[7453]), .I1(ram[7445]), .I2(ram[7437]), .I3(
        ram[7429]), .S0(n27238), .S1(n26763), .ZN(n24343) );
  MUX41 U11366 ( .I0(ram[7549]), .I1(ram[7541]), .I2(ram[7533]), .I3(
        ram[7525]), .S0(n27238), .S1(n26763), .ZN(n24340) );
  MUX41 U11367 ( .I0(n24360), .I1(n24361), .I2(n24362), .I3(n24363), .S0(
        n26248), .S1(n26366), .ZN(n24359) );
  MUX41 U11368 ( .I0(ram[7965]), .I1(ram[7957]), .I2(ram[7949]), .I3(
        ram[7941]), .S0(n27239), .S1(n26764), .ZN(n24363) );
  MUX41 U11369 ( .I0(ram[7997]), .I1(ram[7989]), .I2(ram[7981]), .I3(
        ram[7973]), .S0(n27240), .S1(n26765), .ZN(n24361) );
  MUX41 U11370 ( .I0(ram[8061]), .I1(ram[8053]), .I2(ram[8045]), .I3(
        ram[8037]), .S0(n27240), .S1(n26765), .ZN(n24360) );
  MUX41 U11371 ( .I0(n24300), .I1(n24301), .I2(n24302), .I3(n24303), .S0(
        n26247), .S1(n26365), .ZN(n24299) );
  MUX41 U11372 ( .I0(ram[6429]), .I1(ram[6421]), .I2(ram[6413]), .I3(
        ram[6405]), .S0(n27236), .S1(n26761), .ZN(n24303) );
  MUX41 U11373 ( .I0(ram[6461]), .I1(ram[6453]), .I2(ram[6445]), .I3(
        ram[6437]), .S0(n27236), .S1(n26761), .ZN(n24301) );
  MUX41 U11374 ( .I0(ram[6525]), .I1(ram[6517]), .I2(ram[6509]), .I3(
        ram[6501]), .S0(n27236), .S1(n26761), .ZN(n24300) );
  MUX41 U11375 ( .I0(n24320), .I1(n24321), .I2(n24322), .I3(n24323), .S0(
        n26247), .S1(n26365), .ZN(n24319) );
  MUX41 U11376 ( .I0(ram[6941]), .I1(ram[6933]), .I2(ram[6925]), .I3(
        ram[6917]), .S0(n27237), .S1(n26762), .ZN(n24323) );
  MUX41 U11377 ( .I0(ram[6973]), .I1(ram[6965]), .I2(ram[6957]), .I3(
        ram[6949]), .S0(n27237), .S1(n26762), .ZN(n24321) );
  MUX41 U11378 ( .I0(ram[7037]), .I1(ram[7029]), .I2(ram[7021]), .I3(
        ram[7013]), .S0(n27237), .S1(n26762), .ZN(n24320) );
  MUX41 U11379 ( .I0(n24255), .I1(n24256), .I2(n24257), .I3(n24258), .S0(
        n26246), .S1(n26364), .ZN(n24254) );
  MUX41 U11380 ( .I0(ram[5437]), .I1(ram[5429]), .I2(ram[5421]), .I3(
        ram[5413]), .S0(n27233), .S1(n26758), .ZN(n24256) );
  MUX41 U11381 ( .I0(ram[5405]), .I1(ram[5397]), .I2(ram[5389]), .I3(
        ram[5381]), .S0(n27233), .S1(n26758), .ZN(n24258) );
  MUX41 U11382 ( .I0(ram[5501]), .I1(ram[5493]), .I2(ram[5485]), .I3(
        ram[5477]), .S0(n27234), .S1(n26759), .ZN(n24255) );
  MUX41 U11383 ( .I0(n24275), .I1(n24276), .I2(n24277), .I3(n24278), .S0(
        n26247), .S1(n26365), .ZN(n24274) );
  MUX41 U11384 ( .I0(ram[5949]), .I1(ram[5941]), .I2(ram[5933]), .I3(
        ram[5925]), .S0(n27235), .S1(n26760), .ZN(n24276) );
  MUX41 U11385 ( .I0(ram[5917]), .I1(ram[5909]), .I2(ram[5901]), .I3(
        ram[5893]), .S0(n27235), .S1(n26760), .ZN(n24278) );
  MUX41 U11386 ( .I0(ram[6013]), .I1(ram[6005]), .I2(ram[5997]), .I3(
        ram[5989]), .S0(n27235), .S1(n26760), .ZN(n24275) );
  MUX41 U11387 ( .I0(n24215), .I1(n24216), .I2(n24217), .I3(n24218), .S0(
        n26246), .S1(n26364), .ZN(n24214) );
  MUX41 U11388 ( .I0(ram[4413]), .I1(ram[4405]), .I2(ram[4397]), .I3(
        ram[4389]), .S0(n27231), .S1(n26756), .ZN(n24216) );
  MUX41 U11389 ( .I0(ram[4381]), .I1(ram[4373]), .I2(ram[4365]), .I3(
        ram[4357]), .S0(n27231), .S1(n26756), .ZN(n24218) );
  MUX41 U11390 ( .I0(ram[4477]), .I1(ram[4469]), .I2(ram[4461]), .I3(
        ram[4453]), .S0(n27231), .S1(n26756), .ZN(n24215) );
  MUX41 U11391 ( .I0(n24235), .I1(n24236), .I2(n24237), .I3(n24238), .S0(
        n26246), .S1(n26364), .ZN(n24234) );
  MUX41 U11392 ( .I0(ram[4893]), .I1(ram[4885]), .I2(ram[4877]), .I3(
        ram[4869]), .S0(n27232), .S1(n26757), .ZN(n24238) );
  MUX41 U11393 ( .I0(ram[4925]), .I1(ram[4917]), .I2(ram[4909]), .I3(
        ram[4901]), .S0(n27232), .S1(n26757), .ZN(n24236) );
  MUX41 U11394 ( .I0(ram[4989]), .I1(ram[4981]), .I2(ram[4973]), .I3(
        ram[4965]), .S0(n27232), .S1(n26757), .ZN(n24235) );
  MUX41 U11395 ( .I0(n24511), .I1(n24512), .I2(n24513), .I3(n24514), .S0(
        n26250), .S1(n26368), .ZN(n24510) );
  MUX41 U11396 ( .I0(ram[11581]), .I1(ram[11573]), .I2(ram[11565]), .I3(
        ram[11557]), .S0(n27248), .S1(n26773), .ZN(n24512) );
  MUX41 U11397 ( .I0(ram[11549]), .I1(ram[11541]), .I2(ram[11533]), .I3(
        ram[11525]), .S0(n27248), .S1(n26773), .ZN(n24514) );
  MUX41 U11398 ( .I0(ram[11645]), .I1(ram[11637]), .I2(ram[11629]), .I3(
        ram[11621]), .S0(n27248), .S1(n26773), .ZN(n24511) );
  MUX41 U11399 ( .I0(n24531), .I1(n24532), .I2(n24533), .I3(n24534), .S0(
        n26250), .S1(n26368), .ZN(n24530) );
  MUX41 U11400 ( .I0(ram[12093]), .I1(ram[12085]), .I2(ram[12077]), .I3(
        ram[12069]), .S0(n27249), .S1(n26774), .ZN(n24532) );
  MUX41 U11401 ( .I0(ram[12061]), .I1(ram[12053]), .I2(ram[12045]), .I3(
        ram[12037]), .S0(n27249), .S1(n26774), .ZN(n24534) );
  MUX41 U11402 ( .I0(ram[12157]), .I1(ram[12149]), .I2(ram[12141]), .I3(
        ram[12133]), .S0(n27250), .S1(n26775), .ZN(n24531) );
  MUX41 U11403 ( .I0(n24471), .I1(n24472), .I2(n24473), .I3(n24474), .S0(
        n26249), .S1(n26367), .ZN(n24470) );
  MUX41 U11404 ( .I0(ram[10557]), .I1(ram[10549]), .I2(ram[10541]), .I3(
        ram[10533]), .S0(n27246), .S1(n26771), .ZN(n24472) );
  MUX41 U11405 ( .I0(ram[10525]), .I1(ram[10517]), .I2(ram[10509]), .I3(
        ram[10501]), .S0(n27246), .S1(n26771), .ZN(n24474) );
  MUX41 U11406 ( .I0(ram[10621]), .I1(ram[10613]), .I2(ram[10605]), .I3(
        ram[10597]), .S0(n27246), .S1(n26771), .ZN(n24471) );
  MUX41 U11407 ( .I0(n24491), .I1(n24492), .I2(n24493), .I3(n24494), .S0(
        n26250), .S1(n26368), .ZN(n24490) );
  MUX41 U11408 ( .I0(ram[11037]), .I1(ram[11029]), .I2(ram[11021]), .I3(
        ram[11013]), .S0(n27247), .S1(n26772), .ZN(n24494) );
  MUX41 U11409 ( .I0(ram[11069]), .I1(ram[11061]), .I2(ram[11053]), .I3(
        ram[11045]), .S0(n27247), .S1(n26772), .ZN(n24492) );
  MUX41 U11410 ( .I0(ram[11133]), .I1(ram[11125]), .I2(ram[11117]), .I3(
        ram[11109]), .S0(n27247), .S1(n26772), .ZN(n24491) );
  MUX41 U11411 ( .I0(n24426), .I1(n24427), .I2(n24428), .I3(n24429), .S0(
        n26249), .S1(n26367), .ZN(n24425) );
  MUX41 U11412 ( .I0(ram[9533]), .I1(ram[9525]), .I2(ram[9517]), .I3(
        ram[9509]), .S0(n27243), .S1(n26768), .ZN(n24427) );
  MUX41 U11413 ( .I0(ram[9501]), .I1(ram[9493]), .I2(ram[9485]), .I3(
        ram[9477]), .S0(n27243), .S1(n26768), .ZN(n24429) );
  MUX41 U11414 ( .I0(ram[9597]), .I1(ram[9589]), .I2(ram[9581]), .I3(
        ram[9573]), .S0(n27243), .S1(n26768), .ZN(n24426) );
  MUX41 U11415 ( .I0(n24446), .I1(n24447), .I2(n24448), .I3(n24449), .S0(
        n26249), .S1(n26367), .ZN(n24445) );
  MUX41 U11416 ( .I0(ram[10045]), .I1(ram[10037]), .I2(ram[10029]), .I3(
        ram[10021]), .S0(n27244), .S1(n26769), .ZN(n24447) );
  MUX41 U11417 ( .I0(ram[10013]), .I1(ram[10005]), .I2(ram[9997]), .I3(
        ram[9989]), .S0(n27244), .S1(n26769), .ZN(n24449) );
  MUX41 U11418 ( .I0(ram[10109]), .I1(ram[10101]), .I2(ram[10093]), .I3(
        ram[10085]), .S0(n27245), .S1(n26770), .ZN(n24446) );
  MUX41 U11419 ( .I0(n24386), .I1(n24387), .I2(n24388), .I3(n24389), .S0(
        n26248), .S1(n26366), .ZN(n24385) );
  MUX41 U11420 ( .I0(ram[8509]), .I1(ram[8501]), .I2(ram[8493]), .I3(
        ram[8485]), .S0(n27241), .S1(n26766), .ZN(n24387) );
  MUX41 U11421 ( .I0(ram[8477]), .I1(ram[8469]), .I2(ram[8461]), .I3(
        ram[8453]), .S0(n27241), .S1(n26766), .ZN(n24389) );
  MUX41 U11422 ( .I0(ram[8573]), .I1(ram[8565]), .I2(ram[8557]), .I3(
        ram[8549]), .S0(n27241), .S1(n26766), .ZN(n24386) );
  MUX41 U11423 ( .I0(n24406), .I1(n24407), .I2(n24408), .I3(n24409), .S0(
        n26248), .S1(n26366), .ZN(n24405) );
  MUX41 U11424 ( .I0(ram[8989]), .I1(ram[8981]), .I2(ram[8973]), .I3(
        ram[8965]), .S0(n27242), .S1(n26767), .ZN(n24409) );
  MUX41 U11425 ( .I0(ram[9021]), .I1(ram[9013]), .I2(ram[9005]), .I3(
        ram[8997]), .S0(n27242), .S1(n26767), .ZN(n24407) );
  MUX41 U11426 ( .I0(ram[9085]), .I1(ram[9077]), .I2(ram[9069]), .I3(
        ram[9061]), .S0(n27242), .S1(n26767), .ZN(n24406) );
  MUX41 U11427 ( .I0(n25366), .I1(n25367), .I2(n25368), .I3(n25369), .S0(
        n26262), .S1(n26380), .ZN(n25365) );
  MUX41 U11428 ( .I0(ram[15646]), .I1(ram[15638]), .I2(ram[15630]), .I3(
        ram[15622]), .S0(n27297), .S1(n26822), .ZN(n25369) );
  MUX41 U11429 ( .I0(ram[15678]), .I1(ram[15670]), .I2(ram[15662]), .I3(
        ram[15654]), .S0(n27297), .S1(n26822), .ZN(n25367) );
  MUX41 U11430 ( .I0(ram[15742]), .I1(ram[15734]), .I2(ram[15726]), .I3(
        ram[15718]), .S0(n27298), .S1(n26823), .ZN(n25366) );
  MUX41 U11431 ( .I0(n25386), .I1(n25387), .I2(n25388), .I3(n25389), .S0(
        n26263), .S1(n26381), .ZN(n25385) );
  MUX41 U11432 ( .I0(ram[16158]), .I1(ram[16150]), .I2(ram[16142]), .I3(
        ram[16134]), .S0(n27299), .S1(n26824), .ZN(n25389) );
  MUX41 U11433 ( .I0(ram[16190]), .I1(ram[16182]), .I2(ram[16174]), .I3(
        ram[16166]), .S0(n27299), .S1(n26824), .ZN(n25387) );
  MUX41 U11434 ( .I0(ram[16254]), .I1(ram[16246]), .I2(ram[16238]), .I3(
        ram[16230]), .S0(n27299), .S1(n26824), .ZN(n25386) );
  MUX41 U11435 ( .I0(n25346), .I1(n25347), .I2(n25348), .I3(n25349), .S0(
        n26262), .S1(n26380), .ZN(n25345) );
  MUX41 U11436 ( .I0(ram[15134]), .I1(ram[15126]), .I2(ram[15118]), .I3(
        ram[15110]), .S0(n27296), .S1(n26821), .ZN(n25349) );
  MUX41 U11437 ( .I0(ram[15166]), .I1(ram[15158]), .I2(ram[15150]), .I3(
        ram[15142]), .S0(n27296), .S1(n26821), .ZN(n25347) );
  MUX41 U11438 ( .I0(ram[15230]), .I1(ram[15222]), .I2(ram[15214]), .I3(
        ram[15206]), .S0(n27296), .S1(n26821), .ZN(n25346) );
  MUX41 U11439 ( .I0(n25326), .I1(n25327), .I2(n25328), .I3(n25329), .S0(
        n26262), .S1(n26380), .ZN(n25325) );
  MUX41 U11440 ( .I0(ram[14622]), .I1(ram[14614]), .I2(ram[14606]), .I3(
        ram[14598]), .S0(n27295), .S1(n26820), .ZN(n25329) );
  MUX41 U11441 ( .I0(ram[14654]), .I1(ram[14646]), .I2(ram[14638]), .I3(
        ram[14630]), .S0(n27295), .S1(n26820), .ZN(n25327) );
  MUX41 U11442 ( .I0(ram[14718]), .I1(ram[14710]), .I2(ram[14702]), .I3(
        ram[14694]), .S0(n27295), .S1(n26820), .ZN(n25326) );
  MUX41 U11443 ( .I0(n25281), .I1(n25282), .I2(n25283), .I3(n25284), .S0(
        n26261), .S1(n26379), .ZN(n25280) );
  MUX41 U11444 ( .I0(ram[13598]), .I1(ram[13590]), .I2(ram[13582]), .I3(
        ram[13574]), .S0(n27292), .S1(n26817), .ZN(n25284) );
  MUX41 U11445 ( .I0(ram[13630]), .I1(ram[13622]), .I2(ram[13614]), .I3(
        ram[13606]), .S0(n27292), .S1(n26817), .ZN(n25282) );
  MUX41 U11446 ( .I0(ram[13694]), .I1(ram[13686]), .I2(ram[13678]), .I3(
        ram[13670]), .S0(n27293), .S1(n26818), .ZN(n25281) );
  MUX41 U11447 ( .I0(n25301), .I1(n25302), .I2(n25303), .I3(n25304), .S0(
        n26261), .S1(n26379), .ZN(n25300) );
  MUX41 U11448 ( .I0(ram[14110]), .I1(ram[14102]), .I2(ram[14094]), .I3(
        ram[14086]), .S0(n27294), .S1(n26819), .ZN(n25304) );
  MUX41 U11449 ( .I0(ram[14142]), .I1(ram[14134]), .I2(ram[14126]), .I3(
        ram[14118]), .S0(n27294), .S1(n26819), .ZN(n25302) );
  MUX41 U11450 ( .I0(ram[14206]), .I1(ram[14198]), .I2(ram[14190]), .I3(
        ram[14182]), .S0(n27294), .S1(n26819), .ZN(n25301) );
  MUX41 U11451 ( .I0(n25261), .I1(n25262), .I2(n25263), .I3(n25264), .S0(
        n26261), .S1(n26379), .ZN(n25260) );
  MUX41 U11452 ( .I0(ram[13086]), .I1(ram[13078]), .I2(ram[13070]), .I3(
        ram[13062]), .S0(n27291), .S1(n26816), .ZN(n25264) );
  MUX41 U11453 ( .I0(ram[13118]), .I1(ram[13110]), .I2(ram[13102]), .I3(
        ram[13094]), .S0(n27291), .S1(n26816), .ZN(n25262) );
  MUX41 U11454 ( .I0(ram[13182]), .I1(ram[13174]), .I2(ram[13166]), .I3(
        ram[13158]), .S0(n27291), .S1(n26816), .ZN(n25261) );
  MUX41 U11455 ( .I0(n25241), .I1(n25242), .I2(n25243), .I3(n25244), .S0(
        n26260), .S1(n26378), .ZN(n25240) );
  MUX41 U11456 ( .I0(ram[12574]), .I1(ram[12566]), .I2(ram[12558]), .I3(
        ram[12550]), .S0(n27290), .S1(n26815), .ZN(n25244) );
  MUX41 U11457 ( .I0(ram[12606]), .I1(ram[12598]), .I2(ram[12590]), .I3(
        ram[12582]), .S0(n27290), .S1(n26815), .ZN(n25242) );
  MUX41 U11458 ( .I0(ram[12670]), .I1(ram[12662]), .I2(ram[12654]), .I3(
        ram[12646]), .S0(n27290), .S1(n26815), .ZN(n25241) );
  MUX41 U11459 ( .I0(n25024), .I1(n25025), .I2(n25026), .I3(n25027), .S0(
        n26257), .S1(n26375), .ZN(n25023) );
  MUX41 U11460 ( .I0(ram[7486]), .I1(ram[7478]), .I2(ram[7470]), .I3(
        ram[7462]), .S0(n27278), .S1(n26803), .ZN(n25025) );
  MUX41 U11461 ( .I0(ram[7454]), .I1(ram[7446]), .I2(ram[7438]), .I3(
        ram[7430]), .S0(n27278), .S1(n26803), .ZN(n25027) );
  MUX41 U11462 ( .I0(ram[7550]), .I1(ram[7542]), .I2(ram[7534]), .I3(
        ram[7526]), .S0(n27278), .S1(n26803), .ZN(n25024) );
  MUX41 U11463 ( .I0(n25044), .I1(n25045), .I2(n25046), .I3(n25047), .S0(
        n26258), .S1(n26376), .ZN(n25043) );
  MUX41 U11464 ( .I0(ram[7966]), .I1(ram[7958]), .I2(ram[7950]), .I3(
        ram[7942]), .S0(n27279), .S1(n26804), .ZN(n25047) );
  MUX41 U11465 ( .I0(ram[7998]), .I1(ram[7990]), .I2(ram[7982]), .I3(
        ram[7974]), .S0(n27279), .S1(n26804), .ZN(n25045) );
  MUX41 U11466 ( .I0(ram[8062]), .I1(ram[8054]), .I2(ram[8046]), .I3(
        ram[8038]), .S0(n27279), .S1(n26804), .ZN(n25044) );
  MUX41 U11467 ( .I0(n24984), .I1(n24985), .I2(n24986), .I3(n24987), .S0(
        n26257), .S1(n26375), .ZN(n24983) );
  MUX41 U11468 ( .I0(ram[6430]), .I1(ram[6422]), .I2(ram[6414]), .I3(
        ram[6406]), .S0(n27275), .S1(n26800), .ZN(n24987) );
  MUX41 U11469 ( .I0(ram[6462]), .I1(ram[6454]), .I2(ram[6446]), .I3(
        ram[6438]), .S0(n27275), .S1(n26800), .ZN(n24985) );
  MUX41 U11470 ( .I0(ram[6526]), .I1(ram[6518]), .I2(ram[6510]), .I3(
        ram[6502]), .S0(n27275), .S1(n26800), .ZN(n24984) );
  MUX41 U11471 ( .I0(n25004), .I1(n25005), .I2(n25006), .I3(n25007), .S0(
        n26257), .S1(n26375), .ZN(n25003) );
  MUX41 U11472 ( .I0(ram[6942]), .I1(ram[6934]), .I2(ram[6926]), .I3(
        ram[6918]), .S0(n27276), .S1(n26801), .ZN(n25007) );
  MUX41 U11473 ( .I0(ram[6974]), .I1(ram[6966]), .I2(ram[6958]), .I3(
        ram[6950]), .S0(n27276), .S1(n26801), .ZN(n25005) );
  MUX41 U11474 ( .I0(ram[7038]), .I1(ram[7030]), .I2(ram[7022]), .I3(
        ram[7014]), .S0(n27277), .S1(n26802), .ZN(n25004) );
  MUX41 U11475 ( .I0(n24939), .I1(n24940), .I2(n24941), .I3(n24942), .S0(
        n26256), .S1(n26374), .ZN(n24938) );
  MUX41 U11476 ( .I0(ram[5438]), .I1(ram[5430]), .I2(ram[5422]), .I3(
        ram[5414]), .S0(n27273), .S1(n26798), .ZN(n24940) );
  MUX41 U11477 ( .I0(ram[5406]), .I1(ram[5398]), .I2(ram[5390]), .I3(
        ram[5382]), .S0(n27273), .S1(n26798), .ZN(n24942) );
  MUX41 U11478 ( .I0(ram[5502]), .I1(ram[5494]), .I2(ram[5486]), .I3(
        ram[5478]), .S0(n27273), .S1(n26798), .ZN(n24939) );
  MUX41 U11479 ( .I0(n24959), .I1(n24960), .I2(n24961), .I3(n24962), .S0(
        n26256), .S1(n26374), .ZN(n24958) );
  MUX41 U11480 ( .I0(ram[5950]), .I1(ram[5942]), .I2(ram[5934]), .I3(
        ram[5926]), .S0(n27274), .S1(n26799), .ZN(n24960) );
  MUX41 U11481 ( .I0(ram[5918]), .I1(ram[5910]), .I2(ram[5902]), .I3(
        ram[5894]), .S0(n27274), .S1(n26799), .ZN(n24962) );
  MUX41 U11482 ( .I0(ram[6014]), .I1(ram[6006]), .I2(ram[5998]), .I3(
        ram[5990]), .S0(n27274), .S1(n26799), .ZN(n24959) );
  MUX41 U11483 ( .I0(n24899), .I1(n24900), .I2(n24901), .I3(n24902), .S0(
        n26255), .S1(n26373), .ZN(n24898) );
  MUX41 U11484 ( .I0(ram[4414]), .I1(ram[4406]), .I2(ram[4398]), .I3(
        ram[4390]), .S0(n27270), .S1(n26795), .ZN(n24900) );
  MUX41 U11485 ( .I0(ram[4382]), .I1(ram[4374]), .I2(ram[4366]), .I3(
        ram[4358]), .S0(n27270), .S1(n26795), .ZN(n24902) );
  MUX41 U11486 ( .I0(ram[4478]), .I1(ram[4470]), .I2(ram[4462]), .I3(
        ram[4454]), .S0(n27270), .S1(n26795), .ZN(n24899) );
  MUX41 U11487 ( .I0(n24919), .I1(n24920), .I2(n24921), .I3(n24922), .S0(
        n26256), .S1(n26374), .ZN(n24918) );
  MUX41 U11488 ( .I0(ram[4894]), .I1(ram[4886]), .I2(ram[4878]), .I3(
        ram[4870]), .S0(n27271), .S1(n26796), .ZN(n24922) );
  MUX41 U11489 ( .I0(ram[4926]), .I1(ram[4918]), .I2(ram[4910]), .I3(
        ram[4902]), .S0(n27272), .S1(n26797), .ZN(n24920) );
  MUX41 U11490 ( .I0(ram[4990]), .I1(ram[4982]), .I2(ram[4974]), .I3(
        ram[4966]), .S0(n27272), .S1(n26797), .ZN(n24919) );
  MUX41 U11491 ( .I0(n25195), .I1(n25196), .I2(n25197), .I3(n25198), .S0(
        n26260), .S1(n26378), .ZN(n25194) );
  MUX41 U11492 ( .I0(ram[11582]), .I1(ram[11574]), .I2(ram[11566]), .I3(
        ram[11558]), .S0(n27288), .S1(n26813), .ZN(n25196) );
  MUX41 U11493 ( .I0(ram[11550]), .I1(ram[11542]), .I2(ram[11534]), .I3(
        ram[11526]), .S0(n27287), .S1(n26812), .ZN(n25198) );
  MUX41 U11494 ( .I0(ram[11646]), .I1(ram[11638]), .I2(ram[11630]), .I3(
        ram[11622]), .S0(n27288), .S1(n26813), .ZN(n25195) );
  MUX41 U11495 ( .I0(n25215), .I1(n25216), .I2(n25217), .I3(n25218), .S0(
        n26260), .S1(n26378), .ZN(n25214) );
  MUX41 U11496 ( .I0(ram[12094]), .I1(ram[12086]), .I2(ram[12078]), .I3(
        ram[12070]), .S0(n27289), .S1(n26814), .ZN(n25216) );
  MUX41 U11497 ( .I0(ram[12062]), .I1(ram[12054]), .I2(ram[12046]), .I3(
        ram[12038]), .S0(n27289), .S1(n26814), .ZN(n25218) );
  MUX41 U11498 ( .I0(ram[12158]), .I1(ram[12150]), .I2(ram[12142]), .I3(
        ram[12134]), .S0(n27289), .S1(n26814), .ZN(n25215) );
  MUX41 U11499 ( .I0(n25155), .I1(n25156), .I2(n25157), .I3(n25158), .S0(
        n26259), .S1(n26377), .ZN(n25154) );
  MUX41 U11500 ( .I0(ram[10558]), .I1(ram[10550]), .I2(ram[10542]), .I3(
        ram[10534]), .S0(n27285), .S1(n26810), .ZN(n25156) );
  MUX41 U11501 ( .I0(ram[10526]), .I1(ram[10518]), .I2(ram[10510]), .I3(
        ram[10502]), .S0(n27285), .S1(n26810), .ZN(n25158) );
  MUX41 U11502 ( .I0(ram[10622]), .I1(ram[10614]), .I2(ram[10606]), .I3(
        ram[10598]), .S0(n27285), .S1(n26810), .ZN(n25155) );
  MUX41 U11503 ( .I0(n25175), .I1(n25176), .I2(n25177), .I3(n25178), .S0(
        n26259), .S1(n26377), .ZN(n25174) );
  MUX41 U11504 ( .I0(ram[11038]), .I1(ram[11030]), .I2(ram[11022]), .I3(
        ram[11014]), .S0(n27286), .S1(n26811), .ZN(n25178) );
  MUX41 U11505 ( .I0(ram[11070]), .I1(ram[11062]), .I2(ram[11054]), .I3(
        ram[11046]), .S0(n27286), .S1(n26811), .ZN(n25176) );
  MUX41 U11506 ( .I0(ram[11134]), .I1(ram[11126]), .I2(ram[11118]), .I3(
        ram[11110]), .S0(n27286), .S1(n26811), .ZN(n25175) );
  MUX41 U11507 ( .I0(n25110), .I1(n25111), .I2(n25112), .I3(n25113), .S0(
        n26259), .S1(n26377), .ZN(n25109) );
  MUX41 U11508 ( .I0(ram[9534]), .I1(ram[9526]), .I2(ram[9518]), .I3(
        ram[9510]), .S0(n27283), .S1(n26808), .ZN(n25111) );
  MUX41 U11509 ( .I0(ram[9502]), .I1(ram[9494]), .I2(ram[9486]), .I3(
        ram[9478]), .S0(n27283), .S1(n26808), .ZN(n25113) );
  MUX41 U11510 ( .I0(ram[9598]), .I1(ram[9590]), .I2(ram[9582]), .I3(
        ram[9574]), .S0(n27283), .S1(n26808), .ZN(n25110) );
  MUX41 U11511 ( .I0(n25130), .I1(n25131), .I2(n25132), .I3(n25133), .S0(
        n26259), .S1(n26377), .ZN(n25129) );
  MUX41 U11512 ( .I0(ram[10046]), .I1(ram[10038]), .I2(ram[10030]), .I3(
        ram[10022]), .S0(n27284), .S1(n26809), .ZN(n25131) );
  MUX41 U11513 ( .I0(ram[10014]), .I1(ram[10006]), .I2(ram[9998]), .I3(
        ram[9990]), .S0(n27284), .S1(n26809), .ZN(n25133) );
  MUX41 U11514 ( .I0(ram[10110]), .I1(ram[10102]), .I2(ram[10094]), .I3(
        ram[10086]), .S0(n27284), .S1(n26809), .ZN(n25130) );
  MUX41 U11515 ( .I0(n25070), .I1(n25071), .I2(n25072), .I3(n25073), .S0(
        n26258), .S1(n26376), .ZN(n25069) );
  MUX41 U11516 ( .I0(ram[8510]), .I1(ram[8502]), .I2(ram[8494]), .I3(
        ram[8486]), .S0(n27280), .S1(n26805), .ZN(n25071) );
  MUX41 U11517 ( .I0(ram[8478]), .I1(ram[8470]), .I2(ram[8462]), .I3(
        ram[8454]), .S0(n27280), .S1(n26805), .ZN(n25073) );
  MUX41 U11518 ( .I0(ram[8574]), .I1(ram[8566]), .I2(ram[8558]), .I3(
        ram[8550]), .S0(n27280), .S1(n26805), .ZN(n25070) );
  MUX41 U11519 ( .I0(n25090), .I1(n25091), .I2(n25092), .I3(n25093), .S0(
        n26258), .S1(n26376), .ZN(n25089) );
  MUX41 U11520 ( .I0(ram[8990]), .I1(ram[8982]), .I2(ram[8974]), .I3(
        ram[8966]), .S0(n27281), .S1(n26806), .ZN(n25093) );
  MUX41 U11521 ( .I0(ram[9022]), .I1(ram[9014]), .I2(ram[9006]), .I3(
        ram[8998]), .S0(n27281), .S1(n26806), .ZN(n25091) );
  MUX41 U11522 ( .I0(ram[9086]), .I1(ram[9078]), .I2(ram[9070]), .I3(
        ram[9062]), .S0(n27282), .S1(n26807), .ZN(n25090) );
  MUX41 U11523 ( .I0(n26050), .I1(n26051), .I2(n26052), .I3(n26053), .S0(
        n26272), .S1(n26390), .ZN(n26049) );
  MUX41 U11524 ( .I0(ram[15647]), .I1(ram[15639]), .I2(ram[15631]), .I3(
        ram[15623]), .S0(n27337), .S1(n26862), .ZN(n26053) );
  MUX41 U11525 ( .I0(ram[15679]), .I1(ram[15671]), .I2(ram[15663]), .I3(
        ram[15655]), .S0(n27337), .S1(n26862), .ZN(n26051) );
  MUX41 U11526 ( .I0(ram[15743]), .I1(ram[15735]), .I2(ram[15727]), .I3(
        ram[15719]), .S0(n27337), .S1(n26862), .ZN(n26050) );
  MUX41 U11527 ( .I0(n26070), .I1(n26071), .I2(n26072), .I3(n26073), .S0(
        n26272), .S1(n26390), .ZN(n26069) );
  MUX41 U11528 ( .I0(ram[16159]), .I1(ram[16151]), .I2(ram[16143]), .I3(
        ram[16135]), .S0(n27338), .S1(n26863), .ZN(n26073) );
  MUX41 U11529 ( .I0(ram[16191]), .I1(ram[16183]), .I2(ram[16175]), .I3(
        ram[16167]), .S0(n27338), .S1(n26863), .ZN(n26071) );
  MUX41 U11530 ( .I0(ram[16255]), .I1(ram[16247]), .I2(ram[16239]), .I3(
        ram[16231]), .S0(n27338), .S1(n26863), .ZN(n26070) );
  MUX41 U11531 ( .I0(n26030), .I1(n26031), .I2(n26032), .I3(n26033), .S0(
        n26272), .S1(n26390), .ZN(n26029) );
  MUX41 U11532 ( .I0(ram[15135]), .I1(ram[15127]), .I2(ram[15119]), .I3(
        ram[15111]), .S0(n27335), .S1(n26860), .ZN(n26033) );
  MUX41 U11533 ( .I0(ram[15167]), .I1(ram[15159]), .I2(ram[15151]), .I3(
        ram[15143]), .S0(n27336), .S1(n26861), .ZN(n26031) );
  MUX41 U11534 ( .I0(ram[15231]), .I1(ram[15223]), .I2(ram[15215]), .I3(
        ram[15207]), .S0(n27336), .S1(n26861), .ZN(n26030) );
  MUX41 U11535 ( .I0(n26010), .I1(n26011), .I2(n26012), .I3(n26013), .S0(
        n26271), .S1(n26389), .ZN(n26009) );
  MUX41 U11536 ( .I0(ram[14623]), .I1(ram[14615]), .I2(ram[14607]), .I3(
        ram[14599]), .S0(n27334), .S1(n26859), .ZN(n26013) );
  MUX41 U11537 ( .I0(ram[14655]), .I1(ram[14647]), .I2(ram[14639]), .I3(
        ram[14631]), .S0(n27334), .S1(n26859), .ZN(n26011) );
  MUX41 U11538 ( .I0(ram[14719]), .I1(ram[14711]), .I2(ram[14703]), .I3(
        ram[14695]), .S0(n27334), .S1(n26859), .ZN(n26010) );
  MUX41 U11539 ( .I0(n25965), .I1(n25966), .I2(n25967), .I3(n25968), .S0(
        n26271), .S1(n26389), .ZN(n25964) );
  MUX41 U11540 ( .I0(ram[13599]), .I1(ram[13591]), .I2(ram[13583]), .I3(
        ram[13575]), .S0(n27332), .S1(n26857), .ZN(n25968) );
  MUX41 U11541 ( .I0(ram[13631]), .I1(ram[13623]), .I2(ram[13615]), .I3(
        ram[13607]), .S0(n27332), .S1(n26857), .ZN(n25966) );
  MUX41 U11542 ( .I0(ram[13695]), .I1(ram[13687]), .I2(ram[13679]), .I3(
        ram[13671]), .S0(n27332), .S1(n26857), .ZN(n25965) );
  MUX41 U11543 ( .I0(n25985), .I1(n25986), .I2(n25987), .I3(n25988), .S0(
        n26271), .S1(n26389), .ZN(n25984) );
  MUX41 U11544 ( .I0(ram[14111]), .I1(ram[14103]), .I2(ram[14095]), .I3(
        ram[14087]), .S0(n27333), .S1(n26858), .ZN(n25988) );
  MUX41 U11545 ( .I0(ram[14143]), .I1(ram[14135]), .I2(ram[14127]), .I3(
        ram[14119]), .S0(n27333), .S1(n26858), .ZN(n25986) );
  MUX41 U11546 ( .I0(ram[14207]), .I1(ram[14199]), .I2(ram[14191]), .I3(
        ram[14183]), .S0(n27333), .S1(n26858), .ZN(n25985) );
  MUX41 U11547 ( .I0(n25945), .I1(n25946), .I2(n25947), .I3(n25948), .S0(
        n26271), .S1(n26389), .ZN(n25944) );
  MUX41 U11548 ( .I0(ram[13087]), .I1(ram[13079]), .I2(ram[13071]), .I3(
        ram[13063]), .S0(n27331), .S1(n26856), .ZN(n25948) );
  MUX41 U11549 ( .I0(ram[13119]), .I1(ram[13111]), .I2(ram[13103]), .I3(
        ram[13095]), .S0(n27331), .S1(n26856), .ZN(n25946) );
  MUX41 U11550 ( .I0(ram[13183]), .I1(ram[13175]), .I2(ram[13167]), .I3(
        ram[13159]), .S0(n27331), .S1(n26856), .ZN(n25945) );
  MUX41 U11551 ( .I0(n25925), .I1(n25926), .I2(n25927), .I3(n25928), .S0(
        n26270), .S1(n26388), .ZN(n25924) );
  MUX41 U11552 ( .I0(ram[12575]), .I1(ram[12567]), .I2(ram[12559]), .I3(
        ram[12551]), .S0(n27329), .S1(n26854), .ZN(n25928) );
  MUX41 U11553 ( .I0(ram[12607]), .I1(ram[12599]), .I2(ram[12591]), .I3(
        ram[12583]), .S0(n27329), .S1(n26854), .ZN(n25926) );
  MUX41 U11554 ( .I0(ram[12671]), .I1(ram[12663]), .I2(ram[12655]), .I3(
        ram[12647]), .S0(n27330), .S1(n26855), .ZN(n25925) );
  MUX41 U11555 ( .I0(n25708), .I1(n25709), .I2(n25710), .I3(n25711), .S0(
        n26267), .S1(n26385), .ZN(n25707) );
  MUX41 U11556 ( .I0(ram[7487]), .I1(ram[7479]), .I2(ram[7471]), .I3(
        ram[7463]), .S0(n27317), .S1(n26842), .ZN(n25709) );
  MUX41 U11557 ( .I0(ram[7455]), .I1(ram[7447]), .I2(ram[7439]), .I3(
        ram[7431]), .S0(n27317), .S1(n26842), .ZN(n25711) );
  MUX41 U11558 ( .I0(ram[7551]), .I1(ram[7543]), .I2(ram[7535]), .I3(
        ram[7527]), .S0(n27317), .S1(n26842), .ZN(n25708) );
  MUX41 U11559 ( .I0(n25728), .I1(n25729), .I2(n25730), .I3(n25731), .S0(
        n26267), .S1(n26385), .ZN(n25727) );
  MUX41 U11560 ( .I0(ram[7967]), .I1(ram[7959]), .I2(ram[7951]), .I3(
        ram[7943]), .S0(n27318), .S1(n26843), .ZN(n25731) );
  MUX41 U11561 ( .I0(ram[7999]), .I1(ram[7991]), .I2(ram[7983]), .I3(
        ram[7975]), .S0(n27318), .S1(n26843), .ZN(n25729) );
  MUX41 U11562 ( .I0(ram[8063]), .I1(ram[8055]), .I2(ram[8047]), .I3(
        ram[8039]), .S0(n27318), .S1(n26843), .ZN(n25728) );
  MUX41 U11563 ( .I0(n25668), .I1(n25669), .I2(n25670), .I3(n25671), .S0(
        n26267), .S1(n26385), .ZN(n25667) );
  MUX41 U11564 ( .I0(ram[6431]), .I1(ram[6423]), .I2(ram[6415]), .I3(
        ram[6407]), .S0(n27315), .S1(n26840), .ZN(n25671) );
  MUX41 U11565 ( .I0(ram[6463]), .I1(ram[6455]), .I2(ram[6447]), .I3(
        ram[6439]), .S0(n27315), .S1(n26840), .ZN(n25669) );
  MUX41 U11566 ( .I0(ram[6527]), .I1(ram[6519]), .I2(ram[6511]), .I3(
        ram[6503]), .S0(n27315), .S1(n26840), .ZN(n25668) );
  MUX41 U11567 ( .I0(n25688), .I1(n25689), .I2(n25690), .I3(n25691), .S0(
        n26267), .S1(n26385), .ZN(n25687) );
  MUX41 U11568 ( .I0(ram[6943]), .I1(ram[6935]), .I2(ram[6927]), .I3(
        ram[6919]), .S0(n27316), .S1(n26841), .ZN(n25691) );
  MUX41 U11569 ( .I0(ram[6975]), .I1(ram[6967]), .I2(ram[6959]), .I3(
        ram[6951]), .S0(n27316), .S1(n26841), .ZN(n25689) );
  MUX41 U11570 ( .I0(ram[7039]), .I1(ram[7031]), .I2(ram[7023]), .I3(
        ram[7015]), .S0(n27316), .S1(n26841), .ZN(n25688) );
  MUX41 U11571 ( .I0(n25623), .I1(n25624), .I2(n25625), .I3(n25626), .S0(
        n26266), .S1(n26384), .ZN(n25622) );
  MUX41 U11572 ( .I0(ram[5439]), .I1(ram[5431]), .I2(ram[5423]), .I3(
        ram[5415]), .S0(n27312), .S1(n26837), .ZN(n25624) );
  MUX41 U11573 ( .I0(ram[5407]), .I1(ram[5399]), .I2(ram[5391]), .I3(
        ram[5383]), .S0(n27312), .S1(n26837), .ZN(n25626) );
  MUX41 U11574 ( .I0(ram[5503]), .I1(ram[5495]), .I2(ram[5487]), .I3(
        ram[5479]), .S0(n27312), .S1(n26837), .ZN(n25623) );
  MUX41 U11575 ( .I0(n25643), .I1(n25644), .I2(n25645), .I3(n25646), .S0(
        n26266), .S1(n26384), .ZN(n25642) );
  MUX41 U11576 ( .I0(ram[5951]), .I1(ram[5943]), .I2(ram[5935]), .I3(
        ram[5927]), .S0(n27313), .S1(n26838), .ZN(n25644) );
  MUX41 U11577 ( .I0(ram[5919]), .I1(ram[5911]), .I2(ram[5903]), .I3(
        ram[5895]), .S0(n27313), .S1(n26838), .ZN(n25646) );
  MUX41 U11578 ( .I0(ram[6015]), .I1(ram[6007]), .I2(ram[5999]), .I3(
        ram[5991]), .S0(n27314), .S1(n26839), .ZN(n25643) );
  MUX41 U11579 ( .I0(n25583), .I1(n25584), .I2(n25585), .I3(n25586), .S0(
        n26265), .S1(n26383), .ZN(n25582) );
  MUX41 U11580 ( .I0(ram[4415]), .I1(ram[4407]), .I2(ram[4399]), .I3(
        ram[4391]), .S0(n27310), .S1(n26835), .ZN(n25584) );
  MUX41 U11581 ( .I0(ram[4383]), .I1(ram[4375]), .I2(ram[4367]), .I3(
        ram[4359]), .S0(n27310), .S1(n26835), .ZN(n25586) );
  MUX41 U11582 ( .I0(ram[4479]), .I1(ram[4471]), .I2(ram[4463]), .I3(
        ram[4455]), .S0(n27310), .S1(n26835), .ZN(n25583) );
  MUX41 U11583 ( .I0(n25603), .I1(n25604), .I2(n25605), .I3(n25606), .S0(
        n26266), .S1(n26384), .ZN(n25602) );
  MUX41 U11584 ( .I0(ram[4895]), .I1(ram[4887]), .I2(ram[4879]), .I3(
        ram[4871]), .S0(n27311), .S1(n26836), .ZN(n25606) );
  MUX41 U11585 ( .I0(ram[4927]), .I1(ram[4919]), .I2(ram[4911]), .I3(
        ram[4903]), .S0(n27311), .S1(n26836), .ZN(n25604) );
  MUX41 U11586 ( .I0(ram[4991]), .I1(ram[4983]), .I2(ram[4975]), .I3(
        ram[4967]), .S0(n27311), .S1(n26836), .ZN(n25603) );
  MUX41 U11587 ( .I0(n25879), .I1(n25880), .I2(n25881), .I3(n25882), .S0(
        n26270), .S1(n26388), .ZN(n25878) );
  MUX41 U11588 ( .I0(ram[11583]), .I1(ram[11575]), .I2(ram[11567]), .I3(
        ram[11559]), .S0(n27327), .S1(n26852), .ZN(n25880) );
  MUX41 U11589 ( .I0(ram[11551]), .I1(ram[11543]), .I2(ram[11535]), .I3(
        ram[11527]), .S0(n27327), .S1(n26852), .ZN(n25882) );
  MUX41 U11590 ( .I0(ram[11647]), .I1(ram[11639]), .I2(ram[11631]), .I3(
        ram[11623]), .S0(n27327), .S1(n26852), .ZN(n25879) );
  MUX41 U11591 ( .I0(n25899), .I1(n25900), .I2(n25901), .I3(n25902), .S0(
        n26270), .S1(n26388), .ZN(n25898) );
  MUX41 U11592 ( .I0(ram[12095]), .I1(ram[12087]), .I2(ram[12079]), .I3(
        ram[12071]), .S0(n27328), .S1(n26853), .ZN(n25900) );
  MUX41 U11593 ( .I0(ram[12063]), .I1(ram[12055]), .I2(ram[12047]), .I3(
        ram[12039]), .S0(n27328), .S1(n26853), .ZN(n25902) );
  MUX41 U11594 ( .I0(ram[12159]), .I1(ram[12151]), .I2(ram[12143]), .I3(
        ram[12135]), .S0(n27328), .S1(n26853), .ZN(n25899) );
  MUX41 U11595 ( .I0(n25839), .I1(n25840), .I2(n25841), .I3(n25842), .S0(
        n26269), .S1(n26387), .ZN(n25838) );
  MUX41 U11596 ( .I0(ram[10559]), .I1(ram[10551]), .I2(ram[10543]), .I3(
        ram[10535]), .S0(n27324), .S1(n26849), .ZN(n25840) );
  MUX41 U11597 ( .I0(ram[10527]), .I1(ram[10519]), .I2(ram[10511]), .I3(
        ram[10503]), .S0(n27324), .S1(n26849), .ZN(n25842) );
  MUX41 U11598 ( .I0(ram[10623]), .I1(ram[10615]), .I2(ram[10607]), .I3(
        ram[10599]), .S0(n27325), .S1(n26850), .ZN(n25839) );
  MUX41 U11599 ( .I0(n25859), .I1(n25860), .I2(n25861), .I3(n25862), .S0(
        n26269), .S1(n26387), .ZN(n25858) );
  MUX41 U11600 ( .I0(ram[11039]), .I1(ram[11031]), .I2(ram[11023]), .I3(
        ram[11015]), .S0(n27326), .S1(n26851), .ZN(n25862) );
  MUX41 U11601 ( .I0(ram[11071]), .I1(ram[11063]), .I2(ram[11055]), .I3(
        ram[11047]), .S0(n27326), .S1(n26851), .ZN(n25860) );
  MUX41 U11602 ( .I0(ram[11135]), .I1(ram[11127]), .I2(ram[11119]), .I3(
        ram[11111]), .S0(n27326), .S1(n26851), .ZN(n25859) );
  MUX41 U11603 ( .I0(n25794), .I1(n25795), .I2(n25796), .I3(n25797), .S0(
        n26268), .S1(n26386), .ZN(n25793) );
  MUX41 U11604 ( .I0(ram[9535]), .I1(ram[9527]), .I2(ram[9519]), .I3(
        ram[9511]), .S0(n27322), .S1(n26847), .ZN(n25795) );
  MUX41 U11605 ( .I0(ram[9503]), .I1(ram[9495]), .I2(ram[9487]), .I3(
        ram[9479]), .S0(n27322), .S1(n26847), .ZN(n25797) );
  MUX41 U11606 ( .I0(ram[9599]), .I1(ram[9591]), .I2(ram[9583]), .I3(
        ram[9575]), .S0(n27322), .S1(n26847), .ZN(n25794) );
  MUX41 U11607 ( .I0(n25814), .I1(n25815), .I2(n25816), .I3(n25817), .S0(
        n26269), .S1(n26387), .ZN(n25813) );
  MUX41 U11608 ( .I0(ram[10047]), .I1(ram[10039]), .I2(ram[10031]), .I3(
        ram[10023]), .S0(n27323), .S1(n26848), .ZN(n25815) );
  MUX41 U11609 ( .I0(ram[10015]), .I1(ram[10007]), .I2(ram[9999]), .I3(
        ram[9991]), .S0(n27323), .S1(n26848), .ZN(n25817) );
  MUX41 U11610 ( .I0(ram[10111]), .I1(ram[10103]), .I2(ram[10095]), .I3(
        ram[10087]), .S0(n27323), .S1(n26848), .ZN(n25814) );
  MUX41 U11611 ( .I0(n25754), .I1(n25755), .I2(n25756), .I3(n25757), .S0(
        n26268), .S1(n26386), .ZN(n25753) );
  MUX41 U11612 ( .I0(ram[8511]), .I1(ram[8503]), .I2(ram[8495]), .I3(
        ram[8487]), .S0(n27320), .S1(n26845), .ZN(n25755) );
  MUX41 U11613 ( .I0(ram[8479]), .I1(ram[8471]), .I2(ram[8463]), .I3(
        ram[8455]), .S0(n27319), .S1(n26844), .ZN(n25757) );
  MUX41 U11614 ( .I0(ram[8575]), .I1(ram[8567]), .I2(ram[8559]), .I3(
        ram[8551]), .S0(n27320), .S1(n26845), .ZN(n25754) );
  MUX41 U11615 ( .I0(n25774), .I1(n25775), .I2(n25776), .I3(n25777), .S0(
        n26268), .S1(n26386), .ZN(n25773) );
  MUX41 U11616 ( .I0(ram[8991]), .I1(ram[8983]), .I2(ram[8975]), .I3(
        ram[8967]), .S0(n27321), .S1(n26846), .ZN(n25777) );
  MUX41 U11617 ( .I0(ram[9023]), .I1(ram[9015]), .I2(ram[9007]), .I3(
        ram[8999]), .S0(n27321), .S1(n26846), .ZN(n25775) );
  MUX41 U11618 ( .I0(ram[9087]), .I1(ram[9079]), .I2(ram[9071]), .I3(
        ram[9063]), .S0(n27321), .S1(n26846), .ZN(n25774) );
  MUX41 U11619 ( .I0(n20649), .I1(n20650), .I2(n20651), .I3(n20652), .S0(
        n26194), .S1(n26312), .ZN(n20648) );
  MUX41 U11620 ( .I0(ram[920]), .I1(ram[912]), .I2(ram[904]), .I3(
        ram[896]), .S0(n27026), .S1(n26551), .ZN(n20652) );
  MUX41 U11621 ( .I0(ram[952]), .I1(ram[944]), .I2(ram[936]), .I3(
        ram[928]), .S0(n27026), .S1(n26551), .ZN(n20650) );
  MUX41 U11622 ( .I0(ram[1016]), .I1(ram[1008]), .I2(ram[1000]), .I3(
        ram[992]), .S0(n27026), .S1(n26551), .ZN(n20649) );
  MUX41 U11623 ( .I0(ram[3576]), .I1(ram[3568]), .I2(ram[3560]), .I3(
        ram[3552]), .S0(n27032), .S1(n26557), .ZN(n20754) );
  MUX41 U11624 ( .I0(ram[3320]), .I1(ram[3312]), .I2(ram[3304]), .I3(
        ram[3296]), .S0(n27031), .S1(n26556), .ZN(n20744) );
  MUX41 U11625 ( .I0(ram[3192]), .I1(ram[3184]), .I2(ram[3176]), .I3(
        ram[3168]), .S0(n27031), .S1(n26556), .ZN(n20739) );
  MUX41 U11626 ( .I0(ram[4088]), .I1(ram[4080]), .I2(ram[4072]), .I3(
        ram[4064]), .S0(n27033), .S1(n26558), .ZN(n20774) );
  MUX41 U11627 ( .I0(ram[3832]), .I1(ram[3824]), .I2(ram[3816]), .I3(
        ram[3808]), .S0(n27033), .S1(n26558), .ZN(n20764) );
  MUX41 U11628 ( .I0(ram[3704]), .I1(ram[3696]), .I2(ram[3688]), .I3(
        ram[3680]), .S0(n27032), .S1(n26557), .ZN(n20759) );
  MUX41 U11629 ( .I0(ram[2552]), .I1(ram[2544]), .I2(ram[2536]), .I3(
        ram[2528]), .S0(n27030), .S1(n26555), .ZN(n20714) );
  MUX41 U11630 ( .I0(ram[1528]), .I1(ram[1520]), .I2(ram[1512]), .I3(
        ram[1504]), .S0(n27027), .S1(n26552), .ZN(n20669) );
  MUX41 U11631 ( .I0(ram[1272]), .I1(ram[1264]), .I2(ram[1256]), .I3(
        ram[1248]), .S0(n27026), .S1(n26551), .ZN(n20659) );
  MUX41 U11632 ( .I0(ram[1144]), .I1(ram[1136]), .I2(ram[1128]), .I3(
        ram[1120]), .S0(n27026), .S1(n26551), .ZN(n20654) );
  MUX41 U11633 ( .I0(ram[2040]), .I1(ram[2032]), .I2(ram[2024]), .I3(
        ram[2016]), .S0(n27028), .S1(n26553), .ZN(n20689) );
  MUX41 U11634 ( .I0(ram[1784]), .I1(ram[1776]), .I2(ram[1768]), .I3(
        ram[1760]), .S0(n27028), .S1(n26553), .ZN(n20679) );
  MUX41 U11635 ( .I0(ram[1656]), .I1(ram[1648]), .I2(ram[1640]), .I3(
        ram[1632]), .S0(n27027), .S1(n26552), .ZN(n20674) );
  MUX41 U11636 ( .I0(ram[3577]), .I1(ram[3569]), .I2(ram[3561]), .I3(
        ram[3553]), .S0(n27071), .S1(n26596), .ZN(n21438) );
  MUX41 U11637 ( .I0(ram[3321]), .I1(ram[3313]), .I2(ram[3305]), .I3(
        ram[3297]), .S0(n27071), .S1(n26596), .ZN(n21428) );
  MUX41 U11638 ( .I0(ram[3193]), .I1(ram[3185]), .I2(ram[3177]), .I3(
        ram[3169]), .S0(n27070), .S1(n26595), .ZN(n21423) );
  MUX41 U11639 ( .I0(ram[4089]), .I1(ram[4081]), .I2(ram[4073]), .I3(
        ram[4065]), .S0(n27073), .S1(n26598), .ZN(n21458) );
  MUX41 U11640 ( .I0(ram[3833]), .I1(ram[3825]), .I2(ram[3817]), .I3(
        ram[3809]), .S0(n27072), .S1(n26597), .ZN(n21448) );
  MUX41 U11641 ( .I0(ram[3705]), .I1(ram[3697]), .I2(ram[3689]), .I3(
        ram[3681]), .S0(n27072), .S1(n26597), .ZN(n21443) );
  MUX41 U11642 ( .I0(ram[2553]), .I1(ram[2545]), .I2(ram[2537]), .I3(
        ram[2529]), .S0(n27069), .S1(n26594), .ZN(n21398) );
  MUX41 U11643 ( .I0(ram[1529]), .I1(ram[1521]), .I2(ram[1513]), .I3(
        ram[1505]), .S0(n27066), .S1(n26591), .ZN(n21353) );
  MUX41 U11644 ( .I0(ram[1273]), .I1(ram[1265]), .I2(ram[1257]), .I3(
        ram[1249]), .S0(n27066), .S1(n26591), .ZN(n21343) );
  MUX41 U11645 ( .I0(ram[1145]), .I1(ram[1137]), .I2(ram[1129]), .I3(
        ram[1121]), .S0(n27066), .S1(n26591), .ZN(n21338) );
  MUX41 U11646 ( .I0(ram[2041]), .I1(ram[2033]), .I2(ram[2025]), .I3(
        ram[2017]), .S0(n27068), .S1(n26593), .ZN(n21373) );
  MUX41 U11647 ( .I0(ram[1785]), .I1(ram[1777]), .I2(ram[1769]), .I3(
        ram[1761]), .S0(n27067), .S1(n26592), .ZN(n21363) );
  MUX41 U11648 ( .I0(ram[1657]), .I1(ram[1649]), .I2(ram[1641]), .I3(
        ram[1633]), .S0(n27067), .S1(n26592), .ZN(n21358) );
  MUX41 U11649 ( .I0(ram[505]), .I1(ram[497]), .I2(ram[489]), .I3(
        ram[481]), .S0(n27064), .S1(n26589), .ZN(n21313) );
  MUX41 U11650 ( .I0(ram[3578]), .I1(ram[3570]), .I2(ram[3562]), .I3(
        ram[3554]), .S0(n27111), .S1(n26636), .ZN(n22122) );
  MUX41 U11651 ( .I0(ram[3322]), .I1(ram[3314]), .I2(ram[3306]), .I3(
        ram[3298]), .S0(n27110), .S1(n26635), .ZN(n22112) );
  MUX41 U11652 ( .I0(ram[3194]), .I1(ram[3186]), .I2(ram[3178]), .I3(
        ram[3170]), .S0(n27110), .S1(n26635), .ZN(n22107) );
  MUX41 U11653 ( .I0(ram[4090]), .I1(ram[4082]), .I2(ram[4074]), .I3(
        ram[4066]), .S0(n27112), .S1(n26637), .ZN(n22142) );
  MUX41 U11654 ( .I0(ram[3834]), .I1(ram[3826]), .I2(ram[3818]), .I3(
        ram[3810]), .S0(n27111), .S1(n26636), .ZN(n22132) );
  MUX41 U11655 ( .I0(ram[3706]), .I1(ram[3698]), .I2(ram[3690]), .I3(
        ram[3682]), .S0(n27111), .S1(n26636), .ZN(n22127) );
  MUX41 U11656 ( .I0(ram[2554]), .I1(ram[2546]), .I2(ram[2538]), .I3(
        ram[2530]), .S0(n27108), .S1(n26633), .ZN(n22082) );
  MUX41 U11657 ( .I0(ram[1530]), .I1(ram[1522]), .I2(ram[1514]), .I3(
        ram[1506]), .S0(n27106), .S1(n26631), .ZN(n22037) );
  MUX41 U11658 ( .I0(ram[1274]), .I1(ram[1266]), .I2(ram[1258]), .I3(
        ram[1250]), .S0(n27105), .S1(n26630), .ZN(n22027) );
  MUX41 U11659 ( .I0(ram[1146]), .I1(ram[1138]), .I2(ram[1130]), .I3(
        ram[1122]), .S0(n27105), .S1(n26630), .ZN(n22022) );
  MUX41 U11660 ( .I0(ram[2042]), .I1(ram[2034]), .I2(ram[2026]), .I3(
        ram[2018]), .S0(n27107), .S1(n26632), .ZN(n22057) );
  MUX41 U11661 ( .I0(ram[1786]), .I1(ram[1778]), .I2(ram[1770]), .I3(
        ram[1762]), .S0(n27106), .S1(n26631), .ZN(n22047) );
  MUX41 U11662 ( .I0(ram[1658]), .I1(ram[1650]), .I2(ram[1642]), .I3(
        ram[1634]), .S0(n27106), .S1(n26631), .ZN(n22042) );
  MUX41 U11663 ( .I0(ram[506]), .I1(ram[498]), .I2(ram[490]), .I3(
        ram[482]), .S0(n27103), .S1(n26628), .ZN(n21997) );
  MUX41 U11664 ( .I0(ram[3579]), .I1(ram[3571]), .I2(ram[3563]), .I3(
        ram[3555]), .S0(n27150), .S1(n26675), .ZN(n22806) );
  MUX41 U11665 ( .I0(ram[3323]), .I1(ram[3315]), .I2(ram[3307]), .I3(
        ram[3299]), .S0(n27150), .S1(n26675), .ZN(n22796) );
  MUX41 U11666 ( .I0(ram[3195]), .I1(ram[3187]), .I2(ram[3179]), .I3(
        ram[3171]), .S0(n27149), .S1(n26674), .ZN(n22791) );
  MUX41 U11667 ( .I0(ram[4091]), .I1(ram[4083]), .I2(ram[4075]), .I3(
        ram[4067]), .S0(n27151), .S1(n26676), .ZN(n22826) );
  MUX41 U11668 ( .I0(ram[3835]), .I1(ram[3827]), .I2(ram[3819]), .I3(
        ram[3811]), .S0(n27151), .S1(n26676), .ZN(n22816) );
  MUX41 U11669 ( .I0(ram[3707]), .I1(ram[3699]), .I2(ram[3691]), .I3(
        ram[3683]), .S0(n27150), .S1(n26675), .ZN(n22811) );
  MUX41 U11670 ( .I0(ram[2555]), .I1(ram[2547]), .I2(ram[2539]), .I3(
        ram[2531]), .S0(n27148), .S1(n26673), .ZN(n22766) );
  MUX41 U11671 ( .I0(ram[1531]), .I1(ram[1523]), .I2(ram[1515]), .I3(
        ram[1507]), .S0(n27145), .S1(n26670), .ZN(n22721) );
  MUX41 U11672 ( .I0(ram[1275]), .I1(ram[1267]), .I2(ram[1259]), .I3(
        ram[1251]), .S0(n27145), .S1(n26670), .ZN(n22711) );
  MUX41 U11673 ( .I0(ram[1147]), .I1(ram[1139]), .I2(ram[1131]), .I3(
        ram[1123]), .S0(n27144), .S1(n26669), .ZN(n22706) );
  MUX41 U11674 ( .I0(ram[2043]), .I1(ram[2035]), .I2(ram[2027]), .I3(
        ram[2019]), .S0(n27146), .S1(n26671), .ZN(n22741) );
  MUX41 U11675 ( .I0(ram[1787]), .I1(ram[1779]), .I2(ram[1771]), .I3(
        ram[1763]), .S0(n27146), .S1(n26671), .ZN(n22731) );
  MUX41 U11676 ( .I0(ram[1659]), .I1(ram[1651]), .I2(ram[1643]), .I3(
        ram[1635]), .S0(n27146), .S1(n26671), .ZN(n22726) );
  MUX41 U11677 ( .I0(ram[507]), .I1(ram[499]), .I2(ram[491]), .I3(
        ram[483]), .S0(n27143), .S1(n26668), .ZN(n22681) );
  MUX41 U11678 ( .I0(ram[3580]), .I1(ram[3572]), .I2(ram[3564]), .I3(
        ram[3556]), .S0(n27190), .S1(n26715), .ZN(n23490) );
  MUX41 U11679 ( .I0(ram[3324]), .I1(ram[3316]), .I2(ram[3308]), .I3(
        ram[3300]), .S0(n27189), .S1(n26714), .ZN(n23480) );
  MUX41 U11680 ( .I0(ram[3196]), .I1(ram[3188]), .I2(ram[3180]), .I3(
        ram[3172]), .S0(n27189), .S1(n26714), .ZN(n23475) );
  MUX41 U11681 ( .I0(ram[4092]), .I1(ram[4084]), .I2(ram[4076]), .I3(
        ram[4068]), .S0(n27191), .S1(n26716), .ZN(n23510) );
  MUX41 U11682 ( .I0(ram[3836]), .I1(ram[3828]), .I2(ram[3820]), .I3(
        ram[3812]), .S0(n27190), .S1(n26715), .ZN(n23500) );
  MUX41 U11683 ( .I0(ram[3708]), .I1(ram[3700]), .I2(ram[3692]), .I3(
        ram[3684]), .S0(n27190), .S1(n26715), .ZN(n23495) );
  MUX41 U11684 ( .I0(ram[2556]), .I1(ram[2548]), .I2(ram[2540]), .I3(
        ram[2532]), .S0(n27187), .S1(n26712), .ZN(n23450) );
  MUX41 U11685 ( .I0(ram[1532]), .I1(ram[1524]), .I2(ram[1516]), .I3(
        ram[1508]), .S0(n27185), .S1(n26710), .ZN(n23405) );
  MUX41 U11686 ( .I0(ram[1276]), .I1(ram[1268]), .I2(ram[1260]), .I3(
        ram[1252]), .S0(n27184), .S1(n26709), .ZN(n23395) );
  MUX41 U11687 ( .I0(ram[1148]), .I1(ram[1140]), .I2(ram[1132]), .I3(
        ram[1124]), .S0(n27184), .S1(n26709), .ZN(n23390) );
  MUX41 U11688 ( .I0(ram[2044]), .I1(ram[2036]), .I2(ram[2028]), .I3(
        ram[2020]), .S0(n27186), .S1(n26711), .ZN(n23425) );
  MUX41 U11689 ( .I0(ram[1788]), .I1(ram[1780]), .I2(ram[1772]), .I3(
        ram[1764]), .S0(n27185), .S1(n26710), .ZN(n23415) );
  MUX41 U11690 ( .I0(ram[1660]), .I1(ram[1652]), .I2(ram[1644]), .I3(
        ram[1636]), .S0(n27185), .S1(n26710), .ZN(n23410) );
  MUX41 U11691 ( .I0(ram[508]), .I1(ram[500]), .I2(ram[492]), .I3(
        ram[484]), .S0(n27182), .S1(n26707), .ZN(n23365) );
  MUX41 U11692 ( .I0(ram[3581]), .I1(ram[3573]), .I2(ram[3565]), .I3(
        ram[3557]), .S0(n27229), .S1(n26754), .ZN(n24174) );
  MUX41 U11693 ( .I0(ram[3325]), .I1(ram[3317]), .I2(ram[3309]), .I3(
        ram[3301]), .S0(n27228), .S1(n26753), .ZN(n24164) );
  MUX41 U11694 ( .I0(ram[3197]), .I1(ram[3189]), .I2(ram[3181]), .I3(
        ram[3173]), .S0(n27228), .S1(n26753), .ZN(n24159) );
  MUX41 U11695 ( .I0(ram[4093]), .I1(ram[4085]), .I2(ram[4077]), .I3(
        ram[4069]), .S0(n27230), .S1(n26755), .ZN(n24194) );
  MUX41 U11696 ( .I0(ram[3837]), .I1(ram[3829]), .I2(ram[3821]), .I3(
        ram[3813]), .S0(n27230), .S1(n26755), .ZN(n24184) );
  MUX41 U11697 ( .I0(ram[3709]), .I1(ram[3701]), .I2(ram[3693]), .I3(
        ram[3685]), .S0(n27229), .S1(n26754), .ZN(n24179) );
  MUX41 U11698 ( .I0(ram[2557]), .I1(ram[2549]), .I2(ram[2541]), .I3(
        ram[2533]), .S0(n27226), .S1(n26751), .ZN(n24134) );
  MUX41 U11699 ( .I0(ram[1533]), .I1(ram[1525]), .I2(ram[1517]), .I3(
        ram[1509]), .S0(n27224), .S1(n26749), .ZN(n24089) );
  MUX41 U11700 ( .I0(ram[1277]), .I1(ram[1269]), .I2(ram[1261]), .I3(
        ram[1253]), .S0(n27223), .S1(n26748), .ZN(n24079) );
  MUX41 U11701 ( .I0(ram[1149]), .I1(ram[1141]), .I2(ram[1133]), .I3(
        ram[1125]), .S0(n27223), .S1(n26748), .ZN(n24074) );
  MUX41 U11702 ( .I0(ram[2045]), .I1(ram[2037]), .I2(ram[2029]), .I3(
        ram[2021]), .S0(n27225), .S1(n26750), .ZN(n24109) );
  MUX41 U11703 ( .I0(ram[1789]), .I1(ram[1781]), .I2(ram[1773]), .I3(
        ram[1765]), .S0(n27225), .S1(n26750), .ZN(n24099) );
  MUX41 U11704 ( .I0(ram[1661]), .I1(ram[1653]), .I2(ram[1645]), .I3(
        ram[1637]), .S0(n27224), .S1(n26749), .ZN(n24094) );
  MUX41 U11705 ( .I0(ram[509]), .I1(ram[501]), .I2(ram[493]), .I3(
        ram[485]), .S0(n27222), .S1(n26747), .ZN(n24049) );
  MUX41 U11706 ( .I0(ram[3582]), .I1(ram[3574]), .I2(ram[3566]), .I3(
        ram[3558]), .S0(n27268), .S1(n26793), .ZN(n24858) );
  MUX41 U11707 ( .I0(ram[3326]), .I1(ram[3318]), .I2(ram[3310]), .I3(
        ram[3302]), .S0(n27268), .S1(n26793), .ZN(n24848) );
  MUX41 U11708 ( .I0(ram[3198]), .I1(ram[3190]), .I2(ram[3182]), .I3(
        ram[3174]), .S0(n27267), .S1(n26792), .ZN(n24843) );
  MUX41 U11709 ( .I0(ram[4094]), .I1(ram[4086]), .I2(ram[4078]), .I3(
        ram[4070]), .S0(n27270), .S1(n26795), .ZN(n24878) );
  MUX41 U11710 ( .I0(ram[3838]), .I1(ram[3830]), .I2(ram[3822]), .I3(
        ram[3814]), .S0(n27269), .S1(n26794), .ZN(n24868) );
  MUX41 U11711 ( .I0(ram[3710]), .I1(ram[3702]), .I2(ram[3694]), .I3(
        ram[3686]), .S0(n27269), .S1(n26794), .ZN(n24863) );
  MUX41 U11712 ( .I0(ram[2558]), .I1(ram[2550]), .I2(ram[2542]), .I3(
        ram[2534]), .S0(n27266), .S1(n26791), .ZN(n24818) );
  MUX41 U11713 ( .I0(ram[1534]), .I1(ram[1526]), .I2(ram[1518]), .I3(
        ram[1510]), .S0(n27263), .S1(n26788), .ZN(n24773) );
  MUX41 U11714 ( .I0(ram[1278]), .I1(ram[1270]), .I2(ram[1262]), .I3(
        ram[1254]), .S0(n27263), .S1(n26788), .ZN(n24763) );
  MUX41 U11715 ( .I0(ram[1150]), .I1(ram[1142]), .I2(ram[1134]), .I3(
        ram[1126]), .S0(n27262), .S1(n26787), .ZN(n24758) );
  MUX41 U11716 ( .I0(ram[2046]), .I1(ram[2038]), .I2(ram[2030]), .I3(
        ram[2022]), .S0(n27265), .S1(n26790), .ZN(n24793) );
  MUX41 U11717 ( .I0(ram[1790]), .I1(ram[1782]), .I2(ram[1774]), .I3(
        ram[1766]), .S0(n27264), .S1(n26789), .ZN(n24783) );
  MUX41 U11718 ( .I0(ram[1662]), .I1(ram[1654]), .I2(ram[1646]), .I3(
        ram[1638]), .S0(n27264), .S1(n26789), .ZN(n24778) );
  MUX41 U11719 ( .I0(ram[510]), .I1(ram[502]), .I2(ram[494]), .I3(
        ram[486]), .S0(n27261), .S1(n26786), .ZN(n24733) );
  MUX41 U11720 ( .I0(ram[3583]), .I1(ram[3575]), .I2(ram[3567]), .I3(
        ram[3559]), .S0(n27308), .S1(n26833), .ZN(n25542) );
  MUX41 U11721 ( .I0(ram[3327]), .I1(ram[3319]), .I2(ram[3311]), .I3(
        ram[3303]), .S0(n27307), .S1(n26832), .ZN(n25532) );
  MUX41 U11722 ( .I0(ram[3199]), .I1(ram[3191]), .I2(ram[3183]), .I3(
        ram[3175]), .S0(n27307), .S1(n26832), .ZN(n25527) );
  MUX41 U11723 ( .I0(ram[4095]), .I1(ram[4087]), .I2(ram[4079]), .I3(
        ram[4071]), .S0(n27309), .S1(n26834), .ZN(n25562) );
  MUX41 U11724 ( .I0(ram[3839]), .I1(ram[3831]), .I2(ram[3823]), .I3(
        ram[3815]), .S0(n27308), .S1(n26833), .ZN(n25552) );
  MUX41 U11725 ( .I0(ram[3711]), .I1(ram[3703]), .I2(ram[3695]), .I3(
        ram[3687]), .S0(n27308), .S1(n26833), .ZN(n25547) );
  MUX41 U11726 ( .I0(ram[2559]), .I1(ram[2551]), .I2(ram[2543]), .I3(
        ram[2535]), .S0(n27305), .S1(n26830), .ZN(n25502) );
  MUX41 U11727 ( .I0(ram[1535]), .I1(ram[1527]), .I2(ram[1519]), .I3(
        ram[1511]), .S0(n27303), .S1(n26828), .ZN(n25457) );
  MUX41 U11728 ( .I0(ram[1279]), .I1(ram[1271]), .I2(ram[1263]), .I3(
        ram[1255]), .S0(n27302), .S1(n26827), .ZN(n25447) );
  MUX41 U11729 ( .I0(ram[1151]), .I1(ram[1143]), .I2(ram[1135]), .I3(
        ram[1127]), .S0(n27302), .S1(n26827), .ZN(n25442) );
  MUX41 U11730 ( .I0(ram[2047]), .I1(ram[2039]), .I2(ram[2031]), .I3(
        ram[2023]), .S0(n27304), .S1(n26829), .ZN(n25477) );
  MUX41 U11731 ( .I0(ram[1791]), .I1(ram[1783]), .I2(ram[1775]), .I3(
        ram[1767]), .S0(n27303), .S1(n26828), .ZN(n25467) );
  MUX41 U11732 ( .I0(ram[1663]), .I1(ram[1655]), .I2(ram[1647]), .I3(
        ram[1639]), .S0(n27303), .S1(n26828), .ZN(n25462) );
  MUX41 U11733 ( .I0(ram[511]), .I1(ram[503]), .I2(ram[495]), .I3(
        ram[487]), .S0(n27300), .S1(n26825), .ZN(n25417) );
  MUX41 U11734 ( .I0(ram[15864]), .I1(ram[15856]), .I2(ram[15848]), .I3(
        ram[15840]), .S0(n27062), .S1(n26587), .ZN(n21267) );
  MUX41 U11735 ( .I0(ram[15608]), .I1(ram[15600]), .I2(ram[15592]), .I3(
        ram[15584]), .S0(n27061), .S1(n26586), .ZN(n21257) );
  MUX41 U11736 ( .I0(ram[15480]), .I1(ram[15472]), .I2(ram[15464]), .I3(
        ram[15456]), .S0(n27061), .S1(n26586), .ZN(n21252) );
  MUX41 U11737 ( .I0(ram[13816]), .I1(ram[13808]), .I2(ram[13800]), .I3(
        ram[13792]), .S0(n27057), .S1(n26582), .ZN(n21182) );
  MUX41 U11738 ( .I0(ram[13560]), .I1(ram[13552]), .I2(ram[13544]), .I3(
        ram[13536]), .S0(n27056), .S1(n26581), .ZN(n21172) );
  MUX41 U11739 ( .I0(ram[13432]), .I1(ram[13424]), .I2(ram[13416]), .I3(
        ram[13408]), .S0(n27056), .S1(n26581), .ZN(n21167) );
  MUX41 U11740 ( .I0(ram[7672]), .I1(ram[7664]), .I2(ram[7656]), .I3(
        ram[7648]), .S0(n27042), .S1(n26567), .ZN(n20925) );
  MUX41 U11741 ( .I0(ram[7416]), .I1(ram[7408]), .I2(ram[7400]), .I3(
        ram[7392]), .S0(n27041), .S1(n26566), .ZN(n20915) );
  MUX41 U11742 ( .I0(ram[7288]), .I1(ram[7280]), .I2(ram[7272]), .I3(
        ram[7264]), .S0(n27041), .S1(n26566), .ZN(n20910) );
  MUX41 U11743 ( .I0(ram[5624]), .I1(ram[5616]), .I2(ram[5608]), .I3(
        ram[5600]), .S0(n27037), .S1(n26562), .ZN(n20840) );
  MUX41 U11744 ( .I0(ram[5368]), .I1(ram[5360]), .I2(ram[5352]), .I3(
        ram[5344]), .S0(n27036), .S1(n26561), .ZN(n20830) );
  MUX41 U11745 ( .I0(ram[5240]), .I1(ram[5232]), .I2(ram[5224]), .I3(
        ram[5216]), .S0(n27036), .S1(n26561), .ZN(n20825) );
  MUX41 U11746 ( .I0(ram[11768]), .I1(ram[11760]), .I2(ram[11752]), .I3(
        ram[11744]), .S0(n27052), .S1(n26577), .ZN(n21096) );
  MUX41 U11747 ( .I0(ram[11512]), .I1(ram[11504]), .I2(ram[11496]), .I3(
        ram[11488]), .S0(n27051), .S1(n26576), .ZN(n21086) );
  MUX41 U11748 ( .I0(ram[11384]), .I1(ram[11376]), .I2(ram[11368]), .I3(
        ram[11360]), .S0(n27051), .S1(n26576), .ZN(n21081) );
  MUX41 U11749 ( .I0(ram[9720]), .I1(ram[9712]), .I2(ram[9704]), .I3(
        ram[9696]), .S0(n27047), .S1(n26572), .ZN(n21011) );
  MUX41 U11750 ( .I0(ram[9464]), .I1(ram[9456]), .I2(ram[9448]), .I3(
        ram[9440]), .S0(n27046), .S1(n26571), .ZN(n21001) );
  MUX41 U11751 ( .I0(ram[9336]), .I1(ram[9328]), .I2(ram[9320]), .I3(
        ram[9312]), .S0(n27046), .S1(n26571), .ZN(n20996) );
  MUX41 U11752 ( .I0(ram[15865]), .I1(ram[15857]), .I2(ram[15849]), .I3(
        ram[15841]), .S0(n27101), .S1(n26626), .ZN(n21951) );
  MUX41 U11753 ( .I0(ram[15609]), .I1(ram[15601]), .I2(ram[15593]), .I3(
        ram[15585]), .S0(n27100), .S1(n26625), .ZN(n21941) );
  MUX41 U11754 ( .I0(ram[15481]), .I1(ram[15473]), .I2(ram[15465]), .I3(
        ram[15457]), .S0(n27100), .S1(n26625), .ZN(n21936) );
  MUX41 U11755 ( .I0(ram[13817]), .I1(ram[13809]), .I2(ram[13801]), .I3(
        ram[13793]), .S0(n27096), .S1(n26621), .ZN(n21866) );
  MUX41 U11756 ( .I0(ram[13561]), .I1(ram[13553]), .I2(ram[13545]), .I3(
        ram[13537]), .S0(n27095), .S1(n26620), .ZN(n21856) );
  MUX41 U11757 ( .I0(ram[13433]), .I1(ram[13425]), .I2(ram[13417]), .I3(
        ram[13409]), .S0(n27095), .S1(n26620), .ZN(n21851) );
  MUX41 U11758 ( .I0(n21333), .I1(n21334), .I2(n21335), .I3(n21336), .S0(
        n26204), .S1(n26322), .ZN(n21332) );
  MUX41 U11759 ( .I0(ram[921]), .I1(ram[913]), .I2(ram[905]), .I3(
        ram[897]), .S0(n27065), .S1(n26590), .ZN(n21336) );
  MUX41 U11760 ( .I0(ram[953]), .I1(ram[945]), .I2(ram[937]), .I3(
        ram[929]), .S0(n27065), .S1(n26590), .ZN(n21334) );
  MUX41 U11761 ( .I0(ram[1017]), .I1(ram[1009]), .I2(ram[1001]), .I3(
        ram[993]), .S0(n27065), .S1(n26590), .ZN(n21333) );
  MUX41 U11762 ( .I0(ram[7673]), .I1(ram[7665]), .I2(ram[7657]), .I3(
        ram[7649]), .S0(n27081), .S1(n26606), .ZN(n21609) );
  MUX41 U11763 ( .I0(ram[7417]), .I1(ram[7409]), .I2(ram[7401]), .I3(
        ram[7393]), .S0(n27081), .S1(n26606), .ZN(n21599) );
  MUX41 U11764 ( .I0(ram[7289]), .I1(ram[7281]), .I2(ram[7273]), .I3(
        ram[7265]), .S0(n27080), .S1(n26605), .ZN(n21594) );
  MUX41 U11765 ( .I0(ram[5625]), .I1(ram[5617]), .I2(ram[5609]), .I3(
        ram[5601]), .S0(n27076), .S1(n26601), .ZN(n21524) );
  MUX41 U11766 ( .I0(ram[5369]), .I1(ram[5361]), .I2(ram[5353]), .I3(
        ram[5345]), .S0(n27076), .S1(n26601), .ZN(n21514) );
  MUX41 U11767 ( .I0(ram[5241]), .I1(ram[5233]), .I2(ram[5225]), .I3(
        ram[5217]), .S0(n27075), .S1(n26600), .ZN(n21509) );
  MUX41 U11768 ( .I0(ram[11769]), .I1(ram[11761]), .I2(ram[11753]), .I3(
        ram[11745]), .S0(n27091), .S1(n26616), .ZN(n21780) );
  MUX41 U11769 ( .I0(ram[11513]), .I1(ram[11505]), .I2(ram[11497]), .I3(
        ram[11489]), .S0(n27090), .S1(n26615), .ZN(n21770) );
  MUX41 U11770 ( .I0(ram[11385]), .I1(ram[11377]), .I2(ram[11369]), .I3(
        ram[11361]), .S0(n27090), .S1(n26615), .ZN(n21765) );
  MUX41 U11771 ( .I0(ram[9721]), .I1(ram[9713]), .I2(ram[9705]), .I3(
        ram[9697]), .S0(n27086), .S1(n26611), .ZN(n21695) );
  MUX41 U11772 ( .I0(ram[9465]), .I1(ram[9457]), .I2(ram[9449]), .I3(
        ram[9441]), .S0(n27086), .S1(n26611), .ZN(n21685) );
  MUX41 U11773 ( .I0(ram[9337]), .I1(ram[9329]), .I2(ram[9321]), .I3(
        ram[9313]), .S0(n27085), .S1(n26610), .ZN(n21680) );
  MUX41 U11774 ( .I0(ram[15866]), .I1(ram[15858]), .I2(ram[15850]), .I3(
        ram[15842]), .S0(n27140), .S1(n26665), .ZN(n22635) );
  MUX41 U11775 ( .I0(ram[15610]), .I1(ram[15602]), .I2(ram[15594]), .I3(
        ram[15586]), .S0(n27140), .S1(n26665), .ZN(n22625) );
  MUX41 U11776 ( .I0(ram[15482]), .I1(ram[15474]), .I2(ram[15466]), .I3(
        ram[15458]), .S0(n27139), .S1(n26664), .ZN(n22620) );
  MUX41 U11777 ( .I0(ram[13818]), .I1(ram[13810]), .I2(ram[13802]), .I3(
        ram[13794]), .S0(n27135), .S1(n26660), .ZN(n22550) );
  MUX41 U11778 ( .I0(ram[13562]), .I1(ram[13554]), .I2(ram[13546]), .I3(
        ram[13538]), .S0(n27135), .S1(n26660), .ZN(n22540) );
  MUX41 U11779 ( .I0(ram[13434]), .I1(ram[13426]), .I2(ram[13418]), .I3(
        ram[13410]), .S0(n27134), .S1(n26659), .ZN(n22535) );
  MUX41 U11780 ( .I0(n22017), .I1(n22018), .I2(n22019), .I3(n22020), .S0(
        n26214), .S1(n26332), .ZN(n22016) );
  MUX41 U11781 ( .I0(ram[922]), .I1(ram[914]), .I2(ram[906]), .I3(
        ram[898]), .S0(n27104), .S1(n26629), .ZN(n22020) );
  MUX41 U11782 ( .I0(ram[954]), .I1(ram[946]), .I2(ram[938]), .I3(
        ram[930]), .S0(n27104), .S1(n26629), .ZN(n22018) );
  MUX41 U11783 ( .I0(ram[1018]), .I1(ram[1010]), .I2(ram[1002]), .I3(
        ram[994]), .S0(n27105), .S1(n26630), .ZN(n22017) );
  MUX41 U11784 ( .I0(ram[7674]), .I1(ram[7666]), .I2(ram[7658]), .I3(
        ram[7650]), .S0(n27121), .S1(n26646), .ZN(n22293) );
  MUX41 U11785 ( .I0(ram[7418]), .I1(ram[7410]), .I2(ram[7402]), .I3(
        ram[7394]), .S0(n27120), .S1(n26645), .ZN(n22283) );
  MUX41 U11786 ( .I0(ram[7290]), .I1(ram[7282]), .I2(ram[7274]), .I3(
        ram[7266]), .S0(n27120), .S1(n26645), .ZN(n22278) );
  MUX41 U11787 ( .I0(ram[5626]), .I1(ram[5618]), .I2(ram[5610]), .I3(
        ram[5602]), .S0(n27116), .S1(n26641), .ZN(n22208) );
  MUX41 U11788 ( .I0(ram[5370]), .I1(ram[5362]), .I2(ram[5354]), .I3(
        ram[5346]), .S0(n27115), .S1(n26640), .ZN(n22198) );
  MUX41 U11789 ( .I0(ram[5242]), .I1(ram[5234]), .I2(ram[5226]), .I3(
        ram[5218]), .S0(n27115), .S1(n26640), .ZN(n22193) );
  MUX41 U11790 ( .I0(ram[11770]), .I1(ram[11762]), .I2(ram[11754]), .I3(
        ram[11746]), .S0(n27130), .S1(n26655), .ZN(n22464) );
  MUX41 U11791 ( .I0(ram[11514]), .I1(ram[11506]), .I2(ram[11498]), .I3(
        ram[11490]), .S0(n27130), .S1(n26655), .ZN(n22454) );
  MUX41 U11792 ( .I0(ram[11386]), .I1(ram[11378]), .I2(ram[11370]), .I3(
        ram[11362]), .S0(n27130), .S1(n26655), .ZN(n22449) );
  MUX41 U11793 ( .I0(ram[9722]), .I1(ram[9714]), .I2(ram[9706]), .I3(
        ram[9698]), .S0(n27126), .S1(n26651), .ZN(n22379) );
  MUX41 U11794 ( .I0(ram[9466]), .I1(ram[9458]), .I2(ram[9450]), .I3(
        ram[9442]), .S0(n27125), .S1(n26650), .ZN(n22369) );
  MUX41 U11795 ( .I0(ram[9338]), .I1(ram[9330]), .I2(ram[9322]), .I3(
        ram[9314]), .S0(n27125), .S1(n26650), .ZN(n22364) );
  MUX41 U11796 ( .I0(ram[15867]), .I1(ram[15859]), .I2(ram[15851]), .I3(
        ram[15843]), .S0(n27180), .S1(n26705), .ZN(n23319) );
  MUX41 U11797 ( .I0(ram[15611]), .I1(ram[15603]), .I2(ram[15595]), .I3(
        ram[15587]), .S0(n27179), .S1(n26704), .ZN(n23309) );
  MUX41 U11798 ( .I0(ram[15483]), .I1(ram[15475]), .I2(ram[15467]), .I3(
        ram[15459]), .S0(n27179), .S1(n26704), .ZN(n23304) );
  MUX41 U11799 ( .I0(ram[13819]), .I1(ram[13811]), .I2(ram[13803]), .I3(
        ram[13795]), .S0(n27175), .S1(n26700), .ZN(n23234) );
  MUX41 U11800 ( .I0(ram[13563]), .I1(ram[13555]), .I2(ram[13547]), .I3(
        ram[13539]), .S0(n27174), .S1(n26699), .ZN(n23224) );
  MUX41 U11801 ( .I0(ram[13435]), .I1(ram[13427]), .I2(ram[13419]), .I3(
        ram[13411]), .S0(n27174), .S1(n26699), .ZN(n23219) );
  MUX41 U11802 ( .I0(n22701), .I1(n22702), .I2(n22703), .I3(n22704), .S0(
        n26224), .S1(n26342), .ZN(n22700) );
  MUX41 U11803 ( .I0(ram[923]), .I1(ram[915]), .I2(ram[907]), .I3(
        ram[899]), .S0(n27144), .S1(n26669), .ZN(n22704) );
  MUX41 U11804 ( .I0(ram[955]), .I1(ram[947]), .I2(ram[939]), .I3(
        ram[931]), .S0(n27144), .S1(n26669), .ZN(n22702) );
  MUX41 U11805 ( .I0(ram[1019]), .I1(ram[1011]), .I2(ram[1003]), .I3(
        ram[995]), .S0(n27144), .S1(n26669), .ZN(n22701) );
  MUX41 U11806 ( .I0(ram[7675]), .I1(ram[7667]), .I2(ram[7659]), .I3(
        ram[7651]), .S0(n27160), .S1(n26685), .ZN(n22977) );
  MUX41 U11807 ( .I0(ram[7419]), .I1(ram[7411]), .I2(ram[7403]), .I3(
        ram[7395]), .S0(n27159), .S1(n26684), .ZN(n22967) );
  MUX41 U11808 ( .I0(ram[7291]), .I1(ram[7283]), .I2(ram[7275]), .I3(
        ram[7267]), .S0(n27159), .S1(n26684), .ZN(n22962) );
  MUX41 U11809 ( .I0(ram[5627]), .I1(ram[5619]), .I2(ram[5611]), .I3(
        ram[5603]), .S0(n27155), .S1(n26680), .ZN(n22892) );
  MUX41 U11810 ( .I0(ram[5371]), .I1(ram[5363]), .I2(ram[5355]), .I3(
        ram[5347]), .S0(n27154), .S1(n26679), .ZN(n22882) );
  MUX41 U11811 ( .I0(ram[5243]), .I1(ram[5235]), .I2(ram[5227]), .I3(
        ram[5219]), .S0(n27154), .S1(n26679), .ZN(n22877) );
  MUX41 U11812 ( .I0(ram[11771]), .I1(ram[11763]), .I2(ram[11755]), .I3(
        ram[11747]), .S0(n27170), .S1(n26695), .ZN(n23148) );
  MUX41 U11813 ( .I0(ram[11515]), .I1(ram[11507]), .I2(ram[11499]), .I3(
        ram[11491]), .S0(n27169), .S1(n26694), .ZN(n23138) );
  MUX41 U11814 ( .I0(ram[11387]), .I1(ram[11379]), .I2(ram[11371]), .I3(
        ram[11363]), .S0(n27169), .S1(n26694), .ZN(n23133) );
  MUX41 U11815 ( .I0(ram[9723]), .I1(ram[9715]), .I2(ram[9707]), .I3(
        ram[9699]), .S0(n27165), .S1(n26690), .ZN(n23063) );
  MUX41 U11816 ( .I0(ram[9467]), .I1(ram[9459]), .I2(ram[9451]), .I3(
        ram[9443]), .S0(n27164), .S1(n26689), .ZN(n23053) );
  MUX41 U11817 ( .I0(ram[9339]), .I1(ram[9331]), .I2(ram[9323]), .I3(
        ram[9315]), .S0(n27164), .S1(n26689), .ZN(n23048) );
  MUX41 U11818 ( .I0(ram[15868]), .I1(ram[15860]), .I2(ram[15852]), .I3(
        ram[15844]), .S0(n27219), .S1(n26744), .ZN(n24003) );
  MUX41 U11819 ( .I0(ram[15612]), .I1(ram[15604]), .I2(ram[15596]), .I3(
        ram[15588]), .S0(n27218), .S1(n26743), .ZN(n23993) );
  MUX41 U11820 ( .I0(ram[15484]), .I1(ram[15476]), .I2(ram[15468]), .I3(
        ram[15460]), .S0(n27218), .S1(n26743), .ZN(n23988) );
  MUX41 U11821 ( .I0(ram[13820]), .I1(ram[13812]), .I2(ram[13804]), .I3(
        ram[13796]), .S0(n27214), .S1(n26739), .ZN(n23918) );
  MUX41 U11822 ( .I0(ram[13564]), .I1(ram[13556]), .I2(ram[13548]), .I3(
        ram[13540]), .S0(n27214), .S1(n26739), .ZN(n23908) );
  MUX41 U11823 ( .I0(ram[13436]), .I1(ram[13428]), .I2(ram[13420]), .I3(
        ram[13412]), .S0(n27213), .S1(n26738), .ZN(n23903) );
  MUX41 U11824 ( .I0(n23385), .I1(n23386), .I2(n23387), .I3(n23388), .S0(
        n26234), .S1(n26352), .ZN(n23384) );
  MUX41 U11825 ( .I0(ram[924]), .I1(ram[916]), .I2(ram[908]), .I3(
        ram[900]), .S0(n27183), .S1(n26708), .ZN(n23388) );
  MUX41 U11826 ( .I0(ram[956]), .I1(ram[948]), .I2(ram[940]), .I3(
        ram[932]), .S0(n27183), .S1(n26708), .ZN(n23386) );
  MUX41 U11827 ( .I0(ram[1020]), .I1(ram[1012]), .I2(ram[1004]), .I3(
        ram[996]), .S0(n27183), .S1(n26708), .ZN(n23385) );
  MUX41 U11828 ( .I0(ram[7676]), .I1(ram[7668]), .I2(ram[7660]), .I3(
        ram[7652]), .S0(n27199), .S1(n26724), .ZN(n23661) );
  MUX41 U11829 ( .I0(ram[7420]), .I1(ram[7412]), .I2(ram[7404]), .I3(
        ram[7396]), .S0(n27199), .S1(n26724), .ZN(n23651) );
  MUX41 U11830 ( .I0(ram[7292]), .I1(ram[7284]), .I2(ram[7276]), .I3(
        ram[7268]), .S0(n27198), .S1(n26723), .ZN(n23646) );
  MUX41 U11831 ( .I0(ram[5628]), .I1(ram[5620]), .I2(ram[5612]), .I3(
        ram[5604]), .S0(n27194), .S1(n26719), .ZN(n23576) );
  MUX41 U11832 ( .I0(ram[5372]), .I1(ram[5364]), .I2(ram[5356]), .I3(
        ram[5348]), .S0(n27194), .S1(n26719), .ZN(n23566) );
  MUX41 U11833 ( .I0(ram[5244]), .I1(ram[5236]), .I2(ram[5228]), .I3(
        ram[5220]), .S0(n27194), .S1(n26719), .ZN(n23561) );
  MUX41 U11834 ( .I0(ram[11772]), .I1(ram[11764]), .I2(ram[11756]), .I3(
        ram[11748]), .S0(n27209), .S1(n26734), .ZN(n23832) );
  MUX41 U11835 ( .I0(ram[11516]), .I1(ram[11508]), .I2(ram[11500]), .I3(
        ram[11492]), .S0(n27209), .S1(n26734), .ZN(n23822) );
  MUX41 U11836 ( .I0(ram[11388]), .I1(ram[11380]), .I2(ram[11372]), .I3(
        ram[11364]), .S0(n27208), .S1(n26733), .ZN(n23817) );
  MUX41 U11837 ( .I0(ram[9724]), .I1(ram[9716]), .I2(ram[9708]), .I3(
        ram[9700]), .S0(n27204), .S1(n26729), .ZN(n23747) );
  MUX41 U11838 ( .I0(ram[9468]), .I1(ram[9460]), .I2(ram[9452]), .I3(
        ram[9444]), .S0(n27204), .S1(n26729), .ZN(n23737) );
  MUX41 U11839 ( .I0(ram[9340]), .I1(ram[9332]), .I2(ram[9324]), .I3(
        ram[9316]), .S0(n27203), .S1(n26728), .ZN(n23732) );
  MUX41 U11840 ( .I0(ram[15869]), .I1(ram[15861]), .I2(ram[15853]), .I3(
        ram[15845]), .S0(n27258), .S1(n26783), .ZN(n24687) );
  MUX41 U11841 ( .I0(ram[15613]), .I1(ram[15605]), .I2(ram[15597]), .I3(
        ram[15589]), .S0(n27258), .S1(n26783), .ZN(n24677) );
  MUX41 U11842 ( .I0(ram[15485]), .I1(ram[15477]), .I2(ram[15469]), .I3(
        ram[15461]), .S0(n27258), .S1(n26783), .ZN(n24672) );
  MUX41 U11843 ( .I0(ram[13821]), .I1(ram[13813]), .I2(ram[13805]), .I3(
        ram[13797]), .S0(n27254), .S1(n26779), .ZN(n24602) );
  MUX41 U11844 ( .I0(ram[13565]), .I1(ram[13557]), .I2(ram[13549]), .I3(
        ram[13541]), .S0(n27253), .S1(n26778), .ZN(n24592) );
  MUX41 U11845 ( .I0(ram[13437]), .I1(ram[13429]), .I2(ram[13421]), .I3(
        ram[13413]), .S0(n27253), .S1(n26778), .ZN(n24587) );
  MUX41 U11846 ( .I0(n24069), .I1(n24070), .I2(n24071), .I3(n24072), .S0(
        n26244), .S1(n26362), .ZN(n24068) );
  MUX41 U11847 ( .I0(ram[925]), .I1(ram[917]), .I2(ram[909]), .I3(
        ram[901]), .S0(n27223), .S1(n26748), .ZN(n24072) );
  MUX41 U11848 ( .I0(ram[957]), .I1(ram[949]), .I2(ram[941]), .I3(
        ram[933]), .S0(n27223), .S1(n26748), .ZN(n24070) );
  MUX41 U11849 ( .I0(ram[1021]), .I1(ram[1013]), .I2(ram[1005]), .I3(
        ram[997]), .S0(n27223), .S1(n26748), .ZN(n24069) );
  MUX41 U11850 ( .I0(ram[7677]), .I1(ram[7669]), .I2(ram[7661]), .I3(
        ram[7653]), .S0(n27239), .S1(n26764), .ZN(n24345) );
  MUX41 U11851 ( .I0(ram[7421]), .I1(ram[7413]), .I2(ram[7405]), .I3(
        ram[7397]), .S0(n27238), .S1(n26763), .ZN(n24335) );
  MUX41 U11852 ( .I0(ram[7293]), .I1(ram[7285]), .I2(ram[7277]), .I3(
        ram[7269]), .S0(n27238), .S1(n26763), .ZN(n24330) );
  MUX41 U11853 ( .I0(ram[5629]), .I1(ram[5621]), .I2(ram[5613]), .I3(
        ram[5605]), .S0(n27234), .S1(n26759), .ZN(n24260) );
  MUX41 U11854 ( .I0(ram[5373]), .I1(ram[5365]), .I2(ram[5357]), .I3(
        ram[5349]), .S0(n27233), .S1(n26758), .ZN(n24250) );
  MUX41 U11855 ( .I0(ram[5245]), .I1(ram[5237]), .I2(ram[5229]), .I3(
        ram[5221]), .S0(n27233), .S1(n26758), .ZN(n24245) );
  MUX41 U11856 ( .I0(ram[11773]), .I1(ram[11765]), .I2(ram[11757]), .I3(
        ram[11749]), .S0(n27249), .S1(n26774), .ZN(n24516) );
  MUX41 U11857 ( .I0(ram[11517]), .I1(ram[11509]), .I2(ram[11501]), .I3(
        ram[11493]), .S0(n27248), .S1(n26773), .ZN(n24506) );
  MUX41 U11858 ( .I0(ram[11389]), .I1(ram[11381]), .I2(ram[11373]), .I3(
        ram[11365]), .S0(n27248), .S1(n26773), .ZN(n24501) );
  MUX41 U11859 ( .I0(ram[9725]), .I1(ram[9717]), .I2(ram[9709]), .I3(
        ram[9701]), .S0(n27244), .S1(n26769), .ZN(n24431) );
  MUX41 U11860 ( .I0(ram[9469]), .I1(ram[9461]), .I2(ram[9453]), .I3(
        ram[9445]), .S0(n27243), .S1(n26768), .ZN(n24421) );
  MUX41 U11861 ( .I0(ram[9341]), .I1(ram[9333]), .I2(ram[9325]), .I3(
        ram[9317]), .S0(n27243), .S1(n26768), .ZN(n24416) );
  MUX41 U11862 ( .I0(ram[15870]), .I1(ram[15862]), .I2(ram[15854]), .I3(
        ram[15846]), .S0(n27298), .S1(n26823), .ZN(n25371) );
  MUX41 U11863 ( .I0(ram[15614]), .I1(ram[15606]), .I2(ram[15598]), .I3(
        ram[15590]), .S0(n27297), .S1(n26822), .ZN(n25361) );
  MUX41 U11864 ( .I0(ram[15486]), .I1(ram[15478]), .I2(ram[15470]), .I3(
        ram[15462]), .S0(n27297), .S1(n26822), .ZN(n25356) );
  MUX41 U11865 ( .I0(ram[13822]), .I1(ram[13814]), .I2(ram[13806]), .I3(
        ram[13798]), .S0(n27293), .S1(n26818), .ZN(n25286) );
  MUX41 U11866 ( .I0(ram[13566]), .I1(ram[13558]), .I2(ram[13550]), .I3(
        ram[13542]), .S0(n27292), .S1(n26817), .ZN(n25276) );
  MUX41 U11867 ( .I0(ram[13438]), .I1(ram[13430]), .I2(ram[13422]), .I3(
        ram[13414]), .S0(n27292), .S1(n26817), .ZN(n25271) );
  MUX41 U11868 ( .I0(n24753), .I1(n24754), .I2(n24755), .I3(n24756), .S0(
        n26253), .S1(n26371), .ZN(n24752) );
  MUX41 U11869 ( .I0(ram[926]), .I1(ram[918]), .I2(ram[910]), .I3(
        ram[902]), .S0(n27262), .S1(n26787), .ZN(n24756) );
  MUX41 U11870 ( .I0(ram[958]), .I1(ram[950]), .I2(ram[942]), .I3(
        ram[934]), .S0(n27262), .S1(n26787), .ZN(n24754) );
  MUX41 U11871 ( .I0(ram[1022]), .I1(ram[1014]), .I2(ram[1006]), .I3(
        ram[998]), .S0(n27262), .S1(n26787), .ZN(n24753) );
  MUX41 U11872 ( .I0(ram[7678]), .I1(ram[7670]), .I2(ram[7662]), .I3(
        ram[7654]), .S0(n27278), .S1(n26803), .ZN(n25029) );
  MUX41 U11873 ( .I0(ram[7422]), .I1(ram[7414]), .I2(ram[7406]), .I3(
        ram[7398]), .S0(n27278), .S1(n26803), .ZN(n25019) );
  MUX41 U11874 ( .I0(ram[7294]), .I1(ram[7286]), .I2(ram[7278]), .I3(
        ram[7270]), .S0(n27277), .S1(n26802), .ZN(n25014) );
  MUX41 U11875 ( .I0(ram[5630]), .I1(ram[5622]), .I2(ram[5614]), .I3(
        ram[5606]), .S0(n27273), .S1(n26798), .ZN(n24944) );
  MUX41 U11876 ( .I0(ram[5374]), .I1(ram[5366]), .I2(ram[5358]), .I3(
        ram[5350]), .S0(n27273), .S1(n26798), .ZN(n24934) );
  MUX41 U11877 ( .I0(ram[5246]), .I1(ram[5238]), .I2(ram[5230]), .I3(
        ram[5222]), .S0(n27272), .S1(n26797), .ZN(n24929) );
  MUX41 U11878 ( .I0(ram[11774]), .I1(ram[11766]), .I2(ram[11758]), .I3(
        ram[11750]), .S0(n27288), .S1(n26813), .ZN(n25200) );
  MUX41 U11879 ( .I0(ram[11518]), .I1(ram[11510]), .I2(ram[11502]), .I3(
        ram[11494]), .S0(n27287), .S1(n26812), .ZN(n25190) );
  MUX41 U11880 ( .I0(ram[11390]), .I1(ram[11382]), .I2(ram[11374]), .I3(
        ram[11366]), .S0(n27287), .S1(n26812), .ZN(n25185) );
  MUX41 U11881 ( .I0(ram[9726]), .I1(ram[9718]), .I2(ram[9710]), .I3(
        ram[9702]), .S0(n27283), .S1(n26808), .ZN(n25115) );
  MUX41 U11882 ( .I0(ram[9470]), .I1(ram[9462]), .I2(ram[9454]), .I3(
        ram[9446]), .S0(n27282), .S1(n26807), .ZN(n25105) );
  MUX41 U11883 ( .I0(ram[9342]), .I1(ram[9334]), .I2(ram[9326]), .I3(
        ram[9318]), .S0(n27282), .S1(n26807), .ZN(n25100) );
  MUX41 U11884 ( .I0(ram[15871]), .I1(ram[15863]), .I2(ram[15855]), .I3(
        ram[15847]), .S0(n27337), .S1(n26862), .ZN(n26055) );
  MUX41 U11885 ( .I0(ram[15615]), .I1(ram[15607]), .I2(ram[15599]), .I3(
        ram[15591]), .S0(n27337), .S1(n26862), .ZN(n26045) );
  MUX41 U11886 ( .I0(ram[15487]), .I1(ram[15479]), .I2(ram[15471]), .I3(
        ram[15463]), .S0(n27336), .S1(n26861), .ZN(n26040) );
  MUX41 U11887 ( .I0(ram[13823]), .I1(ram[13815]), .I2(ram[13807]), .I3(
        ram[13799]), .S0(n27332), .S1(n26857), .ZN(n25970) );
  MUX41 U11888 ( .I0(ram[13567]), .I1(ram[13559]), .I2(ram[13551]), .I3(
        ram[13543]), .S0(n27332), .S1(n26857), .ZN(n25960) );
  MUX41 U11889 ( .I0(ram[13439]), .I1(ram[13431]), .I2(ram[13423]), .I3(
        ram[13415]), .S0(n27331), .S1(n26856), .ZN(n25955) );
  MUX41 U11890 ( .I0(n25437), .I1(n25438), .I2(n25439), .I3(n25440), .S0(
        n26263), .S1(n26381), .ZN(n25436) );
  MUX41 U11891 ( .I0(ram[927]), .I1(ram[919]), .I2(ram[911]), .I3(
        ram[903]), .S0(n27301), .S1(n26826), .ZN(n25440) );
  MUX41 U11892 ( .I0(ram[959]), .I1(ram[951]), .I2(ram[943]), .I3(
        ram[935]), .S0(n27301), .S1(n26826), .ZN(n25438) );
  MUX41 U11893 ( .I0(ram[1023]), .I1(ram[1015]), .I2(ram[1007]), .I3(
        ram[999]), .S0(n27302), .S1(n26827), .ZN(n25437) );
  MUX41 U11894 ( .I0(ram[7679]), .I1(ram[7671]), .I2(ram[7663]), .I3(
        ram[7655]), .S0(n27318), .S1(n26843), .ZN(n25713) );
  MUX41 U11895 ( .I0(ram[7423]), .I1(ram[7415]), .I2(ram[7407]), .I3(
        ram[7399]), .S0(n27317), .S1(n26842), .ZN(n25703) );
  MUX41 U11896 ( .I0(ram[7295]), .I1(ram[7287]), .I2(ram[7279]), .I3(
        ram[7271]), .S0(n27317), .S1(n26842), .ZN(n25698) );
  MUX41 U11897 ( .I0(ram[5631]), .I1(ram[5623]), .I2(ram[5615]), .I3(
        ram[5607]), .S0(n27313), .S1(n26838), .ZN(n25628) );
  MUX41 U11898 ( .I0(ram[5375]), .I1(ram[5367]), .I2(ram[5359]), .I3(
        ram[5351]), .S0(n27312), .S1(n26837), .ZN(n25618) );
  MUX41 U11899 ( .I0(ram[5247]), .I1(ram[5239]), .I2(ram[5231]), .I3(
        ram[5223]), .S0(n27312), .S1(n26837), .ZN(n25613) );
  MUX41 U11900 ( .I0(ram[11775]), .I1(ram[11767]), .I2(ram[11759]), .I3(
        ram[11751]), .S0(n27327), .S1(n26852), .ZN(n25884) );
  MUX41 U11901 ( .I0(ram[11519]), .I1(ram[11511]), .I2(ram[11503]), .I3(
        ram[11495]), .S0(n27327), .S1(n26852), .ZN(n25874) );
  MUX41 U11902 ( .I0(ram[11391]), .I1(ram[11383]), .I2(ram[11375]), .I3(
        ram[11367]), .S0(n27326), .S1(n26851), .ZN(n25869) );
  MUX41 U11903 ( .I0(ram[9727]), .I1(ram[9719]), .I2(ram[9711]), .I3(
        ram[9703]), .S0(n27322), .S1(n26847), .ZN(n25799) );
  MUX41 U11904 ( .I0(ram[9471]), .I1(ram[9463]), .I2(ram[9455]), .I3(
        ram[9447]), .S0(n27322), .S1(n26847), .ZN(n25789) );
  MUX41 U11905 ( .I0(ram[9343]), .I1(ram[9335]), .I2(ram[9327]), .I3(
        ram[9319]), .S0(n27322), .S1(n26847), .ZN(n25784) );
  MUX41 U11906 ( .I0(n21287), .I1(n21288), .I2(n21289), .I3(n21290), .S0(
        n26204), .S1(n26322), .ZN(n21286) );
  MUX41 U11907 ( .I0(ram[16280]), .I1(ram[16272]), .I2(ram[16264]), .I3(
        ram[16256]), .S0(n27063), .S1(n26588), .ZN(n21290) );
  MUX41 U11908 ( .I0(ram[16312]), .I1(ram[16304]), .I2(ram[16296]), .I3(
        ram[16288]), .S0(n27063), .S1(n26588), .ZN(n21288) );
  MUX41 U11909 ( .I0(ram[16376]), .I1(ram[16368]), .I2(ram[16360]), .I3(
        ram[16352]), .S0(n27063), .S1(n26588), .ZN(n21287) );
  MUX41 U11910 ( .I0(n21247), .I1(n21248), .I2(n21249), .I3(n21250), .S0(
        n26203), .S1(n26321), .ZN(n21246) );
  MUX41 U11911 ( .I0(ram[15256]), .I1(ram[15248]), .I2(ram[15240]), .I3(
        ram[15232]), .S0(n27060), .S1(n26585), .ZN(n21250) );
  MUX41 U11912 ( .I0(ram[15288]), .I1(ram[15280]), .I2(ram[15272]), .I3(
        ram[15264]), .S0(n27060), .S1(n26585), .ZN(n21248) );
  MUX41 U11913 ( .I0(ram[15352]), .I1(ram[15344]), .I2(ram[15336]), .I3(
        ram[15328]), .S0(n27060), .S1(n26585), .ZN(n21247) );
  MUX41 U11914 ( .I0(n21227), .I1(n21228), .I2(n21229), .I3(n21230), .S0(
        n26203), .S1(n26321), .ZN(n21226) );
  MUX41 U11915 ( .I0(ram[14744]), .I1(ram[14736]), .I2(ram[14728]), .I3(
        ram[14720]), .S0(n27059), .S1(n26584), .ZN(n21230) );
  MUX41 U11916 ( .I0(ram[14776]), .I1(ram[14768]), .I2(ram[14760]), .I3(
        ram[14752]), .S0(n27059), .S1(n26584), .ZN(n21228) );
  MUX41 U11917 ( .I0(ram[14840]), .I1(ram[14832]), .I2(ram[14824]), .I3(
        ram[14816]), .S0(n27059), .S1(n26584), .ZN(n21227) );
  MUX41 U11918 ( .I0(n21202), .I1(n21203), .I2(n21204), .I3(n21205), .S0(
        n26202), .S1(n26320), .ZN(n21201) );
  MUX41 U11919 ( .I0(ram[14232]), .I1(ram[14224]), .I2(ram[14216]), .I3(
        ram[14208]), .S0(n27058), .S1(n26583), .ZN(n21205) );
  MUX41 U11920 ( .I0(ram[14264]), .I1(ram[14256]), .I2(ram[14248]), .I3(
        ram[14240]), .S0(n27058), .S1(n26583), .ZN(n21203) );
  MUX41 U11921 ( .I0(ram[14328]), .I1(ram[14320]), .I2(ram[14312]), .I3(
        ram[14304]), .S0(n27058), .S1(n26583), .ZN(n21202) );
  MUX41 U11922 ( .I0(n21162), .I1(n21163), .I2(n21164), .I3(n21165), .S0(
        n26202), .S1(n26320), .ZN(n21161) );
  MUX41 U11923 ( .I0(ram[13208]), .I1(ram[13200]), .I2(ram[13192]), .I3(
        ram[13184]), .S0(n27055), .S1(n26580), .ZN(n21165) );
  MUX41 U11924 ( .I0(ram[13240]), .I1(ram[13232]), .I2(ram[13224]), .I3(
        ram[13216]), .S0(n27055), .S1(n26580), .ZN(n21163) );
  MUX41 U11925 ( .I0(ram[13304]), .I1(ram[13296]), .I2(ram[13288]), .I3(
        ram[13280]), .S0(n27055), .S1(n26580), .ZN(n21162) );
  MUX41 U11926 ( .I0(n21142), .I1(n21143), .I2(n21144), .I3(n21145), .S0(
        n26201), .S1(n26319), .ZN(n21141) );
  MUX41 U11927 ( .I0(ram[12696]), .I1(ram[12688]), .I2(ram[12680]), .I3(
        ram[12672]), .S0(n27054), .S1(n26579), .ZN(n21145) );
  MUX41 U11928 ( .I0(ram[12728]), .I1(ram[12720]), .I2(ram[12712]), .I3(
        ram[12704]), .S0(n27054), .S1(n26579), .ZN(n21143) );
  MUX41 U11929 ( .I0(ram[12792]), .I1(ram[12784]), .I2(ram[12776]), .I3(
        ram[12768]), .S0(n27054), .S1(n26579), .ZN(n21142) );
  MUX41 U11930 ( .I0(n20945), .I1(n20946), .I2(n20947), .I3(n20948), .S0(
        n26199), .S1(n26317), .ZN(n20944) );
  MUX41 U11931 ( .I0(ram[8120]), .I1(ram[8112]), .I2(ram[8104]), .I3(
        ram[8096]), .S0(n27043), .S1(n26568), .ZN(n20946) );
  MUX41 U11932 ( .I0(ram[8088]), .I1(ram[8080]), .I2(ram[8072]), .I3(
        ram[8064]), .S0(n27043), .S1(n26568), .ZN(n20948) );
  MUX41 U11933 ( .I0(ram[8184]), .I1(ram[8176]), .I2(ram[8168]), .I3(
        ram[8160]), .S0(n27043), .S1(n26568), .ZN(n20945) );
  MUX41 U11934 ( .I0(n20885), .I1(n20886), .I2(n20887), .I3(n20888), .S0(
        n26198), .S1(n26316), .ZN(n20884) );
  MUX41 U11935 ( .I0(ram[6552]), .I1(ram[6544]), .I2(ram[6536]), .I3(
        ram[6528]), .S0(n27039), .S1(n26564), .ZN(n20888) );
  MUX41 U11936 ( .I0(ram[6584]), .I1(ram[6576]), .I2(ram[6568]), .I3(
        ram[6560]), .S0(n27039), .S1(n26564), .ZN(n20886) );
  MUX41 U11937 ( .I0(ram[6648]), .I1(ram[6640]), .I2(ram[6632]), .I3(
        ram[6624]), .S0(n27039), .S1(n26564), .ZN(n20885) );
  MUX41 U11938 ( .I0(n20905), .I1(n20906), .I2(n20907), .I3(n20908), .S0(
        n26198), .S1(n26316), .ZN(n20904) );
  MUX41 U11939 ( .I0(ram[7064]), .I1(ram[7056]), .I2(ram[7048]), .I3(
        ram[7040]), .S0(n27040), .S1(n26565), .ZN(n20908) );
  MUX41 U11940 ( .I0(ram[7096]), .I1(ram[7088]), .I2(ram[7080]), .I3(
        ram[7072]), .S0(n27040), .S1(n26565), .ZN(n20906) );
  MUX41 U11941 ( .I0(ram[7160]), .I1(ram[7152]), .I2(ram[7144]), .I3(
        ram[7136]), .S0(n27041), .S1(n26566), .ZN(n20905) );
  MUX41 U11942 ( .I0(n20860), .I1(n20861), .I2(n20862), .I3(n20863), .S0(
        n26197), .S1(n26315), .ZN(n20859) );
  MUX41 U11943 ( .I0(ram[6072]), .I1(ram[6064]), .I2(ram[6056]), .I3(
        ram[6048]), .S0(n27038), .S1(n26563), .ZN(n20861) );
  MUX41 U11944 ( .I0(ram[6040]), .I1(ram[6032]), .I2(ram[6024]), .I3(
        ram[6016]), .S0(n27038), .S1(n26563), .ZN(n20863) );
  MUX41 U11945 ( .I0(ram[6136]), .I1(ram[6128]), .I2(ram[6120]), .I3(
        ram[6112]), .S0(n27038), .S1(n26563), .ZN(n20860) );
  MUX41 U11946 ( .I0(n20800), .I1(n20801), .I2(n20802), .I3(n20803), .S0(
        n26196), .S1(n26314), .ZN(n20799) );
  MUX41 U11947 ( .I0(ram[4536]), .I1(ram[4528]), .I2(ram[4520]), .I3(
        ram[4512]), .S0(n27034), .S1(n26559), .ZN(n20801) );
  MUX41 U11948 ( .I0(ram[4504]), .I1(ram[4496]), .I2(ram[4488]), .I3(
        ram[4480]), .S0(n27034), .S1(n26559), .ZN(n20803) );
  MUX41 U11949 ( .I0(ram[4600]), .I1(ram[4592]), .I2(ram[4584]), .I3(
        ram[4576]), .S0(n27034), .S1(n26559), .ZN(n20800) );
  MUX41 U11950 ( .I0(n21116), .I1(n21117), .I2(n21118), .I3(n21119), .S0(
        n26201), .S1(n26319), .ZN(n21115) );
  MUX41 U11951 ( .I0(ram[12216]), .I1(ram[12208]), .I2(ram[12200]), .I3(
        ram[12192]), .S0(n27053), .S1(n26578), .ZN(n21117) );
  MUX41 U11952 ( .I0(ram[12184]), .I1(ram[12176]), .I2(ram[12168]), .I3(
        ram[12160]), .S0(n27053), .S1(n26578), .ZN(n21119) );
  MUX41 U11953 ( .I0(ram[12280]), .I1(ram[12272]), .I2(ram[12264]), .I3(
        ram[12256]), .S0(n27053), .S1(n26578), .ZN(n21116) );
  MUX41 U11954 ( .I0(n21056), .I1(n21057), .I2(n21058), .I3(n21059), .S0(
        n26200), .S1(n26318), .ZN(n21055) );
  MUX41 U11955 ( .I0(ram[10680]), .I1(ram[10672]), .I2(ram[10664]), .I3(
        ram[10656]), .S0(n27049), .S1(n26574), .ZN(n21057) );
  MUX41 U11956 ( .I0(ram[10648]), .I1(ram[10640]), .I2(ram[10632]), .I3(
        ram[10624]), .S0(n27049), .S1(n26574), .ZN(n21059) );
  MUX41 U11957 ( .I0(ram[10744]), .I1(ram[10736]), .I2(ram[10728]), .I3(
        ram[10720]), .S0(n27049), .S1(n26574), .ZN(n21056) );
  MUX41 U11958 ( .I0(n21076), .I1(n21077), .I2(n21078), .I3(n21079), .S0(
        n26200), .S1(n26318), .ZN(n21075) );
  MUX41 U11959 ( .I0(ram[11192]), .I1(ram[11184]), .I2(ram[11176]), .I3(
        ram[11168]), .S0(n27050), .S1(n26575), .ZN(n21077) );
  MUX41 U11960 ( .I0(ram[11160]), .I1(ram[11152]), .I2(ram[11144]), .I3(
        ram[11136]), .S0(n27050), .S1(n26575), .ZN(n21079) );
  MUX41 U11961 ( .I0(ram[11256]), .I1(ram[11248]), .I2(ram[11240]), .I3(
        ram[11232]), .S0(n27050), .S1(n26575), .ZN(n21076) );
  MUX41 U11962 ( .I0(n21031), .I1(n21032), .I2(n21033), .I3(n21034), .S0(
        n26200), .S1(n26318), .ZN(n21030) );
  MUX41 U11963 ( .I0(ram[10168]), .I1(ram[10160]), .I2(ram[10152]), .I3(
        ram[10144]), .S0(n27048), .S1(n26573), .ZN(n21032) );
  MUX41 U11964 ( .I0(ram[10136]), .I1(ram[10128]), .I2(ram[10120]), .I3(
        ram[10112]), .S0(n27048), .S1(n26573), .ZN(n21034) );
  MUX41 U11965 ( .I0(ram[10232]), .I1(ram[10224]), .I2(ram[10216]), .I3(
        ram[10208]), .S0(n27048), .S1(n26573), .ZN(n21031) );
  MUX41 U11966 ( .I0(n20971), .I1(n20972), .I2(n20973), .I3(n20974), .S0(
        n26199), .S1(n26317), .ZN(n20970) );
  MUX41 U11967 ( .I0(ram[8632]), .I1(ram[8624]), .I2(ram[8616]), .I3(
        ram[8608]), .S0(n27044), .S1(n26569), .ZN(n20972) );
  MUX41 U11968 ( .I0(ram[8600]), .I1(ram[8592]), .I2(ram[8584]), .I3(
        ram[8576]), .S0(n27044), .S1(n26569), .ZN(n20974) );
  MUX41 U11969 ( .I0(ram[8696]), .I1(ram[8688]), .I2(ram[8680]), .I3(
        ram[8672]), .S0(n27044), .S1(n26569), .ZN(n20971) );
  MUX41 U11970 ( .I0(n20991), .I1(n20992), .I2(n20993), .I3(n20994), .S0(
        n26199), .S1(n26317), .ZN(n20990) );
  MUX41 U11971 ( .I0(ram[9112]), .I1(ram[9104]), .I2(ram[9096]), .I3(
        ram[9088]), .S0(n27045), .S1(n26570), .ZN(n20994) );
  MUX41 U11972 ( .I0(ram[9144]), .I1(ram[9136]), .I2(ram[9128]), .I3(
        ram[9120]), .S0(n27045), .S1(n26570), .ZN(n20992) );
  MUX41 U11973 ( .I0(ram[9208]), .I1(ram[9200]), .I2(ram[9192]), .I3(
        ram[9184]), .S0(n27046), .S1(n26571), .ZN(n20991) );
  MUX41 U11974 ( .I0(n21971), .I1(n21972), .I2(n21973), .I3(n21974), .S0(
        n26213), .S1(n26331), .ZN(n21970) );
  MUX41 U11975 ( .I0(ram[16281]), .I1(ram[16273]), .I2(ram[16265]), .I3(
        ram[16257]), .S0(n27102), .S1(n26627), .ZN(n21974) );
  MUX41 U11976 ( .I0(ram[16313]), .I1(ram[16305]), .I2(ram[16297]), .I3(
        ram[16289]), .S0(n27102), .S1(n26627), .ZN(n21972) );
  MUX41 U11977 ( .I0(ram[16377]), .I1(ram[16369]), .I2(ram[16361]), .I3(
        ram[16353]), .S0(n27102), .S1(n26627), .ZN(n21971) );
  MUX41 U11978 ( .I0(n21931), .I1(n21932), .I2(n21933), .I3(n21934), .S0(
        n26213), .S1(n26331), .ZN(n21930) );
  MUX41 U11979 ( .I0(ram[15257]), .I1(ram[15249]), .I2(ram[15241]), .I3(
        ram[15233]), .S0(n27099), .S1(n26624), .ZN(n21934) );
  MUX41 U11980 ( .I0(ram[15289]), .I1(ram[15281]), .I2(ram[15273]), .I3(
        ram[15265]), .S0(n27100), .S1(n26625), .ZN(n21932) );
  MUX41 U11981 ( .I0(ram[15353]), .I1(ram[15345]), .I2(ram[15337]), .I3(
        ram[15329]), .S0(n27100), .S1(n26625), .ZN(n21931) );
  MUX41 U11982 ( .I0(n21911), .I1(n21912), .I2(n21913), .I3(n21914), .S0(
        n26212), .S1(n26330), .ZN(n21910) );
  MUX41 U11983 ( .I0(ram[14745]), .I1(ram[14737]), .I2(ram[14729]), .I3(
        ram[14721]), .S0(n27098), .S1(n26623), .ZN(n21914) );
  MUX41 U11984 ( .I0(ram[14777]), .I1(ram[14769]), .I2(ram[14761]), .I3(
        ram[14753]), .S0(n27098), .S1(n26623), .ZN(n21912) );
  MUX41 U11985 ( .I0(ram[14841]), .I1(ram[14833]), .I2(ram[14825]), .I3(
        ram[14817]), .S0(n27098), .S1(n26623), .ZN(n21911) );
  MUX41 U11986 ( .I0(n21886), .I1(n21887), .I2(n21888), .I3(n21889), .S0(
        n26212), .S1(n26330), .ZN(n21885) );
  MUX41 U11987 ( .I0(ram[14233]), .I1(ram[14225]), .I2(ram[14217]), .I3(
        ram[14209]), .S0(n27097), .S1(n26622), .ZN(n21889) );
  MUX41 U11988 ( .I0(ram[14265]), .I1(ram[14257]), .I2(ram[14249]), .I3(
        ram[14241]), .S0(n27097), .S1(n26622), .ZN(n21887) );
  MUX41 U11989 ( .I0(ram[14329]), .I1(ram[14321]), .I2(ram[14313]), .I3(
        ram[14305]), .S0(n27097), .S1(n26622), .ZN(n21886) );
  MUX41 U11990 ( .I0(n21846), .I1(n21847), .I2(n21848), .I3(n21849), .S0(
        n26212), .S1(n26330), .ZN(n21845) );
  MUX41 U11991 ( .I0(ram[13209]), .I1(ram[13201]), .I2(ram[13193]), .I3(
        ram[13185]), .S0(n27095), .S1(n26620), .ZN(n21849) );
  MUX41 U11992 ( .I0(ram[13241]), .I1(ram[13233]), .I2(ram[13225]), .I3(
        ram[13217]), .S0(n27095), .S1(n26620), .ZN(n21847) );
  MUX41 U11993 ( .I0(ram[13305]), .I1(ram[13297]), .I2(ram[13289]), .I3(
        ram[13281]), .S0(n27095), .S1(n26620), .ZN(n21846) );
  MUX41 U11994 ( .I0(n21826), .I1(n21827), .I2(n21828), .I3(n21829), .S0(
        n26211), .S1(n26329), .ZN(n21825) );
  MUX41 U11995 ( .I0(ram[12697]), .I1(ram[12689]), .I2(ram[12681]), .I3(
        ram[12673]), .S0(n27093), .S1(n26618), .ZN(n21829) );
  MUX41 U11996 ( .I0(ram[12729]), .I1(ram[12721]), .I2(ram[12713]), .I3(
        ram[12705]), .S0(n27093), .S1(n26618), .ZN(n21827) );
  MUX41 U11997 ( .I0(ram[12793]), .I1(ram[12785]), .I2(ram[12777]), .I3(
        ram[12769]), .S0(n27094), .S1(n26619), .ZN(n21826) );
  MUX41 U11998 ( .I0(n21629), .I1(n21630), .I2(n21631), .I3(n21632), .S0(
        n26208), .S1(n26326), .ZN(n21628) );
  MUX41 U11999 ( .I0(ram[8121]), .I1(ram[8113]), .I2(ram[8105]), .I3(
        ram[8097]), .S0(n27082), .S1(n26607), .ZN(n21630) );
  MUX41 U12000 ( .I0(ram[8089]), .I1(ram[8081]), .I2(ram[8073]), .I3(
        ram[8065]), .S0(n27082), .S1(n26607), .ZN(n21632) );
  MUX41 U12001 ( .I0(ram[8185]), .I1(ram[8177]), .I2(ram[8169]), .I3(
        ram[8161]), .S0(n27082), .S1(n26607), .ZN(n21629) );
  MUX41 U12002 ( .I0(n21569), .I1(n21570), .I2(n21571), .I3(n21572), .S0(
        n26208), .S1(n26326), .ZN(n21568) );
  MUX41 U12003 ( .I0(ram[6553]), .I1(ram[6545]), .I2(ram[6537]), .I3(
        ram[6529]), .S0(n27079), .S1(n26604), .ZN(n21572) );
  MUX41 U12004 ( .I0(ram[6585]), .I1(ram[6577]), .I2(ram[6569]), .I3(
        ram[6561]), .S0(n27079), .S1(n26604), .ZN(n21570) );
  MUX41 U12005 ( .I0(ram[6649]), .I1(ram[6641]), .I2(ram[6633]), .I3(
        ram[6625]), .S0(n27079), .S1(n26604), .ZN(n21569) );
  MUX41 U12006 ( .I0(n21589), .I1(n21590), .I2(n21591), .I3(n21592), .S0(
        n26208), .S1(n26326), .ZN(n21588) );
  MUX41 U12007 ( .I0(ram[7065]), .I1(ram[7057]), .I2(ram[7049]), .I3(
        ram[7041]), .S0(n27080), .S1(n26605), .ZN(n21592) );
  MUX41 U12008 ( .I0(ram[7097]), .I1(ram[7089]), .I2(ram[7081]), .I3(
        ram[7073]), .S0(n27080), .S1(n26605), .ZN(n21590) );
  MUX41 U12009 ( .I0(ram[7161]), .I1(ram[7153]), .I2(ram[7145]), .I3(
        ram[7137]), .S0(n27080), .S1(n26605), .ZN(n21589) );
  MUX41 U12010 ( .I0(n21544), .I1(n21545), .I2(n21546), .I3(n21547), .S0(
        n26207), .S1(n26325), .ZN(n21543) );
  MUX41 U12011 ( .I0(ram[6073]), .I1(ram[6065]), .I2(ram[6057]), .I3(
        ram[6049]), .S0(n27077), .S1(n26602), .ZN(n21545) );
  MUX41 U12012 ( .I0(ram[6041]), .I1(ram[6033]), .I2(ram[6025]), .I3(
        ram[6017]), .S0(n27077), .S1(n26602), .ZN(n21547) );
  MUX41 U12013 ( .I0(ram[6137]), .I1(ram[6129]), .I2(ram[6121]), .I3(
        ram[6113]), .S0(n27078), .S1(n26603), .ZN(n21544) );
  MUX41 U12014 ( .I0(n21484), .I1(n21485), .I2(n21486), .I3(n21487), .S0(
        n26206), .S1(n26324), .ZN(n21483) );
  MUX41 U12015 ( .I0(ram[4537]), .I1(ram[4529]), .I2(ram[4521]), .I3(
        ram[4513]), .S0(n27074), .S1(n26599), .ZN(n21485) );
  MUX41 U12016 ( .I0(ram[4505]), .I1(ram[4497]), .I2(ram[4489]), .I3(
        ram[4481]), .S0(n27074), .S1(n26599), .ZN(n21487) );
  MUX41 U12017 ( .I0(ram[4601]), .I1(ram[4593]), .I2(ram[4585]), .I3(
        ram[4577]), .S0(n27074), .S1(n26599), .ZN(n21484) );
  MUX41 U12018 ( .I0(n21800), .I1(n21801), .I2(n21802), .I3(n21803), .S0(
        n26211), .S1(n26329), .ZN(n21799) );
  MUX41 U12019 ( .I0(ram[12217]), .I1(ram[12209]), .I2(ram[12201]), .I3(
        ram[12193]), .S0(n27092), .S1(n26617), .ZN(n21801) );
  MUX41 U12020 ( .I0(ram[12185]), .I1(ram[12177]), .I2(ram[12169]), .I3(
        ram[12161]), .S0(n27092), .S1(n26617), .ZN(n21803) );
  MUX41 U12021 ( .I0(ram[12281]), .I1(ram[12273]), .I2(ram[12265]), .I3(
        ram[12257]), .S0(n27092), .S1(n26617), .ZN(n21800) );
  MUX41 U12022 ( .I0(n21740), .I1(n21741), .I2(n21742), .I3(n21743), .S0(
        n26210), .S1(n26328), .ZN(n21739) );
  MUX41 U12023 ( .I0(ram[10681]), .I1(ram[10673]), .I2(ram[10665]), .I3(
        ram[10657]), .S0(n27088), .S1(n26613), .ZN(n21741) );
  MUX41 U12024 ( .I0(ram[10649]), .I1(ram[10641]), .I2(ram[10633]), .I3(
        ram[10625]), .S0(n27088), .S1(n26613), .ZN(n21743) );
  MUX41 U12025 ( .I0(ram[10745]), .I1(ram[10737]), .I2(ram[10729]), .I3(
        ram[10721]), .S0(n27089), .S1(n26614), .ZN(n21740) );
  MUX41 U12026 ( .I0(n21760), .I1(n21761), .I2(n21762), .I3(n21763), .S0(
        n26210), .S1(n26328), .ZN(n21759) );
  MUX41 U12027 ( .I0(ram[11193]), .I1(ram[11185]), .I2(ram[11177]), .I3(
        ram[11169]), .S0(n27090), .S1(n26615), .ZN(n21761) );
  MUX41 U12028 ( .I0(ram[11161]), .I1(ram[11153]), .I2(ram[11145]), .I3(
        ram[11137]), .S0(n27090), .S1(n26615), .ZN(n21763) );
  MUX41 U12029 ( .I0(ram[11257]), .I1(ram[11249]), .I2(ram[11241]), .I3(
        ram[11233]), .S0(n27090), .S1(n26615), .ZN(n21760) );
  MUX41 U12030 ( .I0(n21715), .I1(n21716), .I2(n21717), .I3(n21718), .S0(
        n26210), .S1(n26328), .ZN(n21714) );
  MUX41 U12031 ( .I0(ram[10169]), .I1(ram[10161]), .I2(ram[10153]), .I3(
        ram[10145]), .S0(n27087), .S1(n26612), .ZN(n21716) );
  MUX41 U12032 ( .I0(ram[10137]), .I1(ram[10129]), .I2(ram[10121]), .I3(
        ram[10113]), .S0(n27087), .S1(n26612), .ZN(n21718) );
  MUX41 U12033 ( .I0(ram[10233]), .I1(ram[10225]), .I2(ram[10217]), .I3(
        ram[10209]), .S0(n27087), .S1(n26612), .ZN(n21715) );
  MUX41 U12034 ( .I0(n21655), .I1(n21656), .I2(n21657), .I3(n21658), .S0(
        n26209), .S1(n26327), .ZN(n21654) );
  MUX41 U12035 ( .I0(ram[8633]), .I1(ram[8625]), .I2(ram[8617]), .I3(
        ram[8609]), .S0(n27084), .S1(n26609), .ZN(n21656) );
  MUX41 U12036 ( .I0(ram[8601]), .I1(ram[8593]), .I2(ram[8585]), .I3(
        ram[8577]), .S0(n27083), .S1(n26608), .ZN(n21658) );
  MUX41 U12037 ( .I0(ram[8697]), .I1(ram[8689]), .I2(ram[8681]), .I3(
        ram[8673]), .S0(n27084), .S1(n26609), .ZN(n21655) );
  MUX41 U12038 ( .I0(n21675), .I1(n21676), .I2(n21677), .I3(n21678), .S0(
        n26209), .S1(n26327), .ZN(n21674) );
  MUX41 U12039 ( .I0(ram[9113]), .I1(ram[9105]), .I2(ram[9097]), .I3(
        ram[9089]), .S0(n27085), .S1(n26610), .ZN(n21678) );
  MUX41 U12040 ( .I0(ram[9145]), .I1(ram[9137]), .I2(ram[9129]), .I3(
        ram[9121]), .S0(n27085), .S1(n26610), .ZN(n21676) );
  MUX41 U12041 ( .I0(ram[9209]), .I1(ram[9201]), .I2(ram[9193]), .I3(
        ram[9185]), .S0(n27085), .S1(n26610), .ZN(n21675) );
  MUX41 U12042 ( .I0(n22655), .I1(n22656), .I2(n22657), .I3(n22658), .S0(
        n26223), .S1(n26341), .ZN(n22654) );
  MUX41 U12043 ( .I0(ram[16282]), .I1(ram[16274]), .I2(ram[16266]), .I3(
        ram[16258]), .S0(n27141), .S1(n26666), .ZN(n22658) );
  MUX41 U12044 ( .I0(ram[16314]), .I1(ram[16306]), .I2(ram[16298]), .I3(
        ram[16290]), .S0(n27141), .S1(n26666), .ZN(n22656) );
  MUX41 U12045 ( .I0(ram[16378]), .I1(ram[16370]), .I2(ram[16362]), .I3(
        ram[16354]), .S0(n27142), .S1(n26667), .ZN(n22655) );
  MUX41 U12046 ( .I0(n22615), .I1(n22616), .I2(n22617), .I3(n22618), .S0(
        n26223), .S1(n26341), .ZN(n22614) );
  MUX41 U12047 ( .I0(ram[15258]), .I1(ram[15250]), .I2(ram[15242]), .I3(
        ram[15234]), .S0(n27139), .S1(n26664), .ZN(n22618) );
  MUX41 U12048 ( .I0(ram[15290]), .I1(ram[15282]), .I2(ram[15274]), .I3(
        ram[15266]), .S0(n27139), .S1(n26664), .ZN(n22616) );
  MUX41 U12049 ( .I0(ram[15354]), .I1(ram[15346]), .I2(ram[15338]), .I3(
        ram[15330]), .S0(n27139), .S1(n26664), .ZN(n22615) );
  MUX41 U12050 ( .I0(n22595), .I1(n22596), .I2(n22597), .I3(n22598), .S0(
        n26222), .S1(n26340), .ZN(n22594) );
  MUX41 U12051 ( .I0(ram[14746]), .I1(ram[14738]), .I2(ram[14730]), .I3(
        ram[14722]), .S0(n27138), .S1(n26663), .ZN(n22598) );
  MUX41 U12052 ( .I0(ram[14778]), .I1(ram[14770]), .I2(ram[14762]), .I3(
        ram[14754]), .S0(n27138), .S1(n26663), .ZN(n22596) );
  MUX41 U12053 ( .I0(ram[14842]), .I1(ram[14834]), .I2(ram[14826]), .I3(
        ram[14818]), .S0(n27138), .S1(n26663), .ZN(n22595) );
  MUX41 U12054 ( .I0(n22570), .I1(n22571), .I2(n22572), .I3(n22573), .S0(
        n26222), .S1(n26340), .ZN(n22569) );
  MUX41 U12055 ( .I0(ram[14234]), .I1(ram[14226]), .I2(ram[14218]), .I3(
        ram[14210]), .S0(n27136), .S1(n26661), .ZN(n22573) );
  MUX41 U12056 ( .I0(ram[14266]), .I1(ram[14258]), .I2(ram[14250]), .I3(
        ram[14242]), .S0(n27136), .S1(n26661), .ZN(n22571) );
  MUX41 U12057 ( .I0(ram[14330]), .I1(ram[14322]), .I2(ram[14314]), .I3(
        ram[14306]), .S0(n27137), .S1(n26662), .ZN(n22570) );
  MUX41 U12058 ( .I0(n22530), .I1(n22531), .I2(n22532), .I3(n22533), .S0(
        n26221), .S1(n26339), .ZN(n22529) );
  MUX41 U12059 ( .I0(ram[13210]), .I1(ram[13202]), .I2(ram[13194]), .I3(
        ram[13186]), .S0(n27134), .S1(n26659), .ZN(n22533) );
  MUX41 U12060 ( .I0(ram[13242]), .I1(ram[13234]), .I2(ram[13226]), .I3(
        ram[13218]), .S0(n27134), .S1(n26659), .ZN(n22531) );
  MUX41 U12061 ( .I0(ram[13306]), .I1(ram[13298]), .I2(ram[13290]), .I3(
        ram[13282]), .S0(n27134), .S1(n26659), .ZN(n22530) );
  MUX41 U12062 ( .I0(n22510), .I1(n22511), .I2(n22512), .I3(n22513), .S0(
        n26221), .S1(n26339), .ZN(n22509) );
  MUX41 U12063 ( .I0(ram[12698]), .I1(ram[12690]), .I2(ram[12682]), .I3(
        ram[12674]), .S0(n27133), .S1(n26658), .ZN(n22513) );
  MUX41 U12064 ( .I0(ram[12730]), .I1(ram[12722]), .I2(ram[12714]), .I3(
        ram[12706]), .S0(n27133), .S1(n26658), .ZN(n22511) );
  MUX41 U12065 ( .I0(ram[12794]), .I1(ram[12786]), .I2(ram[12778]), .I3(
        ram[12770]), .S0(n27133), .S1(n26658), .ZN(n22510) );
  MUX41 U12066 ( .I0(n22313), .I1(n22314), .I2(n22315), .I3(n22316), .S0(
        n26218), .S1(n26336), .ZN(n22312) );
  MUX41 U12067 ( .I0(ram[8122]), .I1(ram[8114]), .I2(ram[8106]), .I3(
        ram[8098]), .S0(n27122), .S1(n26647), .ZN(n22314) );
  MUX41 U12068 ( .I0(ram[8090]), .I1(ram[8082]), .I2(ram[8074]), .I3(
        ram[8066]), .S0(n27122), .S1(n26647), .ZN(n22316) );
  MUX41 U12069 ( .I0(ram[8186]), .I1(ram[8178]), .I2(ram[8170]), .I3(
        ram[8162]), .S0(n27122), .S1(n26647), .ZN(n22313) );
  MUX41 U12070 ( .I0(n22253), .I1(n22254), .I2(n22255), .I3(n22256), .S0(
        n26217), .S1(n26335), .ZN(n22252) );
  MUX41 U12071 ( .I0(ram[6554]), .I1(ram[6546]), .I2(ram[6538]), .I3(
        ram[6530]), .S0(n27118), .S1(n26643), .ZN(n22256) );
  MUX41 U12072 ( .I0(ram[6586]), .I1(ram[6578]), .I2(ram[6570]), .I3(
        ram[6562]), .S0(n27118), .S1(n26643), .ZN(n22254) );
  MUX41 U12073 ( .I0(ram[6650]), .I1(ram[6642]), .I2(ram[6634]), .I3(
        ram[6626]), .S0(n27118), .S1(n26643), .ZN(n22253) );
  MUX41 U12074 ( .I0(n22273), .I1(n22274), .I2(n22275), .I3(n22276), .S0(
        n26218), .S1(n26336), .ZN(n22272) );
  MUX41 U12075 ( .I0(ram[7066]), .I1(ram[7058]), .I2(ram[7050]), .I3(
        ram[7042]), .S0(n27119), .S1(n26644), .ZN(n22276) );
  MUX41 U12076 ( .I0(ram[7098]), .I1(ram[7090]), .I2(ram[7082]), .I3(
        ram[7074]), .S0(n27119), .S1(n26644), .ZN(n22274) );
  MUX41 U12077 ( .I0(ram[7162]), .I1(ram[7154]), .I2(ram[7146]), .I3(
        ram[7138]), .S0(n27119), .S1(n26644), .ZN(n22273) );
  MUX41 U12078 ( .I0(n22228), .I1(n22229), .I2(n22230), .I3(n22231), .S0(
        n26217), .S1(n26335), .ZN(n22227) );
  MUX41 U12079 ( .I0(ram[6074]), .I1(ram[6066]), .I2(ram[6058]), .I3(
        ram[6050]), .S0(n27117), .S1(n26642), .ZN(n22229) );
  MUX41 U12080 ( .I0(ram[6042]), .I1(ram[6034]), .I2(ram[6026]), .I3(
        ram[6018]), .S0(n27117), .S1(n26642), .ZN(n22231) );
  MUX41 U12081 ( .I0(ram[6138]), .I1(ram[6130]), .I2(ram[6122]), .I3(
        ram[6114]), .S0(n27117), .S1(n26642), .ZN(n22228) );
  MUX41 U12082 ( .I0(n22168), .I1(n22169), .I2(n22170), .I3(n22171), .S0(
        n26216), .S1(n26334), .ZN(n22167) );
  MUX41 U12083 ( .I0(ram[4538]), .I1(ram[4530]), .I2(ram[4522]), .I3(
        ram[4514]), .S0(n27113), .S1(n26638), .ZN(n22169) );
  MUX41 U12084 ( .I0(ram[4506]), .I1(ram[4498]), .I2(ram[4490]), .I3(
        ram[4482]), .S0(n27113), .S1(n26638), .ZN(n22171) );
  MUX41 U12085 ( .I0(ram[4602]), .I1(ram[4594]), .I2(ram[4586]), .I3(
        ram[4578]), .S0(n27113), .S1(n26638), .ZN(n22168) );
  MUX41 U12086 ( .I0(n22484), .I1(n22485), .I2(n22486), .I3(n22487), .S0(
        n26221), .S1(n26339), .ZN(n22483) );
  MUX41 U12087 ( .I0(ram[12218]), .I1(ram[12210]), .I2(ram[12202]), .I3(
        ram[12194]), .S0(n27132), .S1(n26657), .ZN(n22485) );
  MUX41 U12088 ( .I0(ram[12186]), .I1(ram[12178]), .I2(ram[12170]), .I3(
        ram[12162]), .S0(n27131), .S1(n26656), .ZN(n22487) );
  MUX41 U12089 ( .I0(ram[12282]), .I1(ram[12274]), .I2(ram[12266]), .I3(
        ram[12258]), .S0(n27132), .S1(n26657), .ZN(n22484) );
  MUX41 U12090 ( .I0(n22424), .I1(n22425), .I2(n22426), .I3(n22427), .S0(
        n26220), .S1(n26338), .ZN(n22423) );
  MUX41 U12091 ( .I0(ram[10682]), .I1(ram[10674]), .I2(ram[10666]), .I3(
        ram[10658]), .S0(n27128), .S1(n26653), .ZN(n22425) );
  MUX41 U12092 ( .I0(ram[10650]), .I1(ram[10642]), .I2(ram[10634]), .I3(
        ram[10626]), .S0(n27128), .S1(n26653), .ZN(n22427) );
  MUX41 U12093 ( .I0(ram[10746]), .I1(ram[10738]), .I2(ram[10730]), .I3(
        ram[10722]), .S0(n27128), .S1(n26653), .ZN(n22424) );
  MUX41 U12094 ( .I0(n22444), .I1(n22445), .I2(n22446), .I3(n22447), .S0(
        n26220), .S1(n26338), .ZN(n22443) );
  MUX41 U12095 ( .I0(ram[11194]), .I1(ram[11186]), .I2(ram[11178]), .I3(
        ram[11170]), .S0(n27129), .S1(n26654), .ZN(n22445) );
  MUX41 U12096 ( .I0(ram[11162]), .I1(ram[11154]), .I2(ram[11146]), .I3(
        ram[11138]), .S0(n27129), .S1(n26654), .ZN(n22447) );
  MUX41 U12097 ( .I0(ram[11258]), .I1(ram[11250]), .I2(ram[11242]), .I3(
        ram[11234]), .S0(n27129), .S1(n26654), .ZN(n22444) );
  MUX41 U12098 ( .I0(n22399), .I1(n22400), .I2(n22401), .I3(n22402), .S0(
        n26220), .S1(n26338), .ZN(n22398) );
  MUX41 U12099 ( .I0(ram[10170]), .I1(ram[10162]), .I2(ram[10154]), .I3(
        ram[10146]), .S0(n27127), .S1(n26652), .ZN(n22400) );
  MUX41 U12100 ( .I0(ram[10138]), .I1(ram[10130]), .I2(ram[10122]), .I3(
        ram[10114]), .S0(n27127), .S1(n26652), .ZN(n22402) );
  MUX41 U12101 ( .I0(ram[10234]), .I1(ram[10226]), .I2(ram[10218]), .I3(
        ram[10210]), .S0(n27127), .S1(n26652), .ZN(n22399) );
  MUX41 U12102 ( .I0(n22339), .I1(n22340), .I2(n22341), .I3(n22342), .S0(
        n26219), .S1(n26337), .ZN(n22338) );
  MUX41 U12103 ( .I0(ram[8634]), .I1(ram[8626]), .I2(ram[8618]), .I3(
        ram[8610]), .S0(n27123), .S1(n26648), .ZN(n22340) );
  MUX41 U12104 ( .I0(ram[8602]), .I1(ram[8594]), .I2(ram[8586]), .I3(
        ram[8578]), .S0(n27123), .S1(n26648), .ZN(n22342) );
  MUX41 U12105 ( .I0(ram[8698]), .I1(ram[8690]), .I2(ram[8682]), .I3(
        ram[8674]), .S0(n27123), .S1(n26648), .ZN(n22339) );
  MUX41 U12106 ( .I0(n22359), .I1(n22360), .I2(n22361), .I3(n22362), .S0(
        n26219), .S1(n26337), .ZN(n22358) );
  MUX41 U12107 ( .I0(ram[9114]), .I1(ram[9106]), .I2(ram[9098]), .I3(
        ram[9090]), .S0(n27124), .S1(n26649), .ZN(n22362) );
  MUX41 U12108 ( .I0(ram[9146]), .I1(ram[9138]), .I2(ram[9130]), .I3(
        ram[9122]), .S0(n27124), .S1(n26649), .ZN(n22360) );
  MUX41 U12109 ( .I0(ram[9210]), .I1(ram[9202]), .I2(ram[9194]), .I3(
        ram[9186]), .S0(n27124), .S1(n26649), .ZN(n22359) );
  MUX41 U12110 ( .I0(n23339), .I1(n23340), .I2(n23341), .I3(n23342), .S0(
        n26233), .S1(n26351), .ZN(n23338) );
  MUX41 U12111 ( .I0(ram[16283]), .I1(ram[16275]), .I2(ram[16267]), .I3(
        ram[16259]), .S0(n27181), .S1(n26706), .ZN(n23342) );
  MUX41 U12112 ( .I0(ram[16315]), .I1(ram[16307]), .I2(ram[16299]), .I3(
        ram[16291]), .S0(n27181), .S1(n26706), .ZN(n23340) );
  MUX41 U12113 ( .I0(ram[16379]), .I1(ram[16371]), .I2(ram[16363]), .I3(
        ram[16355]), .S0(n27181), .S1(n26706), .ZN(n23339) );
  MUX41 U12114 ( .I0(n23299), .I1(n23300), .I2(n23301), .I3(n23302), .S0(
        n26232), .S1(n26350), .ZN(n23298) );
  MUX41 U12115 ( .I0(ram[15259]), .I1(ram[15251]), .I2(ram[15243]), .I3(
        ram[15235]), .S0(n27178), .S1(n26703), .ZN(n23302) );
  MUX41 U12116 ( .I0(ram[15291]), .I1(ram[15283]), .I2(ram[15275]), .I3(
        ram[15267]), .S0(n27178), .S1(n26703), .ZN(n23300) );
  MUX41 U12117 ( .I0(ram[15355]), .I1(ram[15347]), .I2(ram[15339]), .I3(
        ram[15331]), .S0(n27178), .S1(n26703), .ZN(n23299) );
  MUX41 U12118 ( .I0(n23279), .I1(n23280), .I2(n23281), .I3(n23282), .S0(
        n26232), .S1(n26350), .ZN(n23278) );
  MUX41 U12119 ( .I0(ram[14747]), .I1(ram[14739]), .I2(ram[14731]), .I3(
        ram[14723]), .S0(n27177), .S1(n26702), .ZN(n23282) );
  MUX41 U12120 ( .I0(ram[14779]), .I1(ram[14771]), .I2(ram[14763]), .I3(
        ram[14755]), .S0(n27177), .S1(n26702), .ZN(n23280) );
  MUX41 U12121 ( .I0(ram[14843]), .I1(ram[14835]), .I2(ram[14827]), .I3(
        ram[14819]), .S0(n27177), .S1(n26702), .ZN(n23279) );
  MUX41 U12122 ( .I0(n23254), .I1(n23255), .I2(n23256), .I3(n23257), .S0(
        n26232), .S1(n26350), .ZN(n23253) );
  MUX41 U12123 ( .I0(ram[14235]), .I1(ram[14227]), .I2(ram[14219]), .I3(
        ram[14211]), .S0(n27176), .S1(n26701), .ZN(n23257) );
  MUX41 U12124 ( .I0(ram[14267]), .I1(ram[14259]), .I2(ram[14251]), .I3(
        ram[14243]), .S0(n27176), .S1(n26701), .ZN(n23255) );
  MUX41 U12125 ( .I0(ram[14331]), .I1(ram[14323]), .I2(ram[14315]), .I3(
        ram[14307]), .S0(n27176), .S1(n26701), .ZN(n23254) );
  MUX41 U12126 ( .I0(n23214), .I1(n23215), .I2(n23216), .I3(n23217), .S0(
        n26231), .S1(n26349), .ZN(n23213) );
  MUX41 U12127 ( .I0(ram[13211]), .I1(ram[13203]), .I2(ram[13195]), .I3(
        ram[13187]), .S0(n27173), .S1(n26698), .ZN(n23217) );
  MUX41 U12128 ( .I0(ram[13243]), .I1(ram[13235]), .I2(ram[13227]), .I3(
        ram[13219]), .S0(n27173), .S1(n26698), .ZN(n23215) );
  MUX41 U12129 ( .I0(ram[13307]), .I1(ram[13299]), .I2(ram[13291]), .I3(
        ram[13283]), .S0(n27174), .S1(n26699), .ZN(n23214) );
  MUX41 U12130 ( .I0(n23194), .I1(n23195), .I2(n23196), .I3(n23197), .S0(
        n26231), .S1(n26349), .ZN(n23193) );
  MUX41 U12131 ( .I0(ram[12699]), .I1(ram[12691]), .I2(ram[12683]), .I3(
        ram[12675]), .S0(n27172), .S1(n26697), .ZN(n23197) );
  MUX41 U12132 ( .I0(ram[12731]), .I1(ram[12723]), .I2(ram[12715]), .I3(
        ram[12707]), .S0(n27172), .S1(n26697), .ZN(n23195) );
  MUX41 U12133 ( .I0(ram[12795]), .I1(ram[12787]), .I2(ram[12779]), .I3(
        ram[12771]), .S0(n27172), .S1(n26697), .ZN(n23194) );
  MUX41 U12134 ( .I0(n22997), .I1(n22998), .I2(n22999), .I3(n23000), .S0(
        n26228), .S1(n26346), .ZN(n22996) );
  MUX41 U12135 ( .I0(ram[8123]), .I1(ram[8115]), .I2(ram[8107]), .I3(
        ram[8099]), .S0(n27161), .S1(n26686), .ZN(n22998) );
  MUX41 U12136 ( .I0(ram[8091]), .I1(ram[8083]), .I2(ram[8075]), .I3(
        ram[8067]), .S0(n27161), .S1(n26686), .ZN(n23000) );
  MUX41 U12137 ( .I0(ram[8187]), .I1(ram[8179]), .I2(ram[8171]), .I3(
        ram[8163]), .S0(n27161), .S1(n26686), .ZN(n22997) );
  MUX41 U12138 ( .I0(n22937), .I1(n22938), .I2(n22939), .I3(n22940), .S0(
        n26227), .S1(n26345), .ZN(n22936) );
  MUX41 U12139 ( .I0(ram[6555]), .I1(ram[6547]), .I2(ram[6539]), .I3(
        ram[6531]), .S0(n27157), .S1(n26682), .ZN(n22940) );
  MUX41 U12140 ( .I0(ram[6587]), .I1(ram[6579]), .I2(ram[6571]), .I3(
        ram[6563]), .S0(n27157), .S1(n26682), .ZN(n22938) );
  MUX41 U12141 ( .I0(ram[6651]), .I1(ram[6643]), .I2(ram[6635]), .I3(
        ram[6627]), .S0(n27158), .S1(n26683), .ZN(n22937) );
  MUX41 U12142 ( .I0(n22957), .I1(n22958), .I2(n22959), .I3(n22960), .S0(
        n26228), .S1(n26346), .ZN(n22956) );
  MUX41 U12143 ( .I0(ram[7067]), .I1(ram[7059]), .I2(ram[7051]), .I3(
        ram[7043]), .S0(n27159), .S1(n26684), .ZN(n22960) );
  MUX41 U12144 ( .I0(ram[7099]), .I1(ram[7091]), .I2(ram[7083]), .I3(
        ram[7075]), .S0(n27159), .S1(n26684), .ZN(n22958) );
  MUX41 U12145 ( .I0(ram[7163]), .I1(ram[7155]), .I2(ram[7147]), .I3(
        ram[7139]), .S0(n27159), .S1(n26684), .ZN(n22957) );
  MUX41 U12146 ( .I0(n22912), .I1(n22913), .I2(n22914), .I3(n22915), .S0(
        n26227), .S1(n26345), .ZN(n22911) );
  MUX41 U12147 ( .I0(ram[6075]), .I1(ram[6067]), .I2(ram[6059]), .I3(
        ram[6051]), .S0(n27156), .S1(n26681), .ZN(n22913) );
  MUX41 U12148 ( .I0(ram[6043]), .I1(ram[6035]), .I2(ram[6027]), .I3(
        ram[6019]), .S0(n27156), .S1(n26681), .ZN(n22915) );
  MUX41 U12149 ( .I0(ram[6139]), .I1(ram[6131]), .I2(ram[6123]), .I3(
        ram[6115]), .S0(n27156), .S1(n26681), .ZN(n22912) );
  MUX41 U12150 ( .I0(n22852), .I1(n22853), .I2(n22854), .I3(n22855), .S0(
        n26226), .S1(n26344), .ZN(n22851) );
  MUX41 U12151 ( .I0(ram[4539]), .I1(ram[4531]), .I2(ram[4523]), .I3(
        ram[4515]), .S0(n27152), .S1(n26677), .ZN(n22853) );
  MUX41 U12152 ( .I0(ram[4507]), .I1(ram[4499]), .I2(ram[4491]), .I3(
        ram[4483]), .S0(n27152), .S1(n26677), .ZN(n22855) );
  MUX41 U12153 ( .I0(ram[4603]), .I1(ram[4595]), .I2(ram[4587]), .I3(
        ram[4579]), .S0(n27153), .S1(n26678), .ZN(n22852) );
  MUX41 U12154 ( .I0(n23168), .I1(n23169), .I2(n23170), .I3(n23171), .S0(
        n26231), .S1(n26349), .ZN(n23167) );
  MUX41 U12155 ( .I0(ram[12219]), .I1(ram[12211]), .I2(ram[12203]), .I3(
        ram[12195]), .S0(n27171), .S1(n26696), .ZN(n23169) );
  MUX41 U12156 ( .I0(ram[12187]), .I1(ram[12179]), .I2(ram[12171]), .I3(
        ram[12163]), .S0(n27171), .S1(n26696), .ZN(n23171) );
  MUX41 U12157 ( .I0(ram[12283]), .I1(ram[12275]), .I2(ram[12267]), .I3(
        ram[12259]), .S0(n27171), .S1(n26696), .ZN(n23168) );
  MUX41 U12158 ( .I0(n23108), .I1(n23109), .I2(n23110), .I3(n23111), .S0(
        n26230), .S1(n26348), .ZN(n23107) );
  MUX41 U12159 ( .I0(ram[10683]), .I1(ram[10675]), .I2(ram[10667]), .I3(
        ram[10659]), .S0(n27167), .S1(n26692), .ZN(n23109) );
  MUX41 U12160 ( .I0(ram[10651]), .I1(ram[10643]), .I2(ram[10635]), .I3(
        ram[10627]), .S0(n27167), .S1(n26692), .ZN(n23111) );
  MUX41 U12161 ( .I0(ram[10747]), .I1(ram[10739]), .I2(ram[10731]), .I3(
        ram[10723]), .S0(n27167), .S1(n26692), .ZN(n23108) );
  MUX41 U12162 ( .I0(n23128), .I1(n23129), .I2(n23130), .I3(n23131), .S0(
        n26230), .S1(n26348), .ZN(n23127) );
  MUX41 U12163 ( .I0(ram[11195]), .I1(ram[11187]), .I2(ram[11179]), .I3(
        ram[11171]), .S0(n27168), .S1(n26693), .ZN(n23129) );
  MUX41 U12164 ( .I0(ram[11163]), .I1(ram[11155]), .I2(ram[11147]), .I3(
        ram[11139]), .S0(n27168), .S1(n26693), .ZN(n23131) );
  MUX41 U12165 ( .I0(ram[11259]), .I1(ram[11251]), .I2(ram[11243]), .I3(
        ram[11235]), .S0(n27169), .S1(n26694), .ZN(n23128) );
  MUX41 U12166 ( .I0(n23083), .I1(n23084), .I2(n23085), .I3(n23086), .S0(
        n26229), .S1(n26347), .ZN(n23082) );
  MUX41 U12167 ( .I0(ram[10171]), .I1(ram[10163]), .I2(ram[10155]), .I3(
        ram[10147]), .S0(n27166), .S1(n26691), .ZN(n23084) );
  MUX41 U12168 ( .I0(ram[10139]), .I1(ram[10131]), .I2(ram[10123]), .I3(
        ram[10115]), .S0(n27166), .S1(n26691), .ZN(n23086) );
  MUX41 U12169 ( .I0(ram[10235]), .I1(ram[10227]), .I2(ram[10219]), .I3(
        ram[10211]), .S0(n27166), .S1(n26691), .ZN(n23083) );
  MUX41 U12170 ( .I0(n23023), .I1(n23024), .I2(n23025), .I3(n23026), .S0(
        n26228), .S1(n26346), .ZN(n23022) );
  MUX41 U12171 ( .I0(ram[8635]), .I1(ram[8627]), .I2(ram[8619]), .I3(
        ram[8611]), .S0(n27162), .S1(n26687), .ZN(n23024) );
  MUX41 U12172 ( .I0(ram[8603]), .I1(ram[8595]), .I2(ram[8587]), .I3(
        ram[8579]), .S0(n27162), .S1(n26687), .ZN(n23026) );
  MUX41 U12173 ( .I0(ram[8699]), .I1(ram[8691]), .I2(ram[8683]), .I3(
        ram[8675]), .S0(n27162), .S1(n26687), .ZN(n23023) );
  MUX41 U12174 ( .I0(n23043), .I1(n23044), .I2(n23045), .I3(n23046), .S0(
        n26229), .S1(n26347), .ZN(n23042) );
  MUX41 U12175 ( .I0(ram[9115]), .I1(ram[9107]), .I2(ram[9099]), .I3(
        ram[9091]), .S0(n27163), .S1(n26688), .ZN(n23046) );
  MUX41 U12176 ( .I0(ram[9147]), .I1(ram[9139]), .I2(ram[9131]), .I3(
        ram[9123]), .S0(n27164), .S1(n26689), .ZN(n23044) );
  MUX41 U12177 ( .I0(ram[9211]), .I1(ram[9203]), .I2(ram[9195]), .I3(
        ram[9187]), .S0(n27164), .S1(n26689), .ZN(n23043) );
  MUX41 U12178 ( .I0(n24023), .I1(n24024), .I2(n24025), .I3(n24026), .S0(
        n26243), .S1(n26361), .ZN(n24022) );
  MUX41 U12179 ( .I0(ram[16284]), .I1(ram[16276]), .I2(ram[16268]), .I3(
        ram[16260]), .S0(n27220), .S1(n26745), .ZN(n24026) );
  MUX41 U12180 ( .I0(ram[16316]), .I1(ram[16308]), .I2(ram[16300]), .I3(
        ram[16292]), .S0(n27220), .S1(n26745), .ZN(n24024) );
  MUX41 U12181 ( .I0(ram[16380]), .I1(ram[16372]), .I2(ram[16364]), .I3(
        ram[16356]), .S0(n27220), .S1(n26745), .ZN(n24023) );
  MUX41 U12182 ( .I0(n23983), .I1(n23984), .I2(n23985), .I3(n23986), .S0(
        n26242), .S1(n26360), .ZN(n23982) );
  MUX41 U12183 ( .I0(ram[15260]), .I1(ram[15252]), .I2(ram[15244]), .I3(
        ram[15236]), .S0(n27218), .S1(n26743), .ZN(n23986) );
  MUX41 U12184 ( .I0(ram[15292]), .I1(ram[15284]), .I2(ram[15276]), .I3(
        ram[15268]), .S0(n27218), .S1(n26743), .ZN(n23984) );
  MUX41 U12185 ( .I0(ram[15356]), .I1(ram[15348]), .I2(ram[15340]), .I3(
        ram[15332]), .S0(n27218), .S1(n26743), .ZN(n23983) );
  MUX41 U12186 ( .I0(n23963), .I1(n23964), .I2(n23965), .I3(n23966), .S0(
        n26242), .S1(n26360), .ZN(n23962) );
  MUX41 U12187 ( .I0(ram[14748]), .I1(ram[14740]), .I2(ram[14732]), .I3(
        ram[14724]), .S0(n27216), .S1(n26741), .ZN(n23966) );
  MUX41 U12188 ( .I0(ram[14780]), .I1(ram[14772]), .I2(ram[14764]), .I3(
        ram[14756]), .S0(n27216), .S1(n26741), .ZN(n23964) );
  MUX41 U12189 ( .I0(ram[14844]), .I1(ram[14836]), .I2(ram[14828]), .I3(
        ram[14820]), .S0(n27217), .S1(n26742), .ZN(n23963) );
  MUX41 U12190 ( .I0(n23938), .I1(n23939), .I2(n23940), .I3(n23941), .S0(
        n26242), .S1(n26360), .ZN(n23937) );
  MUX41 U12191 ( .I0(ram[14236]), .I1(ram[14228]), .I2(ram[14220]), .I3(
        ram[14212]), .S0(n27215), .S1(n26740), .ZN(n23941) );
  MUX41 U12192 ( .I0(ram[14268]), .I1(ram[14260]), .I2(ram[14252]), .I3(
        ram[14244]), .S0(n27215), .S1(n26740), .ZN(n23939) );
  MUX41 U12193 ( .I0(ram[14332]), .I1(ram[14324]), .I2(ram[14316]), .I3(
        ram[14308]), .S0(n27215), .S1(n26740), .ZN(n23938) );
  MUX41 U12194 ( .I0(n23898), .I1(n23899), .I2(n23900), .I3(n23901), .S0(
        n26241), .S1(n26359), .ZN(n23897) );
  MUX41 U12195 ( .I0(ram[13212]), .I1(ram[13204]), .I2(ram[13196]), .I3(
        ram[13188]), .S0(n27213), .S1(n26738), .ZN(n23901) );
  MUX41 U12196 ( .I0(ram[13244]), .I1(ram[13236]), .I2(ram[13228]), .I3(
        ram[13220]), .S0(n27213), .S1(n26738), .ZN(n23899) );
  MUX41 U12197 ( .I0(ram[13308]), .I1(ram[13300]), .I2(ram[13292]), .I3(
        ram[13284]), .S0(n27213), .S1(n26738), .ZN(n23898) );
  MUX41 U12198 ( .I0(n23878), .I1(n23879), .I2(n23880), .I3(n23881), .S0(
        n26241), .S1(n26359), .ZN(n23877) );
  MUX41 U12199 ( .I0(ram[12700]), .I1(ram[12692]), .I2(ram[12684]), .I3(
        ram[12676]), .S0(n27211), .S1(n26736), .ZN(n23881) );
  MUX41 U12200 ( .I0(ram[12732]), .I1(ram[12724]), .I2(ram[12716]), .I3(
        ram[12708]), .S0(n27212), .S1(n26737), .ZN(n23879) );
  MUX41 U12201 ( .I0(ram[12796]), .I1(ram[12788]), .I2(ram[12780]), .I3(
        ram[12772]), .S0(n27212), .S1(n26737), .ZN(n23878) );
  MUX41 U12202 ( .I0(n23681), .I1(n23682), .I2(n23683), .I3(n23684), .S0(
        n26238), .S1(n26356), .ZN(n23680) );
  MUX41 U12203 ( .I0(ram[8124]), .I1(ram[8116]), .I2(ram[8108]), .I3(
        ram[8100]), .S0(n27200), .S1(n26725), .ZN(n23682) );
  MUX41 U12204 ( .I0(ram[8092]), .I1(ram[8084]), .I2(ram[8076]), .I3(
        ram[8068]), .S0(n27200), .S1(n26725), .ZN(n23684) );
  MUX41 U12205 ( .I0(ram[8188]), .I1(ram[8180]), .I2(ram[8172]), .I3(
        ram[8164]), .S0(n27201), .S1(n26726), .ZN(n23681) );
  MUX41 U12206 ( .I0(n23621), .I1(n23622), .I2(n23623), .I3(n23624), .S0(
        n26237), .S1(n26355), .ZN(n23620) );
  MUX41 U12207 ( .I0(ram[6556]), .I1(ram[6548]), .I2(ram[6540]), .I3(
        ram[6532]), .S0(n27197), .S1(n26722), .ZN(n23624) );
  MUX41 U12208 ( .I0(ram[6588]), .I1(ram[6580]), .I2(ram[6572]), .I3(
        ram[6564]), .S0(n27197), .S1(n26722), .ZN(n23622) );
  MUX41 U12209 ( .I0(ram[6652]), .I1(ram[6644]), .I2(ram[6636]), .I3(
        ram[6628]), .S0(n27197), .S1(n26722), .ZN(n23621) );
  MUX41 U12210 ( .I0(n23641), .I1(n23642), .I2(n23643), .I3(n23644), .S0(
        n26237), .S1(n26355), .ZN(n23640) );
  MUX41 U12211 ( .I0(ram[7068]), .I1(ram[7060]), .I2(ram[7052]), .I3(
        ram[7044]), .S0(n27198), .S1(n26723), .ZN(n23644) );
  MUX41 U12212 ( .I0(ram[7100]), .I1(ram[7092]), .I2(ram[7084]), .I3(
        ram[7076]), .S0(n27198), .S1(n26723), .ZN(n23642) );
  MUX41 U12213 ( .I0(ram[7164]), .I1(ram[7156]), .I2(ram[7148]), .I3(
        ram[7140]), .S0(n27198), .S1(n26723), .ZN(n23641) );
  MUX41 U12214 ( .I0(n23596), .I1(n23597), .I2(n23598), .I3(n23599), .S0(
        n26237), .S1(n26355), .ZN(n23595) );
  MUX41 U12215 ( .I0(ram[6076]), .I1(ram[6068]), .I2(ram[6060]), .I3(
        ram[6052]), .S0(n27196), .S1(n26721), .ZN(n23597) );
  MUX41 U12216 ( .I0(ram[6044]), .I1(ram[6036]), .I2(ram[6028]), .I3(
        ram[6020]), .S0(n27195), .S1(n26720), .ZN(n23599) );
  MUX41 U12217 ( .I0(ram[6140]), .I1(ram[6132]), .I2(ram[6124]), .I3(
        ram[6116]), .S0(n27196), .S1(n26721), .ZN(n23596) );
  MUX41 U12218 ( .I0(n23536), .I1(n23537), .I2(n23538), .I3(n23539), .S0(
        n26236), .S1(n26354), .ZN(n23535) );
  MUX41 U12219 ( .I0(ram[4540]), .I1(ram[4532]), .I2(ram[4524]), .I3(
        ram[4516]), .S0(n27192), .S1(n26717), .ZN(n23537) );
  MUX41 U12220 ( .I0(ram[4508]), .I1(ram[4500]), .I2(ram[4492]), .I3(
        ram[4484]), .S0(n27192), .S1(n26717), .ZN(n23539) );
  MUX41 U12221 ( .I0(ram[4604]), .I1(ram[4596]), .I2(ram[4588]), .I3(
        ram[4580]), .S0(n27192), .S1(n26717), .ZN(n23536) );
  MUX41 U12222 ( .I0(n23852), .I1(n23853), .I2(n23854), .I3(n23855), .S0(
        n26240), .S1(n26358), .ZN(n23851) );
  MUX41 U12223 ( .I0(ram[12220]), .I1(ram[12212]), .I2(ram[12204]), .I3(
        ram[12196]), .S0(n27210), .S1(n26735), .ZN(n23853) );
  MUX41 U12224 ( .I0(ram[12188]), .I1(ram[12180]), .I2(ram[12172]), .I3(
        ram[12164]), .S0(n27210), .S1(n26735), .ZN(n23855) );
  MUX41 U12225 ( .I0(ram[12284]), .I1(ram[12276]), .I2(ram[12268]), .I3(
        ram[12260]), .S0(n27210), .S1(n26735), .ZN(n23852) );
  MUX41 U12226 ( .I0(n23792), .I1(n23793), .I2(n23794), .I3(n23795), .S0(
        n26240), .S1(n26358), .ZN(n23791) );
  MUX41 U12227 ( .I0(ram[10684]), .I1(ram[10676]), .I2(ram[10668]), .I3(
        ram[10660]), .S0(n27207), .S1(n26732), .ZN(n23793) );
  MUX41 U12228 ( .I0(ram[10652]), .I1(ram[10644]), .I2(ram[10636]), .I3(
        ram[10628]), .S0(n27207), .S1(n26732), .ZN(n23795) );
  MUX41 U12229 ( .I0(ram[10748]), .I1(ram[10740]), .I2(ram[10732]), .I3(
        ram[10724]), .S0(n27207), .S1(n26732), .ZN(n23792) );
  MUX41 U12230 ( .I0(n23812), .I1(n23813), .I2(n23814), .I3(n23815), .S0(
        n26240), .S1(n26358), .ZN(n23811) );
  MUX41 U12231 ( .I0(ram[11196]), .I1(ram[11188]), .I2(ram[11180]), .I3(
        ram[11172]), .S0(n27208), .S1(n26733), .ZN(n23813) );
  MUX41 U12232 ( .I0(ram[11164]), .I1(ram[11156]), .I2(ram[11148]), .I3(
        ram[11140]), .S0(n27208), .S1(n26733), .ZN(n23815) );
  MUX41 U12233 ( .I0(ram[11260]), .I1(ram[11252]), .I2(ram[11244]), .I3(
        ram[11236]), .S0(n27208), .S1(n26733), .ZN(n23812) );
  MUX41 U12234 ( .I0(n23767), .I1(n23768), .I2(n23769), .I3(n23770), .S0(
        n26239), .S1(n26357), .ZN(n23766) );
  MUX41 U12235 ( .I0(ram[10172]), .I1(ram[10164]), .I2(ram[10156]), .I3(
        ram[10148]), .S0(n27205), .S1(n26730), .ZN(n23768) );
  MUX41 U12236 ( .I0(ram[10140]), .I1(ram[10132]), .I2(ram[10124]), .I3(
        ram[10116]), .S0(n27205), .S1(n26730), .ZN(n23770) );
  MUX41 U12237 ( .I0(ram[10236]), .I1(ram[10228]), .I2(ram[10220]), .I3(
        ram[10212]), .S0(n27206), .S1(n26731), .ZN(n23767) );
  MUX41 U12238 ( .I0(n23707), .I1(n23708), .I2(n23709), .I3(n23710), .S0(
        n26238), .S1(n26356), .ZN(n23706) );
  MUX41 U12239 ( .I0(ram[8636]), .I1(ram[8628]), .I2(ram[8620]), .I3(
        ram[8612]), .S0(n27202), .S1(n26727), .ZN(n23708) );
  MUX41 U12240 ( .I0(ram[8604]), .I1(ram[8596]), .I2(ram[8588]), .I3(
        ram[8580]), .S0(n27202), .S1(n26727), .ZN(n23710) );
  MUX41 U12241 ( .I0(ram[8700]), .I1(ram[8692]), .I2(ram[8684]), .I3(
        ram[8676]), .S0(n27202), .S1(n26727), .ZN(n23707) );
  MUX41 U12242 ( .I0(n23727), .I1(n23728), .I2(n23729), .I3(n23730), .S0(
        n26239), .S1(n26357), .ZN(n23726) );
  MUX41 U12243 ( .I0(ram[9116]), .I1(ram[9108]), .I2(ram[9100]), .I3(
        ram[9092]), .S0(n27203), .S1(n26728), .ZN(n23730) );
  MUX41 U12244 ( .I0(ram[9148]), .I1(ram[9140]), .I2(ram[9132]), .I3(
        ram[9124]), .S0(n27203), .S1(n26728), .ZN(n23728) );
  MUX41 U12245 ( .I0(ram[9212]), .I1(ram[9204]), .I2(ram[9196]), .I3(
        ram[9188]), .S0(n27203), .S1(n26728), .ZN(n23727) );
  MUX41 U12246 ( .I0(n24707), .I1(n24708), .I2(n24709), .I3(n24710), .S0(
        n26253), .S1(n26371), .ZN(n24706) );
  MUX41 U12247 ( .I0(ram[16285]), .I1(ram[16277]), .I2(ram[16269]), .I3(
        ram[16261]), .S0(n27259), .S1(n26784), .ZN(n24710) );
  MUX41 U12248 ( .I0(ram[16317]), .I1(ram[16309]), .I2(ram[16301]), .I3(
        ram[16293]), .S0(n27260), .S1(n26785), .ZN(n24708) );
  MUX41 U12249 ( .I0(ram[16381]), .I1(ram[16373]), .I2(ram[16365]), .I3(
        ram[16357]), .S0(n27260), .S1(n26785), .ZN(n24707) );
  MUX41 U12250 ( .I0(n24667), .I1(n24668), .I2(n24669), .I3(n24670), .S0(
        n26252), .S1(n26370), .ZN(n24666) );
  MUX41 U12251 ( .I0(ram[15261]), .I1(ram[15253]), .I2(ram[15245]), .I3(
        ram[15237]), .S0(n27257), .S1(n26782), .ZN(n24670) );
  MUX41 U12252 ( .I0(ram[15293]), .I1(ram[15285]), .I2(ram[15277]), .I3(
        ram[15269]), .S0(n27257), .S1(n26782), .ZN(n24668) );
  MUX41 U12253 ( .I0(ram[15357]), .I1(ram[15349]), .I2(ram[15341]), .I3(
        ram[15333]), .S0(n27257), .S1(n26782), .ZN(n24667) );
  MUX41 U12254 ( .I0(n24647), .I1(n24648), .I2(n24649), .I3(n24650), .S0(
        n26252), .S1(n26370), .ZN(n24646) );
  MUX41 U12255 ( .I0(ram[14749]), .I1(ram[14741]), .I2(ram[14733]), .I3(
        ram[14725]), .S0(n27256), .S1(n26781), .ZN(n24650) );
  MUX41 U12256 ( .I0(ram[14781]), .I1(ram[14773]), .I2(ram[14765]), .I3(
        ram[14757]), .S0(n27256), .S1(n26781), .ZN(n24648) );
  MUX41 U12257 ( .I0(ram[14845]), .I1(ram[14837]), .I2(ram[14829]), .I3(
        ram[14821]), .S0(n27256), .S1(n26781), .ZN(n24647) );
  MUX41 U12258 ( .I0(n24622), .I1(n24623), .I2(n24624), .I3(n24625), .S0(
        n26252), .S1(n26370), .ZN(n24621) );
  MUX41 U12259 ( .I0(ram[14237]), .I1(ram[14229]), .I2(ram[14221]), .I3(
        ram[14213]), .S0(n27255), .S1(n26780), .ZN(n24625) );
  MUX41 U12260 ( .I0(ram[14269]), .I1(ram[14261]), .I2(ram[14253]), .I3(
        ram[14245]), .S0(n27255), .S1(n26780), .ZN(n24623) );
  MUX41 U12261 ( .I0(ram[14333]), .I1(ram[14325]), .I2(ram[14317]), .I3(
        ram[14309]), .S0(n27255), .S1(n26780), .ZN(n24622) );
  MUX41 U12262 ( .I0(n24582), .I1(n24583), .I2(n24584), .I3(n24585), .S0(
        n26251), .S1(n26369), .ZN(n24581) );
  MUX41 U12263 ( .I0(ram[13213]), .I1(ram[13205]), .I2(ram[13197]), .I3(
        ram[13189]), .S0(n27252), .S1(n26777), .ZN(n24585) );
  MUX41 U12264 ( .I0(ram[13245]), .I1(ram[13237]), .I2(ram[13229]), .I3(
        ram[13221]), .S0(n27252), .S1(n26777), .ZN(n24583) );
  MUX41 U12265 ( .I0(ram[13309]), .I1(ram[13301]), .I2(ram[13293]), .I3(
        ram[13285]), .S0(n27252), .S1(n26777), .ZN(n24582) );
  MUX41 U12266 ( .I0(n24562), .I1(n24563), .I2(n24564), .I3(n24565), .S0(
        n26251), .S1(n26369), .ZN(n24561) );
  MUX41 U12267 ( .I0(ram[12701]), .I1(ram[12693]), .I2(ram[12685]), .I3(
        ram[12677]), .S0(n27251), .S1(n26776), .ZN(n24565) );
  MUX41 U12268 ( .I0(ram[12733]), .I1(ram[12725]), .I2(ram[12717]), .I3(
        ram[12709]), .S0(n27251), .S1(n26776), .ZN(n24563) );
  MUX41 U12269 ( .I0(ram[12797]), .I1(ram[12789]), .I2(ram[12781]), .I3(
        ram[12773]), .S0(n27251), .S1(n26776), .ZN(n24562) );
  MUX41 U12270 ( .I0(n24365), .I1(n24366), .I2(n24367), .I3(n24368), .S0(
        n26248), .S1(n26366), .ZN(n24364) );
  MUX41 U12271 ( .I0(ram[8125]), .I1(ram[8117]), .I2(ram[8109]), .I3(
        ram[8101]), .S0(n27240), .S1(n26765), .ZN(n24366) );
  MUX41 U12272 ( .I0(ram[8093]), .I1(ram[8085]), .I2(ram[8077]), .I3(
        ram[8069]), .S0(n27240), .S1(n26765), .ZN(n24368) );
  MUX41 U12273 ( .I0(ram[8189]), .I1(ram[8181]), .I2(ram[8173]), .I3(
        ram[8165]), .S0(n27240), .S1(n26765), .ZN(n24365) );
  MUX41 U12274 ( .I0(n24305), .I1(n24306), .I2(n24307), .I3(n24308), .S0(
        n26247), .S1(n26365), .ZN(n24304) );
  MUX41 U12275 ( .I0(ram[6557]), .I1(ram[6549]), .I2(ram[6541]), .I3(
        ram[6533]), .S0(n27236), .S1(n26761), .ZN(n24308) );
  MUX41 U12276 ( .I0(ram[6589]), .I1(ram[6581]), .I2(ram[6573]), .I3(
        ram[6565]), .S0(n27236), .S1(n26761), .ZN(n24306) );
  MUX41 U12277 ( .I0(ram[6653]), .I1(ram[6645]), .I2(ram[6637]), .I3(
        ram[6629]), .S0(n27236), .S1(n26761), .ZN(n24305) );
  MUX41 U12278 ( .I0(n24325), .I1(n24326), .I2(n24327), .I3(n24328), .S0(
        n26247), .S1(n26365), .ZN(n24324) );
  MUX41 U12279 ( .I0(ram[7069]), .I1(ram[7061]), .I2(ram[7053]), .I3(
        ram[7045]), .S0(n27237), .S1(n26762), .ZN(n24328) );
  MUX41 U12280 ( .I0(ram[7101]), .I1(ram[7093]), .I2(ram[7085]), .I3(
        ram[7077]), .S0(n27237), .S1(n26762), .ZN(n24326) );
  MUX41 U12281 ( .I0(ram[7165]), .I1(ram[7157]), .I2(ram[7149]), .I3(
        ram[7141]), .S0(n27238), .S1(n26763), .ZN(n24325) );
  MUX41 U12282 ( .I0(n24280), .I1(n24281), .I2(n24282), .I3(n24283), .S0(
        n26247), .S1(n26365), .ZN(n24279) );
  MUX41 U12283 ( .I0(ram[6077]), .I1(ram[6069]), .I2(ram[6061]), .I3(
        ram[6053]), .S0(n27235), .S1(n26760), .ZN(n24281) );
  MUX41 U12284 ( .I0(ram[6045]), .I1(ram[6037]), .I2(ram[6029]), .I3(
        ram[6021]), .S0(n27235), .S1(n26760), .ZN(n24283) );
  MUX41 U12285 ( .I0(ram[6141]), .I1(ram[6133]), .I2(ram[6125]), .I3(
        ram[6117]), .S0(n27235), .S1(n26760), .ZN(n24280) );
  MUX41 U12286 ( .I0(n24220), .I1(n24221), .I2(n24222), .I3(n24223), .S0(
        n26246), .S1(n26364), .ZN(n24219) );
  MUX41 U12287 ( .I0(ram[4541]), .I1(ram[4533]), .I2(ram[4525]), .I3(
        ram[4517]), .S0(n27231), .S1(n26756), .ZN(n24221) );
  MUX41 U12288 ( .I0(ram[4509]), .I1(ram[4501]), .I2(ram[4493]), .I3(
        ram[4485]), .S0(n27231), .S1(n26756), .ZN(n24223) );
  MUX41 U12289 ( .I0(ram[4605]), .I1(ram[4597]), .I2(ram[4589]), .I3(
        ram[4581]), .S0(n27231), .S1(n26756), .ZN(n24220) );
  MUX41 U12290 ( .I0(n24536), .I1(n24537), .I2(n24538), .I3(n24539), .S0(
        n26250), .S1(n26368), .ZN(n24535) );
  MUX41 U12291 ( .I0(ram[12221]), .I1(ram[12213]), .I2(ram[12205]), .I3(
        ram[12197]), .S0(n27250), .S1(n26775), .ZN(n24537) );
  MUX41 U12292 ( .I0(ram[12189]), .I1(ram[12181]), .I2(ram[12173]), .I3(
        ram[12165]), .S0(n27250), .S1(n26775), .ZN(n24539) );
  MUX41 U12293 ( .I0(ram[12285]), .I1(ram[12277]), .I2(ram[12269]), .I3(
        ram[12261]), .S0(n27250), .S1(n26775), .ZN(n24536) );
  MUX41 U12294 ( .I0(n24476), .I1(n24477), .I2(n24478), .I3(n24479), .S0(
        n26249), .S1(n26367), .ZN(n24475) );
  MUX41 U12295 ( .I0(ram[10685]), .I1(ram[10677]), .I2(ram[10669]), .I3(
        ram[10661]), .S0(n27246), .S1(n26771), .ZN(n24477) );
  MUX41 U12296 ( .I0(ram[10653]), .I1(ram[10645]), .I2(ram[10637]), .I3(
        ram[10629]), .S0(n27246), .S1(n26771), .ZN(n24479) );
  MUX41 U12297 ( .I0(ram[10749]), .I1(ram[10741]), .I2(ram[10733]), .I3(
        ram[10725]), .S0(n27246), .S1(n26771), .ZN(n24476) );
  MUX41 U12298 ( .I0(n24496), .I1(n24497), .I2(n24498), .I3(n24499), .S0(
        n26250), .S1(n26368), .ZN(n24495) );
  MUX41 U12299 ( .I0(ram[11197]), .I1(ram[11189]), .I2(ram[11181]), .I3(
        ram[11173]), .S0(n27247), .S1(n26772), .ZN(n24497) );
  MUX41 U12300 ( .I0(ram[11165]), .I1(ram[11157]), .I2(ram[11149]), .I3(
        ram[11141]), .S0(n27247), .S1(n26772), .ZN(n24499) );
  MUX41 U12301 ( .I0(ram[11261]), .I1(ram[11253]), .I2(ram[11245]), .I3(
        ram[11237]), .S0(n27247), .S1(n26772), .ZN(n24496) );
  MUX41 U12302 ( .I0(n24451), .I1(n24452), .I2(n24453), .I3(n24454), .S0(
        n26249), .S1(n26367), .ZN(n24450) );
  MUX41 U12303 ( .I0(ram[10173]), .I1(ram[10165]), .I2(ram[10157]), .I3(
        ram[10149]), .S0(n27245), .S1(n26770), .ZN(n24452) );
  MUX41 U12304 ( .I0(ram[10141]), .I1(ram[10133]), .I2(ram[10125]), .I3(
        ram[10117]), .S0(n27245), .S1(n26770), .ZN(n24454) );
  MUX41 U12305 ( .I0(ram[10237]), .I1(ram[10229]), .I2(ram[10221]), .I3(
        ram[10213]), .S0(n27245), .S1(n26770), .ZN(n24451) );
  MUX41 U12306 ( .I0(n24391), .I1(n24392), .I2(n24393), .I3(n24394), .S0(
        n26248), .S1(n26366), .ZN(n24390) );
  MUX41 U12307 ( .I0(ram[8637]), .I1(ram[8629]), .I2(ram[8621]), .I3(
        ram[8613]), .S0(n27241), .S1(n26766), .ZN(n24392) );
  MUX41 U12308 ( .I0(ram[8605]), .I1(ram[8597]), .I2(ram[8589]), .I3(
        ram[8581]), .S0(n27241), .S1(n26766), .ZN(n24394) );
  MUX41 U12309 ( .I0(ram[8701]), .I1(ram[8693]), .I2(ram[8685]), .I3(
        ram[8677]), .S0(n27241), .S1(n26766), .ZN(n24391) );
  MUX41 U12310 ( .I0(n24411), .I1(n24412), .I2(n24413), .I3(n24414), .S0(
        n26248), .S1(n26366), .ZN(n24410) );
  MUX41 U12311 ( .I0(ram[9117]), .I1(ram[9109]), .I2(ram[9101]), .I3(
        ram[9093]), .S0(n27242), .S1(n26767), .ZN(n24414) );
  MUX41 U12312 ( .I0(ram[9149]), .I1(ram[9141]), .I2(ram[9133]), .I3(
        ram[9125]), .S0(n27242), .S1(n26767), .ZN(n24412) );
  MUX41 U12313 ( .I0(ram[9213]), .I1(ram[9205]), .I2(ram[9197]), .I3(
        ram[9189]), .S0(n27242), .S1(n26767), .ZN(n24411) );
  MUX41 U12314 ( .I0(n25391), .I1(n25392), .I2(n25393), .I3(n25394), .S0(
        n26263), .S1(n26381), .ZN(n25390) );
  MUX41 U12315 ( .I0(ram[16286]), .I1(ram[16278]), .I2(ram[16270]), .I3(
        ram[16262]), .S0(n27299), .S1(n26824), .ZN(n25394) );
  MUX41 U12316 ( .I0(ram[16318]), .I1(ram[16310]), .I2(ram[16302]), .I3(
        ram[16294]), .S0(n27299), .S1(n26824), .ZN(n25392) );
  MUX41 U12317 ( .I0(ram[16382]), .I1(ram[16374]), .I2(ram[16366]), .I3(
        ram[16358]), .S0(n27299), .S1(n26824), .ZN(n25391) );
  MUX41 U12318 ( .I0(n25351), .I1(n25352), .I2(n25353), .I3(n25354), .S0(
        n26262), .S1(n26380), .ZN(n25350) );
  MUX41 U12319 ( .I0(ram[15262]), .I1(ram[15254]), .I2(ram[15246]), .I3(
        ram[15238]), .S0(n27296), .S1(n26821), .ZN(n25354) );
  MUX41 U12320 ( .I0(ram[15294]), .I1(ram[15286]), .I2(ram[15278]), .I3(
        ram[15270]), .S0(n27296), .S1(n26821), .ZN(n25352) );
  MUX41 U12321 ( .I0(ram[15358]), .I1(ram[15350]), .I2(ram[15342]), .I3(
        ram[15334]), .S0(n27297), .S1(n26822), .ZN(n25351) );
  MUX41 U12322 ( .I0(n25331), .I1(n25332), .I2(n25333), .I3(n25334), .S0(
        n26262), .S1(n26380), .ZN(n25330) );
  MUX41 U12323 ( .I0(ram[14750]), .I1(ram[14742]), .I2(ram[14734]), .I3(
        ram[14726]), .S0(n27295), .S1(n26820), .ZN(n25334) );
  MUX41 U12324 ( .I0(ram[14782]), .I1(ram[14774]), .I2(ram[14766]), .I3(
        ram[14758]), .S0(n27295), .S1(n26820), .ZN(n25332) );
  MUX41 U12325 ( .I0(ram[14846]), .I1(ram[14838]), .I2(ram[14830]), .I3(
        ram[14822]), .S0(n27295), .S1(n26820), .ZN(n25331) );
  MUX41 U12326 ( .I0(n25306), .I1(n25307), .I2(n25308), .I3(n25309), .S0(
        n26261), .S1(n26379), .ZN(n25305) );
  MUX41 U12327 ( .I0(ram[14238]), .I1(ram[14230]), .I2(ram[14222]), .I3(
        ram[14214]), .S0(n27294), .S1(n26819), .ZN(n25309) );
  MUX41 U12328 ( .I0(ram[14270]), .I1(ram[14262]), .I2(ram[14254]), .I3(
        ram[14246]), .S0(n27294), .S1(n26819), .ZN(n25307) );
  MUX41 U12329 ( .I0(ram[14334]), .I1(ram[14326]), .I2(ram[14318]), .I3(
        ram[14310]), .S0(n27294), .S1(n26819), .ZN(n25306) );
  MUX41 U12330 ( .I0(n25266), .I1(n25267), .I2(n25268), .I3(n25269), .S0(
        n26261), .S1(n26379), .ZN(n25265) );
  MUX41 U12331 ( .I0(ram[13214]), .I1(ram[13206]), .I2(ram[13198]), .I3(
        ram[13190]), .S0(n27291), .S1(n26816), .ZN(n25269) );
  MUX41 U12332 ( .I0(ram[13246]), .I1(ram[13238]), .I2(ram[13230]), .I3(
        ram[13222]), .S0(n27292), .S1(n26817), .ZN(n25267) );
  MUX41 U12333 ( .I0(ram[13310]), .I1(ram[13302]), .I2(ram[13294]), .I3(
        ram[13286]), .S0(n27292), .S1(n26817), .ZN(n25266) );
  MUX41 U12334 ( .I0(n25246), .I1(n25247), .I2(n25248), .I3(n25249), .S0(
        n26260), .S1(n26378), .ZN(n25245) );
  MUX41 U12335 ( .I0(ram[12702]), .I1(ram[12694]), .I2(ram[12686]), .I3(
        ram[12678]), .S0(n27290), .S1(n26815), .ZN(n25249) );
  MUX41 U12336 ( .I0(ram[12734]), .I1(ram[12726]), .I2(ram[12718]), .I3(
        ram[12710]), .S0(n27290), .S1(n26815), .ZN(n25247) );
  MUX41 U12337 ( .I0(ram[12798]), .I1(ram[12790]), .I2(ram[12782]), .I3(
        ram[12774]), .S0(n27290), .S1(n26815), .ZN(n25246) );
  MUX41 U12338 ( .I0(n25049), .I1(n25050), .I2(n25051), .I3(n25052), .S0(
        n26258), .S1(n26376), .ZN(n25048) );
  MUX41 U12339 ( .I0(ram[8126]), .I1(ram[8118]), .I2(ram[8110]), .I3(
        ram[8102]), .S0(n27279), .S1(n26804), .ZN(n25050) );
  MUX41 U12340 ( .I0(ram[8094]), .I1(ram[8086]), .I2(ram[8078]), .I3(
        ram[8070]), .S0(n27279), .S1(n26804), .ZN(n25052) );
  MUX41 U12341 ( .I0(ram[8190]), .I1(ram[8182]), .I2(ram[8174]), .I3(
        ram[8166]), .S0(n27279), .S1(n26804), .ZN(n25049) );
  MUX41 U12342 ( .I0(n24989), .I1(n24990), .I2(n24991), .I3(n24992), .S0(
        n26257), .S1(n26375), .ZN(n24988) );
  MUX41 U12343 ( .I0(ram[6558]), .I1(ram[6550]), .I2(ram[6542]), .I3(
        ram[6534]), .S0(n27275), .S1(n26800), .ZN(n24992) );
  MUX41 U12344 ( .I0(ram[6590]), .I1(ram[6582]), .I2(ram[6574]), .I3(
        ram[6566]), .S0(n27276), .S1(n26801), .ZN(n24990) );
  MUX41 U12345 ( .I0(ram[6654]), .I1(ram[6646]), .I2(ram[6638]), .I3(
        ram[6630]), .S0(n27276), .S1(n26801), .ZN(n24989) );
  MUX41 U12346 ( .I0(n25009), .I1(n25010), .I2(n25011), .I3(n25012), .S0(
        n26257), .S1(n26375), .ZN(n25008) );
  MUX41 U12347 ( .I0(ram[7070]), .I1(ram[7062]), .I2(ram[7054]), .I3(
        ram[7046]), .S0(n27277), .S1(n26802), .ZN(n25012) );
  MUX41 U12348 ( .I0(ram[7102]), .I1(ram[7094]), .I2(ram[7086]), .I3(
        ram[7078]), .S0(n27277), .S1(n26802), .ZN(n25010) );
  MUX41 U12349 ( .I0(ram[7166]), .I1(ram[7158]), .I2(ram[7150]), .I3(
        ram[7142]), .S0(n27277), .S1(n26802), .ZN(n25009) );
  MUX41 U12350 ( .I0(n24964), .I1(n24965), .I2(n24966), .I3(n24967), .S0(
        n26256), .S1(n26374), .ZN(n24963) );
  MUX41 U12351 ( .I0(ram[6078]), .I1(ram[6070]), .I2(ram[6062]), .I3(
        ram[6054]), .S0(n27274), .S1(n26799), .ZN(n24965) );
  MUX41 U12352 ( .I0(ram[6046]), .I1(ram[6038]), .I2(ram[6030]), .I3(
        ram[6022]), .S0(n27274), .S1(n26799), .ZN(n24967) );
  MUX41 U12353 ( .I0(ram[6142]), .I1(ram[6134]), .I2(ram[6126]), .I3(
        ram[6118]), .S0(n27274), .S1(n26799), .ZN(n24964) );
  MUX41 U12354 ( .I0(n24904), .I1(n24905), .I2(n24906), .I3(n24907), .S0(
        n26256), .S1(n26374), .ZN(n24903) );
  MUX41 U12355 ( .I0(ram[4542]), .I1(ram[4534]), .I2(ram[4526]), .I3(
        ram[4518]), .S0(n27271), .S1(n26796), .ZN(n24905) );
  MUX41 U12356 ( .I0(ram[4510]), .I1(ram[4502]), .I2(ram[4494]), .I3(
        ram[4486]), .S0(n27271), .S1(n26796), .ZN(n24907) );
  MUX41 U12357 ( .I0(ram[4606]), .I1(ram[4598]), .I2(ram[4590]), .I3(
        ram[4582]), .S0(n27271), .S1(n26796), .ZN(n24904) );
  MUX41 U12358 ( .I0(n25220), .I1(n25221), .I2(n25222), .I3(n25223), .S0(
        n26260), .S1(n26378), .ZN(n25219) );
  MUX41 U12359 ( .I0(ram[12222]), .I1(ram[12214]), .I2(ram[12206]), .I3(
        ram[12198]), .S0(n27289), .S1(n26814), .ZN(n25221) );
  MUX41 U12360 ( .I0(ram[12190]), .I1(ram[12182]), .I2(ram[12174]), .I3(
        ram[12166]), .S0(n27289), .S1(n26814), .ZN(n25223) );
  MUX41 U12361 ( .I0(ram[12286]), .I1(ram[12278]), .I2(ram[12270]), .I3(
        ram[12262]), .S0(n27289), .S1(n26814), .ZN(n25220) );
  MUX41 U12362 ( .I0(n25160), .I1(n25161), .I2(n25162), .I3(n25163), .S0(
        n26259), .S1(n26377), .ZN(n25159) );
  MUX41 U12363 ( .I0(ram[10686]), .I1(ram[10678]), .I2(ram[10670]), .I3(
        ram[10662]), .S0(n27285), .S1(n26810), .ZN(n25161) );
  MUX41 U12364 ( .I0(ram[10654]), .I1(ram[10646]), .I2(ram[10638]), .I3(
        ram[10630]), .S0(n27285), .S1(n26810), .ZN(n25163) );
  MUX41 U12365 ( .I0(ram[10750]), .I1(ram[10742]), .I2(ram[10734]), .I3(
        ram[10726]), .S0(n27286), .S1(n26811), .ZN(n25160) );
  MUX41 U12366 ( .I0(n25180), .I1(n25181), .I2(n25182), .I3(n25183), .S0(
        n26260), .S1(n26378), .ZN(n25179) );
  MUX41 U12367 ( .I0(ram[11198]), .I1(ram[11190]), .I2(ram[11182]), .I3(
        ram[11174]), .S0(n27287), .S1(n26812), .ZN(n25181) );
  MUX41 U12368 ( .I0(ram[11166]), .I1(ram[11158]), .I2(ram[11150]), .I3(
        ram[11142]), .S0(n27287), .S1(n26812), .ZN(n25183) );
  MUX41 U12369 ( .I0(ram[11262]), .I1(ram[11254]), .I2(ram[11246]), .I3(
        ram[11238]), .S0(n27287), .S1(n26812), .ZN(n25180) );
  MUX41 U12370 ( .I0(n25135), .I1(n25136), .I2(n25137), .I3(n25138), .S0(
        n26259), .S1(n26377), .ZN(n25134) );
  MUX41 U12371 ( .I0(ram[10174]), .I1(ram[10166]), .I2(ram[10158]), .I3(
        ram[10150]), .S0(n27284), .S1(n26809), .ZN(n25136) );
  MUX41 U12372 ( .I0(ram[10142]), .I1(ram[10134]), .I2(ram[10126]), .I3(
        ram[10118]), .S0(n27284), .S1(n26809), .ZN(n25138) );
  MUX41 U12373 ( .I0(ram[10238]), .I1(ram[10230]), .I2(ram[10222]), .I3(
        ram[10214]), .S0(n27284), .S1(n26809), .ZN(n25135) );
  MUX41 U12374 ( .I0(n25075), .I1(n25076), .I2(n25077), .I3(n25078), .S0(
        n26258), .S1(n26376), .ZN(n25074) );
  MUX41 U12375 ( .I0(ram[8638]), .I1(ram[8630]), .I2(ram[8622]), .I3(
        ram[8614]), .S0(n27280), .S1(n26805), .ZN(n25076) );
  MUX41 U12376 ( .I0(ram[8606]), .I1(ram[8598]), .I2(ram[8590]), .I3(
        ram[8582]), .S0(n27280), .S1(n26805), .ZN(n25078) );
  MUX41 U12377 ( .I0(ram[8702]), .I1(ram[8694]), .I2(ram[8686]), .I3(
        ram[8678]), .S0(n27281), .S1(n26806), .ZN(n25075) );
  MUX41 U12378 ( .I0(n25095), .I1(n25096), .I2(n25097), .I3(n25098), .S0(
        n26258), .S1(n26376), .ZN(n25094) );
  MUX41 U12379 ( .I0(ram[9118]), .I1(ram[9110]), .I2(ram[9102]), .I3(
        ram[9094]), .S0(n27282), .S1(n26807), .ZN(n25098) );
  MUX41 U12380 ( .I0(ram[9150]), .I1(ram[9142]), .I2(ram[9134]), .I3(
        ram[9126]), .S0(n27282), .S1(n26807), .ZN(n25096) );
  MUX41 U12381 ( .I0(ram[9214]), .I1(ram[9206]), .I2(ram[9198]), .I3(
        ram[9190]), .S0(n27282), .S1(n26807), .ZN(n25095) );
  MUX41 U12382 ( .I0(n26075), .I1(n26076), .I2(n26077), .I3(n26078), .S0(
        n26272), .S1(n26390), .ZN(n26074) );
  MUX41 U12383 ( .I0(ram[16287]), .I1(ram[16279]), .I2(ram[16271]), .I3(
        ram[16263]), .S0(n27338), .S1(n26863), .ZN(n26078) );
  MUX41 U12384 ( .I0(ram[16319]), .I1(ram[16311]), .I2(ram[16303]), .I3(
        ram[16295]), .S0(n27338), .S1(n26863), .ZN(n26076) );
  MUX41 U12385 ( .I0(ram[16383]), .I1(ram[16375]), .I2(ram[16367]), .I3(
        ram[16359]), .S0(n27338), .S1(n26863), .ZN(n26075) );
  MUX41 U12386 ( .I0(n26035), .I1(n26036), .I2(n26037), .I3(n26038), .S0(
        n26272), .S1(n26390), .ZN(n26034) );
  MUX41 U12387 ( .I0(ram[15263]), .I1(ram[15255]), .I2(ram[15247]), .I3(
        ram[15239]), .S0(n27336), .S1(n26861), .ZN(n26038) );
  MUX41 U12388 ( .I0(ram[15295]), .I1(ram[15287]), .I2(ram[15279]), .I3(
        ram[15271]), .S0(n27336), .S1(n26861), .ZN(n26036) );
  MUX41 U12389 ( .I0(ram[15359]), .I1(ram[15351]), .I2(ram[15343]), .I3(
        ram[15335]), .S0(n27336), .S1(n26861), .ZN(n26035) );
  MUX41 U12390 ( .I0(n26015), .I1(n26016), .I2(n26017), .I3(n26018), .S0(
        n26272), .S1(n26390), .ZN(n26014) );
  MUX41 U12391 ( .I0(ram[14751]), .I1(ram[14743]), .I2(ram[14735]), .I3(
        ram[14727]), .S0(n27335), .S1(n26860), .ZN(n26018) );
  MUX41 U12392 ( .I0(ram[14783]), .I1(ram[14775]), .I2(ram[14767]), .I3(
        ram[14759]), .S0(n27335), .S1(n26860), .ZN(n26016) );
  MUX41 U12393 ( .I0(ram[14847]), .I1(ram[14839]), .I2(ram[14831]), .I3(
        ram[14823]), .S0(n27335), .S1(n26860), .ZN(n26015) );
  MUX41 U12394 ( .I0(n25990), .I1(n25991), .I2(n25992), .I3(n25993), .S0(
        n26271), .S1(n26389), .ZN(n25989) );
  MUX41 U12395 ( .I0(ram[14239]), .I1(ram[14231]), .I2(ram[14223]), .I3(
        ram[14215]), .S0(n27333), .S1(n26858), .ZN(n25993) );
  MUX41 U12396 ( .I0(ram[14271]), .I1(ram[14263]), .I2(ram[14255]), .I3(
        ram[14247]), .S0(n27333), .S1(n26858), .ZN(n25991) );
  MUX41 U12397 ( .I0(ram[14335]), .I1(ram[14327]), .I2(ram[14319]), .I3(
        ram[14311]), .S0(n27334), .S1(n26859), .ZN(n25990) );
  MUX41 U12398 ( .I0(n25950), .I1(n25951), .I2(n25952), .I3(n25953), .S0(
        n26271), .S1(n26389), .ZN(n25949) );
  MUX41 U12399 ( .I0(ram[13215]), .I1(ram[13207]), .I2(ram[13199]), .I3(
        ram[13191]), .S0(n27331), .S1(n26856), .ZN(n25953) );
  MUX41 U12400 ( .I0(ram[13247]), .I1(ram[13239]), .I2(ram[13231]), .I3(
        ram[13223]), .S0(n27331), .S1(n26856), .ZN(n25951) );
  MUX41 U12401 ( .I0(ram[13311]), .I1(ram[13303]), .I2(ram[13295]), .I3(
        ram[13287]), .S0(n27331), .S1(n26856), .ZN(n25950) );
  MUX41 U12402 ( .I0(n25930), .I1(n25931), .I2(n25932), .I3(n25933), .S0(
        n26270), .S1(n26388), .ZN(n25929) );
  MUX41 U12403 ( .I0(ram[12703]), .I1(ram[12695]), .I2(ram[12687]), .I3(
        ram[12679]), .S0(n27330), .S1(n26855), .ZN(n25933) );
  MUX41 U12404 ( .I0(ram[12735]), .I1(ram[12727]), .I2(ram[12719]), .I3(
        ram[12711]), .S0(n27330), .S1(n26855), .ZN(n25931) );
  MUX41 U12405 ( .I0(ram[12799]), .I1(ram[12791]), .I2(ram[12783]), .I3(
        ram[12775]), .S0(n27330), .S1(n26855), .ZN(n25930) );
  MUX41 U12406 ( .I0(n25733), .I1(n25734), .I2(n25735), .I3(n25736), .S0(
        n26268), .S1(n26386), .ZN(n25732) );
  MUX41 U12407 ( .I0(ram[8127]), .I1(ram[8119]), .I2(ram[8111]), .I3(
        ram[8103]), .S0(n27319), .S1(n26844), .ZN(n25734) );
  MUX41 U12408 ( .I0(ram[8095]), .I1(ram[8087]), .I2(ram[8079]), .I3(
        ram[8071]), .S0(n27319), .S1(n26844), .ZN(n25736) );
  MUX41 U12409 ( .I0(ram[8191]), .I1(ram[8183]), .I2(ram[8175]), .I3(
        ram[8167]), .S0(n27319), .S1(n26844), .ZN(n25733) );
  MUX41 U12410 ( .I0(n25673), .I1(n25674), .I2(n25675), .I3(n25676), .S0(
        n26267), .S1(n26385), .ZN(n25672) );
  MUX41 U12411 ( .I0(ram[6559]), .I1(ram[6551]), .I2(ram[6543]), .I3(
        ram[6535]), .S0(n27315), .S1(n26840), .ZN(n25676) );
  MUX41 U12412 ( .I0(ram[6591]), .I1(ram[6583]), .I2(ram[6575]), .I3(
        ram[6567]), .S0(n27315), .S1(n26840), .ZN(n25674) );
  MUX41 U12413 ( .I0(ram[6655]), .I1(ram[6647]), .I2(ram[6639]), .I3(
        ram[6631]), .S0(n27315), .S1(n26840), .ZN(n25673) );
  MUX41 U12414 ( .I0(n25693), .I1(n25694), .I2(n25695), .I3(n25696), .S0(
        n26267), .S1(n26385), .ZN(n25692) );
  MUX41 U12415 ( .I0(ram[7071]), .I1(ram[7063]), .I2(ram[7055]), .I3(
        ram[7047]), .S0(n27316), .S1(n26841), .ZN(n25696) );
  MUX41 U12416 ( .I0(ram[7103]), .I1(ram[7095]), .I2(ram[7087]), .I3(
        ram[7079]), .S0(n27316), .S1(n26841), .ZN(n25694) );
  MUX41 U12417 ( .I0(ram[7167]), .I1(ram[7159]), .I2(ram[7151]), .I3(
        ram[7143]), .S0(n27316), .S1(n26841), .ZN(n25693) );
  MUX41 U12418 ( .I0(n25648), .I1(n25649), .I2(n25650), .I3(n25651), .S0(
        n26266), .S1(n26384), .ZN(n25647) );
  MUX41 U12419 ( .I0(ram[6079]), .I1(ram[6071]), .I2(ram[6063]), .I3(
        ram[6055]), .S0(n27314), .S1(n26839), .ZN(n25649) );
  MUX41 U12420 ( .I0(ram[6047]), .I1(ram[6039]), .I2(ram[6031]), .I3(
        ram[6023]), .S0(n27314), .S1(n26839), .ZN(n25651) );
  MUX41 U12421 ( .I0(ram[6143]), .I1(ram[6135]), .I2(ram[6127]), .I3(
        ram[6119]), .S0(n27314), .S1(n26839), .ZN(n25648) );
  MUX41 U12422 ( .I0(n25588), .I1(n25589), .I2(n25590), .I3(n25591), .S0(
        n26265), .S1(n26383), .ZN(n25587) );
  MUX41 U12423 ( .I0(ram[4543]), .I1(ram[4535]), .I2(ram[4527]), .I3(
        ram[4519]), .S0(n27310), .S1(n26835), .ZN(n25589) );
  MUX41 U12424 ( .I0(ram[4511]), .I1(ram[4503]), .I2(ram[4495]), .I3(
        ram[4487]), .S0(n27310), .S1(n26835), .ZN(n25591) );
  MUX41 U12425 ( .I0(ram[4607]), .I1(ram[4599]), .I2(ram[4591]), .I3(
        ram[4583]), .S0(n27310), .S1(n26835), .ZN(n25588) );
  MUX41 U12426 ( .I0(n25904), .I1(n25905), .I2(n25906), .I3(n25907), .S0(
        n26270), .S1(n26388), .ZN(n25903) );
  MUX41 U12427 ( .I0(ram[12223]), .I1(ram[12215]), .I2(ram[12207]), .I3(
        ram[12199]), .S0(n27328), .S1(n26853), .ZN(n25905) );
  MUX41 U12428 ( .I0(ram[12191]), .I1(ram[12183]), .I2(ram[12175]), .I3(
        ram[12167]), .S0(n27328), .S1(n26853), .ZN(n25907) );
  MUX41 U12429 ( .I0(ram[12287]), .I1(ram[12279]), .I2(ram[12271]), .I3(
        ram[12263]), .S0(n27329), .S1(n26854), .ZN(n25904) );
  MUX41 U12430 ( .I0(n25844), .I1(n25845), .I2(n25846), .I3(n25847), .S0(
        n26269), .S1(n26387), .ZN(n25843) );
  MUX41 U12431 ( .I0(ram[10687]), .I1(ram[10679]), .I2(ram[10671]), .I3(
        ram[10663]), .S0(n27325), .S1(n26850), .ZN(n25845) );
  MUX41 U12432 ( .I0(ram[10655]), .I1(ram[10647]), .I2(ram[10639]), .I3(
        ram[10631]), .S0(n27325), .S1(n26850), .ZN(n25847) );
  MUX41 U12433 ( .I0(ram[10751]), .I1(ram[10743]), .I2(ram[10735]), .I3(
        ram[10727]), .S0(n27325), .S1(n26850), .ZN(n25844) );
  MUX41 U12434 ( .I0(n25864), .I1(n25865), .I2(n25866), .I3(n25867), .S0(
        n26269), .S1(n26387), .ZN(n25863) );
  MUX41 U12435 ( .I0(ram[11199]), .I1(ram[11191]), .I2(ram[11183]), .I3(
        ram[11175]), .S0(n27326), .S1(n26851), .ZN(n25865) );
  MUX41 U12436 ( .I0(ram[11167]), .I1(ram[11159]), .I2(ram[11151]), .I3(
        ram[11143]), .S0(n27326), .S1(n26851), .ZN(n25867) );
  MUX41 U12437 ( .I0(ram[11263]), .I1(ram[11255]), .I2(ram[11247]), .I3(
        ram[11239]), .S0(n27326), .S1(n26851), .ZN(n25864) );
  MUX41 U12438 ( .I0(n25819), .I1(n25820), .I2(n25821), .I3(n25822), .S0(
        n26269), .S1(n26387), .ZN(n25818) );
  MUX41 U12439 ( .I0(ram[10175]), .I1(ram[10167]), .I2(ram[10159]), .I3(
        ram[10151]), .S0(n27324), .S1(n26849), .ZN(n25820) );
  MUX41 U12440 ( .I0(ram[10143]), .I1(ram[10135]), .I2(ram[10127]), .I3(
        ram[10119]), .S0(n27323), .S1(n26848), .ZN(n25822) );
  MUX41 U12441 ( .I0(ram[10239]), .I1(ram[10231]), .I2(ram[10223]), .I3(
        ram[10215]), .S0(n27324), .S1(n26849), .ZN(n25819) );
  MUX41 U12442 ( .I0(n25759), .I1(n25760), .I2(n25761), .I3(n25762), .S0(
        n26268), .S1(n26386), .ZN(n25758) );
  MUX41 U12443 ( .I0(ram[8639]), .I1(ram[8631]), .I2(ram[8623]), .I3(
        ram[8615]), .S0(n27320), .S1(n26845), .ZN(n25760) );
  MUX41 U12444 ( .I0(ram[8607]), .I1(ram[8599]), .I2(ram[8591]), .I3(
        ram[8583]), .S0(n27320), .S1(n26845), .ZN(n25762) );
  MUX41 U12445 ( .I0(ram[8703]), .I1(ram[8695]), .I2(ram[8687]), .I3(
        ram[8679]), .S0(n27320), .S1(n26845), .ZN(n25759) );
  MUX41 U12446 ( .I0(n25779), .I1(n25780), .I2(n25781), .I3(n25782), .S0(
        n26268), .S1(n26386), .ZN(n25778) );
  MUX41 U12447 ( .I0(ram[9119]), .I1(ram[9111]), .I2(ram[9103]), .I3(
        ram[9095]), .S0(n27321), .S1(n26846), .ZN(n25782) );
  MUX41 U12448 ( .I0(ram[9151]), .I1(ram[9143]), .I2(ram[9135]), .I3(
        ram[9127]), .S0(n27321), .S1(n26846), .ZN(n25780) );
  MUX41 U12449 ( .I0(ram[9215]), .I1(ram[9207]), .I2(ram[9199]), .I3(
        ram[9191]), .S0(n27321), .S1(n26846), .ZN(n25779) );
  MUX41 U12450 ( .I0(n20634), .I1(n20635), .I2(n20636), .I3(n20637), .S0(
        n26194), .S1(n26312), .ZN(n20633) );
  MUX41 U12451 ( .I0(ram[536]), .I1(ram[528]), .I2(ram[520]), .I3(
        ram[512]), .S0(n27025), .S1(n26550), .ZN(n20637) );
  MUX41 U12452 ( .I0(ram[568]), .I1(ram[560]), .I2(ram[552]), .I3(
        ram[544]), .S0(n27025), .S1(n26550), .ZN(n20635) );
  MUX41 U12453 ( .I0(ram[632]), .I1(ram[624]), .I2(ram[616]), .I3(
        ram[608]), .S0(n27025), .S1(n26550), .ZN(n20634) );
  MUX41 U12454 ( .I0(ram[3736]), .I1(ram[3728]), .I2(ram[3720]), .I3(
        ram[3712]), .S0(n27032), .S1(n26557), .ZN(n20767) );
  MUX41 U12455 ( .I0(ram[3608]), .I1(ram[3600]), .I2(ram[3592]), .I3(
        ram[3584]), .S0(n27032), .S1(n26557), .ZN(n20762) );
  MUX41 U12456 ( .I0(ram[2456]), .I1(ram[2448]), .I2(ram[2440]), .I3(
        ram[2432]), .S0(n27029), .S1(n26554), .ZN(n20717) );
  MUX41 U12457 ( .I0(ram[2200]), .I1(ram[2192]), .I2(ram[2184]), .I3(
        ram[2176]), .S0(n27029), .S1(n26554), .ZN(n20707) );
  MUX41 U12458 ( .I0(ram[2072]), .I1(ram[2064]), .I2(ram[2056]), .I3(
        ram[2048]), .S0(n27028), .S1(n26553), .ZN(n20702) );
  MUX41 U12459 ( .I0(ram[2968]), .I1(ram[2960]), .I2(ram[2952]), .I3(
        ram[2944]), .S0(n27031), .S1(n26556), .ZN(n20737) );
  MUX41 U12460 ( .I0(ram[2712]), .I1(ram[2704]), .I2(ram[2696]), .I3(
        ram[2688]), .S0(n27030), .S1(n26555), .ZN(n20727) );
  MUX41 U12461 ( .I0(ram[2584]), .I1(ram[2576]), .I2(ram[2568]), .I3(
        ram[2560]), .S0(n27030), .S1(n26555), .ZN(n20722) );
  MUX41 U12462 ( .I0(ram[1688]), .I1(ram[1680]), .I2(ram[1672]), .I3(
        ram[1664]), .S0(n27027), .S1(n26552), .ZN(n20682) );
  MUX41 U12463 ( .I0(ram[1560]), .I1(ram[1552]), .I2(ram[1544]), .I3(
        ram[1536]), .S0(n27027), .S1(n26552), .ZN(n20677) );
  MUX41 U12464 ( .I0(ram[408]), .I1(ram[400]), .I2(ram[392]), .I3(
        ram[384]), .S0(n27024), .S1(n26549), .ZN(n20632) );
  MUX41 U12465 ( .I0(ram[152]), .I1(ram[144]), .I2(ram[136]), .I3(
        ram[128]), .S0(n27024), .S1(n26549), .ZN(n3840) );
  MUX41 U12466 ( .I0(ram[3737]), .I1(ram[3729]), .I2(ram[3721]), .I3(
        ram[3713]), .S0(n27072), .S1(n26597), .ZN(n21451) );
  MUX41 U12467 ( .I0(ram[3609]), .I1(ram[3601]), .I2(ram[3593]), .I3(
        ram[3585]), .S0(n27071), .S1(n26596), .ZN(n21446) );
  MUX41 U12468 ( .I0(ram[2457]), .I1(ram[2449]), .I2(ram[2441]), .I3(
        ram[2433]), .S0(n27069), .S1(n26594), .ZN(n21401) );
  MUX41 U12469 ( .I0(ram[2201]), .I1(ram[2193]), .I2(ram[2185]), .I3(
        ram[2177]), .S0(n27068), .S1(n26593), .ZN(n21391) );
  MUX41 U12470 ( .I0(ram[2073]), .I1(ram[2065]), .I2(ram[2057]), .I3(
        ram[2049]), .S0(n27068), .S1(n26593), .ZN(n21386) );
  MUX41 U12471 ( .I0(ram[2969]), .I1(ram[2961]), .I2(ram[2953]), .I3(
        ram[2945]), .S0(n27070), .S1(n26595), .ZN(n21421) );
  MUX41 U12472 ( .I0(ram[2713]), .I1(ram[2705]), .I2(ram[2697]), .I3(
        ram[2689]), .S0(n27069), .S1(n26594), .ZN(n21411) );
  MUX41 U12473 ( .I0(ram[2585]), .I1(ram[2577]), .I2(ram[2569]), .I3(
        ram[2561]), .S0(n27069), .S1(n26594), .ZN(n21406) );
  MUX41 U12474 ( .I0(ram[1689]), .I1(ram[1681]), .I2(ram[1673]), .I3(
        ram[1665]), .S0(n27067), .S1(n26592), .ZN(n21366) );
  MUX41 U12475 ( .I0(ram[1561]), .I1(ram[1553]), .I2(ram[1545]), .I3(
        ram[1537]), .S0(n27067), .S1(n26592), .ZN(n21361) );
  MUX41 U12476 ( .I0(ram[409]), .I1(ram[401]), .I2(ram[393]), .I3(
        ram[385]), .S0(n27064), .S1(n26589), .ZN(n21316) );
  MUX41 U12477 ( .I0(ram[153]), .I1(ram[145]), .I2(ram[137]), .I3(
        ram[129]), .S0(n27063), .S1(n26588), .ZN(n21306) );
  MUX41 U12478 ( .I0(ram[25]), .I1(ram[17]), .I2(ram[9]), .I3(ram[1]), 
        .S0(n27063), .S1(n26588), .ZN(n21301) );
  MUX41 U12479 ( .I0(ram[3738]), .I1(ram[3730]), .I2(ram[3722]), .I3(
        ram[3714]), .S0(n27111), .S1(n26636), .ZN(n22135) );
  MUX41 U12480 ( .I0(ram[3610]), .I1(ram[3602]), .I2(ram[3594]), .I3(
        ram[3586]), .S0(n27111), .S1(n26636), .ZN(n22130) );
  MUX41 U12481 ( .I0(ram[2458]), .I1(ram[2450]), .I2(ram[2442]), .I3(
        ram[2434]), .S0(n27108), .S1(n26633), .ZN(n22085) );
  MUX41 U12482 ( .I0(ram[2202]), .I1(ram[2194]), .I2(ram[2186]), .I3(
        ram[2178]), .S0(n27107), .S1(n26632), .ZN(n22075) );
  MUX41 U12483 ( .I0(ram[2074]), .I1(ram[2066]), .I2(ram[2058]), .I3(
        ram[2050]), .S0(n27107), .S1(n26632), .ZN(n22070) );
  MUX41 U12484 ( .I0(ram[2970]), .I1(ram[2962]), .I2(ram[2954]), .I3(
        ram[2946]), .S0(n27109), .S1(n26634), .ZN(n22105) );
  MUX41 U12485 ( .I0(ram[2714]), .I1(ram[2706]), .I2(ram[2698]), .I3(
        ram[2690]), .S0(n27109), .S1(n26634), .ZN(n22095) );
  MUX41 U12486 ( .I0(ram[2586]), .I1(ram[2578]), .I2(ram[2570]), .I3(
        ram[2562]), .S0(n27108), .S1(n26633), .ZN(n22090) );
  MUX41 U12487 ( .I0(ram[1690]), .I1(ram[1682]), .I2(ram[1674]), .I3(
        ram[1666]), .S0(n27106), .S1(n26631), .ZN(n22050) );
  MUX41 U12488 ( .I0(ram[1562]), .I1(ram[1554]), .I2(ram[1546]), .I3(
        ram[1538]), .S0(n27106), .S1(n26631), .ZN(n22045) );
  MUX41 U12489 ( .I0(ram[410]), .I1(ram[402]), .I2(ram[394]), .I3(
        ram[386]), .S0(n27103), .S1(n26628), .ZN(n22000) );
  MUX41 U12490 ( .I0(ram[154]), .I1(ram[146]), .I2(ram[138]), .I3(
        ram[130]), .S0(n27103), .S1(n26628), .ZN(n21990) );
  MUX41 U12491 ( .I0(ram[26]), .I1(ram[18]), .I2(ram[10]), .I3(ram[2]), 
        .S0(n27102), .S1(n26627), .ZN(n21985) );
  MUX41 U12492 ( .I0(ram[3739]), .I1(ram[3731]), .I2(ram[3723]), .I3(
        ram[3715]), .S0(n27151), .S1(n26676), .ZN(n22819) );
  MUX41 U12493 ( .I0(ram[3611]), .I1(ram[3603]), .I2(ram[3595]), .I3(
        ram[3587]), .S0(n27150), .S1(n26675), .ZN(n22814) );
  MUX41 U12494 ( .I0(ram[2459]), .I1(ram[2451]), .I2(ram[2443]), .I3(
        ram[2435]), .S0(n27147), .S1(n26672), .ZN(n22769) );
  MUX41 U12495 ( .I0(ram[2203]), .I1(ram[2195]), .I2(ram[2187]), .I3(
        ram[2179]), .S0(n27147), .S1(n26672), .ZN(n22759) );
  MUX41 U12496 ( .I0(ram[2075]), .I1(ram[2067]), .I2(ram[2059]), .I3(
        ram[2051]), .S0(n27147), .S1(n26672), .ZN(n22754) );
  MUX41 U12497 ( .I0(ram[2971]), .I1(ram[2963]), .I2(ram[2955]), .I3(
        ram[2947]), .S0(n27149), .S1(n26674), .ZN(n22789) );
  MUX41 U12498 ( .I0(ram[2715]), .I1(ram[2707]), .I2(ram[2699]), .I3(
        ram[2691]), .S0(n27148), .S1(n26673), .ZN(n22779) );
  MUX41 U12499 ( .I0(ram[2587]), .I1(ram[2579]), .I2(ram[2571]), .I3(
        ram[2563]), .S0(n27148), .S1(n26673), .ZN(n22774) );
  MUX41 U12500 ( .I0(ram[1691]), .I1(ram[1683]), .I2(ram[1675]), .I3(
        ram[1667]), .S0(n27146), .S1(n26671), .ZN(n22734) );
  MUX41 U12501 ( .I0(ram[1563]), .I1(ram[1555]), .I2(ram[1547]), .I3(
        ram[1539]), .S0(n27145), .S1(n26670), .ZN(n22729) );
  MUX41 U12502 ( .I0(ram[411]), .I1(ram[403]), .I2(ram[395]), .I3(
        ram[387]), .S0(n27143), .S1(n26668), .ZN(n22684) );
  MUX41 U12503 ( .I0(ram[155]), .I1(ram[147]), .I2(ram[139]), .I3(
        ram[131]), .S0(n27142), .S1(n26667), .ZN(n22674) );
  MUX41 U12504 ( .I0(ram[27]), .I1(ram[19]), .I2(ram[11]), .I3(ram[3]), 
        .S0(n27142), .S1(n26667), .ZN(n22669) );
  MUX41 U12505 ( .I0(ram[3740]), .I1(ram[3732]), .I2(ram[3724]), .I3(
        ram[3716]), .S0(n27190), .S1(n26715), .ZN(n23503) );
  MUX41 U12506 ( .I0(ram[3612]), .I1(ram[3604]), .I2(ram[3596]), .I3(
        ram[3588]), .S0(n27190), .S1(n26715), .ZN(n23498) );
  MUX41 U12507 ( .I0(ram[2460]), .I1(ram[2452]), .I2(ram[2444]), .I3(
        ram[2436]), .S0(n27187), .S1(n26712), .ZN(n23453) );
  MUX41 U12508 ( .I0(ram[2204]), .I1(ram[2196]), .I2(ram[2188]), .I3(
        ram[2180]), .S0(n27186), .S1(n26711), .ZN(n23443) );
  MUX41 U12509 ( .I0(ram[2076]), .I1(ram[2068]), .I2(ram[2060]), .I3(
        ram[2052]), .S0(n27186), .S1(n26711), .ZN(n23438) );
  MUX41 U12510 ( .I0(ram[2972]), .I1(ram[2964]), .I2(ram[2956]), .I3(
        ram[2948]), .S0(n27188), .S1(n26713), .ZN(n23473) );
  MUX41 U12511 ( .I0(ram[2716]), .I1(ram[2708]), .I2(ram[2700]), .I3(
        ram[2692]), .S0(n27187), .S1(n26712), .ZN(n23463) );
  MUX41 U12512 ( .I0(ram[2588]), .I1(ram[2580]), .I2(ram[2572]), .I3(
        ram[2564]), .S0(n27187), .S1(n26712), .ZN(n23458) );
  MUX41 U12513 ( .I0(ram[1692]), .I1(ram[1684]), .I2(ram[1676]), .I3(
        ram[1668]), .S0(n27185), .S1(n26710), .ZN(n23418) );
  MUX41 U12514 ( .I0(ram[1564]), .I1(ram[1556]), .I2(ram[1548]), .I3(
        ram[1540]), .S0(n27185), .S1(n26710), .ZN(n23413) );
  MUX41 U12515 ( .I0(ram[412]), .I1(ram[404]), .I2(ram[396]), .I3(
        ram[388]), .S0(n27182), .S1(n26707), .ZN(n23368) );
  MUX41 U12516 ( .I0(ram[156]), .I1(ram[148]), .I2(ram[140]), .I3(
        ram[132]), .S0(n27181), .S1(n26706), .ZN(n23358) );
  MUX41 U12517 ( .I0(ram[28]), .I1(ram[20]), .I2(ram[12]), .I3(ram[4]), 
        .S0(n27181), .S1(n26706), .ZN(n23353) );
  MUX41 U12518 ( .I0(ram[3741]), .I1(ram[3733]), .I2(ram[3725]), .I3(
        ram[3717]), .S0(n27229), .S1(n26754), .ZN(n24187) );
  MUX41 U12519 ( .I0(ram[3613]), .I1(ram[3605]), .I2(ram[3597]), .I3(
        ram[3589]), .S0(n27229), .S1(n26754), .ZN(n24182) );
  MUX41 U12520 ( .I0(ram[2461]), .I1(ram[2453]), .I2(ram[2445]), .I3(
        ram[2437]), .S0(n27226), .S1(n26751), .ZN(n24137) );
  MUX41 U12521 ( .I0(ram[2205]), .I1(ram[2197]), .I2(ram[2189]), .I3(
        ram[2181]), .S0(n27226), .S1(n26751), .ZN(n24127) );
  MUX41 U12522 ( .I0(ram[2077]), .I1(ram[2069]), .I2(ram[2061]), .I3(
        ram[2053]), .S0(n27225), .S1(n26750), .ZN(n24122) );
  MUX41 U12523 ( .I0(ram[2973]), .I1(ram[2965]), .I2(ram[2957]), .I3(
        ram[2949]), .S0(n27227), .S1(n26752), .ZN(n24157) );
  MUX41 U12524 ( .I0(ram[2717]), .I1(ram[2709]), .I2(ram[2701]), .I3(
        ram[2693]), .S0(n27227), .S1(n26752), .ZN(n24147) );
  MUX41 U12525 ( .I0(ram[2589]), .I1(ram[2581]), .I2(ram[2573]), .I3(
        ram[2565]), .S0(n27227), .S1(n26752), .ZN(n24142) );
  MUX41 U12526 ( .I0(ram[1693]), .I1(ram[1685]), .I2(ram[1677]), .I3(
        ram[1669]), .S0(n27224), .S1(n26749), .ZN(n24102) );
  MUX41 U12527 ( .I0(ram[1565]), .I1(ram[1557]), .I2(ram[1549]), .I3(
        ram[1541]), .S0(n27224), .S1(n26749), .ZN(n24097) );
  MUX41 U12528 ( .I0(ram[413]), .I1(ram[405]), .I2(ram[397]), .I3(
        ram[389]), .S0(n27221), .S1(n26746), .ZN(n24052) );
  MUX41 U12529 ( .I0(ram[157]), .I1(ram[149]), .I2(ram[141]), .I3(
        ram[133]), .S0(n27221), .S1(n26746), .ZN(n24042) );
  MUX41 U12530 ( .I0(ram[29]), .I1(ram[21]), .I2(ram[13]), .I3(ram[5]), 
        .S0(n27220), .S1(n26745), .ZN(n24037) );
  MUX41 U12531 ( .I0(ram[3742]), .I1(ram[3734]), .I2(ram[3726]), .I3(
        ram[3718]), .S0(n27269), .S1(n26794), .ZN(n24871) );
  MUX41 U12532 ( .I0(ram[3614]), .I1(ram[3606]), .I2(ram[3598]), .I3(
        ram[3590]), .S0(n27268), .S1(n26793), .ZN(n24866) );
  MUX41 U12533 ( .I0(ram[2462]), .I1(ram[2454]), .I2(ram[2446]), .I3(
        ram[2438]), .S0(n27266), .S1(n26791), .ZN(n24821) );
  MUX41 U12534 ( .I0(ram[2206]), .I1(ram[2198]), .I2(ram[2190]), .I3(
        ram[2182]), .S0(n27265), .S1(n26790), .ZN(n24811) );
  MUX41 U12535 ( .I0(ram[2078]), .I1(ram[2070]), .I2(ram[2062]), .I3(
        ram[2054]), .S0(n27265), .S1(n26790), .ZN(n24806) );
  MUX41 U12536 ( .I0(ram[2974]), .I1(ram[2966]), .I2(ram[2958]), .I3(
        ram[2950]), .S0(n27267), .S1(n26792), .ZN(n24841) );
  MUX41 U12537 ( .I0(ram[2718]), .I1(ram[2710]), .I2(ram[2702]), .I3(
        ram[2694]), .S0(n27266), .S1(n26791), .ZN(n24831) );
  MUX41 U12538 ( .I0(ram[2590]), .I1(ram[2582]), .I2(ram[2574]), .I3(
        ram[2566]), .S0(n27266), .S1(n26791), .ZN(n24826) );
  MUX41 U12539 ( .I0(ram[1694]), .I1(ram[1686]), .I2(ram[1678]), .I3(
        ram[1670]), .S0(n27264), .S1(n26789), .ZN(n24786) );
  MUX41 U12540 ( .I0(ram[1566]), .I1(ram[1558]), .I2(ram[1550]), .I3(
        ram[1542]), .S0(n27263), .S1(n26788), .ZN(n24781) );
  MUX41 U12541 ( .I0(ram[414]), .I1(ram[406]), .I2(ram[398]), .I3(
        ram[390]), .S0(n27261), .S1(n26786), .ZN(n24736) );
  MUX41 U12542 ( .I0(ram[158]), .I1(ram[150]), .I2(ram[142]), .I3(
        ram[134]), .S0(n27260), .S1(n26785), .ZN(n24726) );
  MUX41 U12543 ( .I0(ram[30]), .I1(ram[22]), .I2(ram[14]), .I3(ram[6]), 
        .S0(n27260), .S1(n26785), .ZN(n24721) );
  MUX41 U12544 ( .I0(ram[3743]), .I1(ram[3735]), .I2(ram[3727]), .I3(
        ram[3719]), .S0(n27308), .S1(n26833), .ZN(n25555) );
  MUX41 U12545 ( .I0(ram[3615]), .I1(ram[3607]), .I2(ram[3599]), .I3(
        ram[3591]), .S0(n27308), .S1(n26833), .ZN(n25550) );
  MUX41 U12546 ( .I0(ram[2463]), .I1(ram[2455]), .I2(ram[2447]), .I3(
        ram[2439]), .S0(n27305), .S1(n26830), .ZN(n25505) );
  MUX41 U12547 ( .I0(ram[2207]), .I1(ram[2199]), .I2(ram[2191]), .I3(
        ram[2183]), .S0(n27304), .S1(n26829), .ZN(n25495) );
  MUX41 U12548 ( .I0(ram[2079]), .I1(ram[2071]), .I2(ram[2063]), .I3(
        ram[2055]), .S0(n27304), .S1(n26829), .ZN(n25490) );
  MUX41 U12549 ( .I0(ram[2975]), .I1(ram[2967]), .I2(ram[2959]), .I3(
        ram[2951]), .S0(n27306), .S1(n26831), .ZN(n25525) );
  MUX41 U12550 ( .I0(ram[2719]), .I1(ram[2711]), .I2(ram[2703]), .I3(
        ram[2695]), .S0(n27306), .S1(n26831), .ZN(n25515) );
  MUX41 U12551 ( .I0(ram[2591]), .I1(ram[2583]), .I2(ram[2575]), .I3(
        ram[2567]), .S0(n27305), .S1(n26830), .ZN(n25510) );
  MUX41 U12552 ( .I0(ram[1695]), .I1(ram[1687]), .I2(ram[1679]), .I3(
        ram[1671]), .S0(n27303), .S1(n26828), .ZN(n25470) );
  MUX41 U12553 ( .I0(ram[1567]), .I1(ram[1559]), .I2(ram[1551]), .I3(
        ram[1543]), .S0(n27303), .S1(n26828), .ZN(n25465) );
  MUX41 U12554 ( .I0(ram[415]), .I1(ram[407]), .I2(ram[399]), .I3(
        ram[391]), .S0(n27300), .S1(n26825), .ZN(n25420) );
  MUX41 U12555 ( .I0(ram[159]), .I1(ram[151]), .I2(ram[143]), .I3(
        ram[135]), .S0(n27299), .S1(n26824), .ZN(n25410) );
  MUX41 U12556 ( .I0(ram[31]), .I1(ram[23]), .I2(ram[15]), .I3(ram[7]), 
        .S0(n27299), .S1(n26824), .ZN(n25405) );
  MUX41 U12557 ( .I0(ram[5272]), .I1(ram[5264]), .I2(ram[5256]), .I3(
        ram[5248]), .S0(n27036), .S1(n26561), .ZN(n20833) );
  MUX41 U12558 ( .I0(ram[5144]), .I1(ram[5136]), .I2(ram[5128]), .I3(
        ram[5120]), .S0(n27036), .S1(n26561), .ZN(n20828) );
  MUX41 U12559 ( .I0(ram[9240]), .I1(ram[9232]), .I2(ram[9224]), .I3(
        ram[9216]), .S0(n27046), .S1(n26571), .ZN(n20999) );
  MUX41 U12560 ( .I0(n21318), .I1(n21319), .I2(n21320), .I3(n21321), .S0(
        n26204), .S1(n26322), .ZN(n21317) );
  MUX41 U12561 ( .I0(ram[537]), .I1(ram[529]), .I2(ram[521]), .I3(
        ram[513]), .S0(n27064), .S1(n26589), .ZN(n21321) );
  MUX41 U12562 ( .I0(ram[569]), .I1(ram[561]), .I2(ram[553]), .I3(
        ram[545]), .S0(n27064), .S1(n26589), .ZN(n21319) );
  MUX41 U12563 ( .I0(ram[633]), .I1(ram[625]), .I2(ram[617]), .I3(
        ram[609]), .S0(n27064), .S1(n26589), .ZN(n21318) );
  MUX41 U12564 ( .I0(ram[5273]), .I1(ram[5265]), .I2(ram[5257]), .I3(
        ram[5249]), .S0(n27075), .S1(n26600), .ZN(n21517) );
  MUX41 U12565 ( .I0(ram[5145]), .I1(ram[5137]), .I2(ram[5129]), .I3(
        ram[5121]), .S0(n27075), .S1(n26600), .ZN(n21512) );
  MUX41 U12566 ( .I0(ram[9241]), .I1(ram[9233]), .I2(ram[9225]), .I3(
        ram[9217]), .S0(n27085), .S1(n26610), .ZN(n21683) );
  MUX41 U12567 ( .I0(ram[5274]), .I1(ram[5266]), .I2(ram[5258]), .I3(
        ram[5250]), .S0(n27115), .S1(n26640), .ZN(n22201) );
  MUX41 U12568 ( .I0(ram[5146]), .I1(ram[5138]), .I2(ram[5130]), .I3(
        ram[5122]), .S0(n27115), .S1(n26640), .ZN(n22196) );
  MUX41 U12569 ( .I0(ram[5275]), .I1(ram[5267]), .I2(ram[5259]), .I3(
        ram[5251]), .S0(n27154), .S1(n26679), .ZN(n22885) );
  MUX41 U12570 ( .I0(ram[5147]), .I1(ram[5139]), .I2(ram[5131]), .I3(
        ram[5123]), .S0(n27154), .S1(n26679), .ZN(n22880) );
  MUX41 U12571 ( .I0(ram[5276]), .I1(ram[5268]), .I2(ram[5260]), .I3(
        ram[5252]), .S0(n27194), .S1(n26719), .ZN(n23569) );
  MUX41 U12572 ( .I0(ram[5148]), .I1(ram[5140]), .I2(ram[5132]), .I3(
        ram[5124]), .S0(n27193), .S1(n26718), .ZN(n23564) );
  MUX41 U12573 ( .I0(ram[5277]), .I1(ram[5269]), .I2(ram[5261]), .I3(
        ram[5253]), .S0(n27233), .S1(n26758), .ZN(n24253) );
  MUX41 U12574 ( .I0(ram[5149]), .I1(ram[5141]), .I2(ram[5133]), .I3(
        ram[5125]), .S0(n27233), .S1(n26758), .ZN(n24248) );
  MUX41 U12575 ( .I0(ram[5278]), .I1(ram[5270]), .I2(ram[5262]), .I3(
        ram[5254]), .S0(n27272), .S1(n26797), .ZN(n24937) );
  MUX41 U12576 ( .I0(ram[5150]), .I1(ram[5142]), .I2(ram[5134]), .I3(
        ram[5126]), .S0(n27272), .S1(n26797), .ZN(n24932) );
  MUX41 U12577 ( .I0(ram[5279]), .I1(ram[5271]), .I2(ram[5263]), .I3(
        ram[5255]), .S0(n27312), .S1(n26837), .ZN(n25621) );
  MUX41 U12578 ( .I0(ram[5151]), .I1(ram[5143]), .I2(ram[5135]), .I3(
        ram[5127]), .S0(n27311), .S1(n26836), .ZN(n25616) );
  MUX41 U12579 ( .I0(n20890), .I1(n20891), .I2(n20892), .I3(n20893), .S0(
        n26198), .S1(n26316), .ZN(n20889) );
  MUX41 U12580 ( .I0(ram[6680]), .I1(ram[6672]), .I2(ram[6664]), .I3(
        ram[6656]), .S0(n27039), .S1(n26564), .ZN(n20893) );
  MUX41 U12581 ( .I0(ram[6712]), .I1(ram[6704]), .I2(ram[6696]), .I3(
        ram[6688]), .S0(n27040), .S1(n26565), .ZN(n20891) );
  MUX41 U12582 ( .I0(ram[6776]), .I1(ram[6768]), .I2(ram[6760]), .I3(
        ram[6752]), .S0(n27040), .S1(n26565), .ZN(n20890) );
  MUX41 U12583 ( .I0(n20785), .I1(n20786), .I2(n20787), .I3(n20788), .S0(
        n26196), .S1(n26314), .ZN(n20784) );
  MUX41 U12584 ( .I0(ram[4152]), .I1(ram[4144]), .I2(ram[4136]), .I3(
        ram[4128]), .S0(n27033), .S1(n26558), .ZN(n20786) );
  MUX41 U12585 ( .I0(ram[4120]), .I1(ram[4112]), .I2(ram[4104]), .I3(
        ram[4096]), .S0(n27033), .S1(n26558), .ZN(n20788) );
  MUX41 U12586 ( .I0(ram[4216]), .I1(ram[4208]), .I2(ram[4200]), .I3(
        ram[4192]), .S0(n27034), .S1(n26559), .ZN(n20785) );
  MUX41 U12587 ( .I0(n20805), .I1(n20806), .I2(n20807), .I3(n20808), .S0(
        n26197), .S1(n26315), .ZN(n20804) );
  MUX41 U12588 ( .I0(ram[4664]), .I1(ram[4656]), .I2(ram[4648]), .I3(
        ram[4640]), .S0(n27035), .S1(n26560), .ZN(n20806) );
  MUX41 U12589 ( .I0(ram[4632]), .I1(ram[4624]), .I2(ram[4616]), .I3(
        ram[4608]), .S0(n27035), .S1(n26560), .ZN(n20808) );
  MUX41 U12590 ( .I0(ram[4728]), .I1(ram[4720]), .I2(ram[4712]), .I3(
        ram[4704]), .S0(n27035), .S1(n26560), .ZN(n20805) );
  MUX41 U12591 ( .I0(n21061), .I1(n21062), .I2(n21063), .I3(n21064), .S0(
        n26200), .S1(n26318), .ZN(n21060) );
  MUX41 U12592 ( .I0(ram[10808]), .I1(ram[10800]), .I2(ram[10792]), .I3(
        ram[10784]), .S0(n27049), .S1(n26574), .ZN(n21062) );
  MUX41 U12593 ( .I0(ram[10776]), .I1(ram[10768]), .I2(ram[10760]), .I3(
        ram[10752]), .S0(n27049), .S1(n26574), .ZN(n21064) );
  MUX41 U12594 ( .I0(ram[10872]), .I1(ram[10864]), .I2(ram[10856]), .I3(
        ram[10848]), .S0(n27050), .S1(n26575), .ZN(n21061) );
  MUX41 U12595 ( .I0(n20956), .I1(n20957), .I2(n20958), .I3(n20959), .S0(
        n26199), .S1(n26317), .ZN(n20955) );
  MUX41 U12596 ( .I0(ram[8248]), .I1(ram[8240]), .I2(ram[8232]), .I3(
        ram[8224]), .S0(n27043), .S1(n26568), .ZN(n20957) );
  MUX41 U12597 ( .I0(ram[8216]), .I1(ram[8208]), .I2(ram[8200]), .I3(
        ram[8192]), .S0(n27043), .S1(n26568), .ZN(n20959) );
  MUX41 U12598 ( .I0(ram[8312]), .I1(ram[8304]), .I2(ram[8296]), .I3(
        ram[8288]), .S0(n27043), .S1(n26568), .ZN(n20956) );
  MUX41 U12599 ( .I0(n20976), .I1(n20977), .I2(n20978), .I3(n20979), .S0(
        n26199), .S1(n26317), .ZN(n20975) );
  MUX41 U12600 ( .I0(ram[8760]), .I1(ram[8752]), .I2(ram[8744]), .I3(
        ram[8736]), .S0(n27044), .S1(n26569), .ZN(n20977) );
  MUX41 U12601 ( .I0(ram[8728]), .I1(ram[8720]), .I2(ram[8712]), .I3(
        ram[8704]), .S0(n27044), .S1(n26569), .ZN(n20979) );
  MUX41 U12602 ( .I0(ram[8824]), .I1(ram[8816]), .I2(ram[8808]), .I3(
        ram[8800]), .S0(n27045), .S1(n26570), .ZN(n20976) );
  MUX41 U12603 ( .I0(n21574), .I1(n21575), .I2(n21576), .I3(n21577), .S0(
        n26208), .S1(n26326), .ZN(n21573) );
  MUX41 U12604 ( .I0(ram[6681]), .I1(ram[6673]), .I2(ram[6665]), .I3(
        ram[6657]), .S0(n27079), .S1(n26604), .ZN(n21577) );
  MUX41 U12605 ( .I0(ram[6713]), .I1(ram[6705]), .I2(ram[6697]), .I3(
        ram[6689]), .S0(n27079), .S1(n26604), .ZN(n21575) );
  MUX41 U12606 ( .I0(ram[6777]), .I1(ram[6769]), .I2(ram[6761]), .I3(
        ram[6753]), .S0(n27079), .S1(n26604), .ZN(n21574) );
  MUX41 U12607 ( .I0(n21469), .I1(n21470), .I2(n21471), .I3(n21472), .S0(
        n26206), .S1(n26324), .ZN(n21468) );
  MUX41 U12608 ( .I0(ram[4153]), .I1(ram[4145]), .I2(ram[4137]), .I3(
        ram[4129]), .S0(n27073), .S1(n26598), .ZN(n21470) );
  MUX41 U12609 ( .I0(ram[4121]), .I1(ram[4113]), .I2(ram[4105]), .I3(
        ram[4097]), .S0(n27073), .S1(n26598), .ZN(n21472) );
  MUX41 U12610 ( .I0(ram[4217]), .I1(ram[4209]), .I2(ram[4201]), .I3(
        ram[4193]), .S0(n27073), .S1(n26598), .ZN(n21469) );
  MUX41 U12611 ( .I0(n21489), .I1(n21490), .I2(n21491), .I3(n21492), .S0(
        n26206), .S1(n26324), .ZN(n21488) );
  MUX41 U12612 ( .I0(ram[4665]), .I1(ram[4657]), .I2(ram[4649]), .I3(
        ram[4641]), .S0(n27074), .S1(n26599), .ZN(n21490) );
  MUX41 U12613 ( .I0(ram[4633]), .I1(ram[4625]), .I2(ram[4617]), .I3(
        ram[4609]), .S0(n27074), .S1(n26599), .ZN(n21492) );
  MUX41 U12614 ( .I0(ram[4729]), .I1(ram[4721]), .I2(ram[4713]), .I3(
        ram[4705]), .S0(n27074), .S1(n26599), .ZN(n21489) );
  MUX41 U12615 ( .I0(n21745), .I1(n21746), .I2(n21747), .I3(n21748), .S0(
        n26210), .S1(n26328), .ZN(n21744) );
  MUX41 U12616 ( .I0(ram[10809]), .I1(ram[10801]), .I2(ram[10793]), .I3(
        ram[10785]), .S0(n27089), .S1(n26614), .ZN(n21746) );
  MUX41 U12617 ( .I0(ram[10777]), .I1(ram[10769]), .I2(ram[10761]), .I3(
        ram[10753]), .S0(n27089), .S1(n26614), .ZN(n21748) );
  MUX41 U12618 ( .I0(ram[10873]), .I1(ram[10865]), .I2(ram[10857]), .I3(
        ram[10849]), .S0(n27089), .S1(n26614), .ZN(n21745) );
  MUX41 U12619 ( .I0(n21640), .I1(n21641), .I2(n21642), .I3(n21643), .S0(
        n26209), .S1(n26327), .ZN(n21639) );
  MUX41 U12620 ( .I0(ram[8249]), .I1(ram[8241]), .I2(ram[8233]), .I3(
        ram[8225]), .S0(n27083), .S1(n26608), .ZN(n21641) );
  MUX41 U12621 ( .I0(ram[8217]), .I1(ram[8209]), .I2(ram[8201]), .I3(
        ram[8193]), .S0(n27083), .S1(n26608), .ZN(n21643) );
  MUX41 U12622 ( .I0(ram[8313]), .I1(ram[8305]), .I2(ram[8297]), .I3(
        ram[8289]), .S0(n27083), .S1(n26608), .ZN(n21640) );
  MUX41 U12623 ( .I0(n21660), .I1(n21661), .I2(n21662), .I3(n21663), .S0(
        n26209), .S1(n26327), .ZN(n21659) );
  MUX41 U12624 ( .I0(ram[8761]), .I1(ram[8753]), .I2(ram[8745]), .I3(
        ram[8737]), .S0(n27084), .S1(n26609), .ZN(n21661) );
  MUX41 U12625 ( .I0(ram[8729]), .I1(ram[8721]), .I2(ram[8713]), .I3(
        ram[8705]), .S0(n27084), .S1(n26609), .ZN(n21663) );
  MUX41 U12626 ( .I0(ram[8825]), .I1(ram[8817]), .I2(ram[8809]), .I3(
        ram[8801]), .S0(n27084), .S1(n26609), .ZN(n21660) );
  MUX41 U12627 ( .I0(n22153), .I1(n22154), .I2(n22155), .I3(n22156), .S0(
        n26216), .S1(n26334), .ZN(n22152) );
  MUX41 U12628 ( .I0(ram[4154]), .I1(ram[4146]), .I2(ram[4138]), .I3(
        ram[4130]), .S0(n27112), .S1(n26637), .ZN(n22154) );
  MUX41 U12629 ( .I0(ram[4122]), .I1(ram[4114]), .I2(ram[4106]), .I3(
        ram[4098]), .S0(n27112), .S1(n26637), .ZN(n22156) );
  MUX41 U12630 ( .I0(ram[4218]), .I1(ram[4210]), .I2(ram[4202]), .I3(
        ram[4194]), .S0(n27112), .S1(n26637), .ZN(n22153) );
  MUX41 U12631 ( .I0(n22173), .I1(n22174), .I2(n22175), .I3(n22176), .S0(
        n26216), .S1(n26334), .ZN(n22172) );
  MUX41 U12632 ( .I0(ram[4666]), .I1(ram[4658]), .I2(ram[4650]), .I3(
        ram[4642]), .S0(n27113), .S1(n26638), .ZN(n22174) );
  MUX41 U12633 ( .I0(ram[4634]), .I1(ram[4626]), .I2(ram[4618]), .I3(
        ram[4610]), .S0(n27113), .S1(n26638), .ZN(n22176) );
  MUX41 U12634 ( .I0(ram[4730]), .I1(ram[4722]), .I2(ram[4714]), .I3(
        ram[4706]), .S0(n27114), .S1(n26639), .ZN(n22173) );
  MUX41 U12635 ( .I0(n22429), .I1(n22430), .I2(n22431), .I3(n22432), .S0(
        n26220), .S1(n26338), .ZN(n22428) );
  MUX41 U12636 ( .I0(ram[10810]), .I1(ram[10802]), .I2(ram[10794]), .I3(
        ram[10786]), .S0(n27128), .S1(n26653), .ZN(n22430) );
  MUX41 U12637 ( .I0(ram[10778]), .I1(ram[10770]), .I2(ram[10762]), .I3(
        ram[10754]), .S0(n27128), .S1(n26653), .ZN(n22432) );
  MUX41 U12638 ( .I0(ram[10874]), .I1(ram[10866]), .I2(ram[10858]), .I3(
        ram[10850]), .S0(n27128), .S1(n26653), .ZN(n22429) );
  MUX41 U12639 ( .I0(n22344), .I1(n22345), .I2(n22346), .I3(n22347), .S0(
        n26219), .S1(n26337), .ZN(n22343) );
  MUX41 U12640 ( .I0(ram[8762]), .I1(ram[8754]), .I2(ram[8746]), .I3(
        ram[8738]), .S0(n27123), .S1(n26648), .ZN(n22345) );
  MUX41 U12641 ( .I0(ram[8730]), .I1(ram[8722]), .I2(ram[8714]), .I3(
        ram[8706]), .S0(n27123), .S1(n26648), .ZN(n22347) );
  MUX41 U12642 ( .I0(ram[8826]), .I1(ram[8818]), .I2(ram[8810]), .I3(
        ram[8802]), .S0(n27123), .S1(n26648), .ZN(n22344) );
  MUX41 U12643 ( .I0(n22837), .I1(n22838), .I2(n22839), .I3(n22840), .S0(
        n26226), .S1(n26344), .ZN(n22836) );
  MUX41 U12644 ( .I0(ram[4155]), .I1(ram[4147]), .I2(ram[4139]), .I3(
        ram[4131]), .S0(n27152), .S1(n26677), .ZN(n22838) );
  MUX41 U12645 ( .I0(ram[4123]), .I1(ram[4115]), .I2(ram[4107]), .I3(
        ram[4099]), .S0(n27151), .S1(n26676), .ZN(n22840) );
  MUX41 U12646 ( .I0(ram[4219]), .I1(ram[4211]), .I2(ram[4203]), .I3(
        ram[4195]), .S0(n27152), .S1(n26677), .ZN(n22837) );
  MUX41 U12647 ( .I0(n22857), .I1(n22858), .I2(n22859), .I3(n22860), .S0(
        n26226), .S1(n26344), .ZN(n22856) );
  MUX41 U12648 ( .I0(ram[4667]), .I1(ram[4659]), .I2(ram[4651]), .I3(
        ram[4643]), .S0(n27153), .S1(n26678), .ZN(n22858) );
  MUX41 U12649 ( .I0(ram[4635]), .I1(ram[4627]), .I2(ram[4619]), .I3(
        ram[4611]), .S0(n27153), .S1(n26678), .ZN(n22860) );
  MUX41 U12650 ( .I0(ram[4731]), .I1(ram[4723]), .I2(ram[4715]), .I3(
        ram[4707]), .S0(n27153), .S1(n26678), .ZN(n22857) );
  MUX41 U12651 ( .I0(n23113), .I1(n23114), .I2(n23115), .I3(n23116), .S0(
        n26230), .S1(n26348), .ZN(n23112) );
  MUX41 U12652 ( .I0(ram[10811]), .I1(ram[10803]), .I2(ram[10795]), .I3(
        ram[10787]), .S0(n27168), .S1(n26693), .ZN(n23114) );
  MUX41 U12653 ( .I0(ram[10779]), .I1(ram[10771]), .I2(ram[10763]), .I3(
        ram[10755]), .S0(n27167), .S1(n26692), .ZN(n23116) );
  MUX41 U12654 ( .I0(ram[10875]), .I1(ram[10867]), .I2(ram[10859]), .I3(
        ram[10851]), .S0(n27168), .S1(n26693), .ZN(n23113) );
  MUX41 U12655 ( .I0(n23028), .I1(n23029), .I2(n23030), .I3(n23031), .S0(
        n26229), .S1(n26347), .ZN(n23027) );
  MUX41 U12656 ( .I0(ram[8763]), .I1(ram[8755]), .I2(ram[8747]), .I3(
        ram[8739]), .S0(n27163), .S1(n26688), .ZN(n23029) );
  MUX41 U12657 ( .I0(ram[8731]), .I1(ram[8723]), .I2(ram[8715]), .I3(
        ram[8707]), .S0(n27163), .S1(n26688), .ZN(n23031) );
  MUX41 U12658 ( .I0(ram[8827]), .I1(ram[8819]), .I2(ram[8811]), .I3(
        ram[8803]), .S0(n27163), .S1(n26688), .ZN(n23028) );
  MUX41 U12659 ( .I0(n23521), .I1(n23522), .I2(n23523), .I3(n23524), .S0(
        n26236), .S1(n26354), .ZN(n23520) );
  MUX41 U12660 ( .I0(ram[4156]), .I1(ram[4148]), .I2(ram[4140]), .I3(
        ram[4132]), .S0(n27191), .S1(n26716), .ZN(n23522) );
  MUX41 U12661 ( .I0(ram[4124]), .I1(ram[4116]), .I2(ram[4108]), .I3(
        ram[4100]), .S0(n27191), .S1(n26716), .ZN(n23524) );
  MUX41 U12662 ( .I0(ram[4220]), .I1(ram[4212]), .I2(ram[4204]), .I3(
        ram[4196]), .S0(n27191), .S1(n26716), .ZN(n23521) );
  MUX41 U12663 ( .I0(n23541), .I1(n23542), .I2(n23543), .I3(n23544), .S0(
        n26236), .S1(n26354), .ZN(n23540) );
  MUX41 U12664 ( .I0(ram[4668]), .I1(ram[4660]), .I2(ram[4652]), .I3(
        ram[4644]), .S0(n27192), .S1(n26717), .ZN(n23542) );
  MUX41 U12665 ( .I0(ram[4636]), .I1(ram[4628]), .I2(ram[4620]), .I3(
        ram[4612]), .S0(n27192), .S1(n26717), .ZN(n23544) );
  MUX41 U12666 ( .I0(ram[4732]), .I1(ram[4724]), .I2(ram[4716]), .I3(
        ram[4708]), .S0(n27192), .S1(n26717), .ZN(n23541) );
  MUX41 U12667 ( .I0(n23797), .I1(n23798), .I2(n23799), .I3(n23800), .S0(
        n26240), .S1(n26358), .ZN(n23796) );
  MUX41 U12668 ( .I0(ram[10812]), .I1(ram[10804]), .I2(ram[10796]), .I3(
        ram[10788]), .S0(n27207), .S1(n26732), .ZN(n23798) );
  MUX41 U12669 ( .I0(ram[10780]), .I1(ram[10772]), .I2(ram[10764]), .I3(
        ram[10756]), .S0(n27207), .S1(n26732), .ZN(n23800) );
  MUX41 U12670 ( .I0(ram[10876]), .I1(ram[10868]), .I2(ram[10860]), .I3(
        ram[10852]), .S0(n27207), .S1(n26732), .ZN(n23797) );
  MUX41 U12671 ( .I0(n23712), .I1(n23713), .I2(n23714), .I3(n23715), .S0(
        n26238), .S1(n26356), .ZN(n23711) );
  MUX41 U12672 ( .I0(ram[8764]), .I1(ram[8756]), .I2(ram[8748]), .I3(
        ram[8740]), .S0(n27202), .S1(n26727), .ZN(n23713) );
  MUX41 U12673 ( .I0(ram[8732]), .I1(ram[8724]), .I2(ram[8716]), .I3(
        ram[8708]), .S0(n27202), .S1(n26727), .ZN(n23715) );
  MUX41 U12674 ( .I0(ram[8828]), .I1(ram[8820]), .I2(ram[8812]), .I3(
        ram[8804]), .S0(n27202), .S1(n26727), .ZN(n23712) );
  MUX41 U12675 ( .I0(n24205), .I1(n24206), .I2(n24207), .I3(n24208), .S0(
        n26245), .S1(n26363), .ZN(n24204) );
  MUX41 U12676 ( .I0(ram[4157]), .I1(ram[4149]), .I2(ram[4141]), .I3(
        ram[4133]), .S0(n27230), .S1(n26755), .ZN(n24206) );
  MUX41 U12677 ( .I0(ram[4125]), .I1(ram[4117]), .I2(ram[4109]), .I3(
        ram[4101]), .S0(n27230), .S1(n26755), .ZN(n24208) );
  MUX41 U12678 ( .I0(ram[4221]), .I1(ram[4213]), .I2(ram[4205]), .I3(
        ram[4197]), .S0(n27230), .S1(n26755), .ZN(n24205) );
  MUX41 U12679 ( .I0(n24225), .I1(n24226), .I2(n24227), .I3(n24228), .S0(
        n26246), .S1(n26364), .ZN(n24224) );
  MUX41 U12680 ( .I0(ram[4669]), .I1(ram[4661]), .I2(ram[4653]), .I3(
        ram[4645]), .S0(n27232), .S1(n26757), .ZN(n24226) );
  MUX41 U12681 ( .I0(ram[4637]), .I1(ram[4629]), .I2(ram[4621]), .I3(
        ram[4613]), .S0(n27231), .S1(n26756), .ZN(n24228) );
  MUX41 U12682 ( .I0(ram[4733]), .I1(ram[4725]), .I2(ram[4717]), .I3(
        ram[4709]), .S0(n27232), .S1(n26757), .ZN(n24225) );
  MUX41 U12683 ( .I0(n24481), .I1(n24482), .I2(n24483), .I3(n24484), .S0(
        n26249), .S1(n26367), .ZN(n24480) );
  MUX41 U12684 ( .I0(ram[10813]), .I1(ram[10805]), .I2(ram[10797]), .I3(
        ram[10789]), .S0(n27246), .S1(n26771), .ZN(n24482) );
  MUX41 U12685 ( .I0(ram[10781]), .I1(ram[10773]), .I2(ram[10765]), .I3(
        ram[10757]), .S0(n27246), .S1(n26771), .ZN(n24484) );
  MUX41 U12686 ( .I0(ram[10877]), .I1(ram[10869]), .I2(ram[10861]), .I3(
        ram[10853]), .S0(n27246), .S1(n26771), .ZN(n24481) );
  MUX41 U12687 ( .I0(n24396), .I1(n24397), .I2(n24398), .I3(n24399), .S0(
        n26248), .S1(n26366), .ZN(n24395) );
  MUX41 U12688 ( .I0(ram[8765]), .I1(ram[8757]), .I2(ram[8749]), .I3(
        ram[8741]), .S0(n27241), .S1(n26766), .ZN(n24397) );
  MUX41 U12689 ( .I0(ram[8733]), .I1(ram[8725]), .I2(ram[8717]), .I3(
        ram[8709]), .S0(n27241), .S1(n26766), .ZN(n24399) );
  MUX41 U12690 ( .I0(ram[8829]), .I1(ram[8821]), .I2(ram[8813]), .I3(
        ram[8805]), .S0(n27242), .S1(n26767), .ZN(n24396) );
  MUX41 U12691 ( .I0(n24889), .I1(n24890), .I2(n24891), .I3(n24892), .S0(
        n26255), .S1(n26373), .ZN(n24888) );
  MUX41 U12692 ( .I0(ram[4158]), .I1(ram[4150]), .I2(ram[4142]), .I3(
        ram[4134]), .S0(n27270), .S1(n26795), .ZN(n24890) );
  MUX41 U12693 ( .I0(ram[4126]), .I1(ram[4118]), .I2(ram[4110]), .I3(
        ram[4102]), .S0(n27270), .S1(n26795), .ZN(n24892) );
  MUX41 U12694 ( .I0(ram[4222]), .I1(ram[4214]), .I2(ram[4206]), .I3(
        ram[4198]), .S0(n27270), .S1(n26795), .ZN(n24889) );
  MUX41 U12695 ( .I0(n24909), .I1(n24910), .I2(n24911), .I3(n24912), .S0(
        n26256), .S1(n26374), .ZN(n24908) );
  MUX41 U12696 ( .I0(ram[4670]), .I1(ram[4662]), .I2(ram[4654]), .I3(
        ram[4646]), .S0(n27271), .S1(n26796), .ZN(n24910) );
  MUX41 U12697 ( .I0(ram[4638]), .I1(ram[4630]), .I2(ram[4622]), .I3(
        ram[4614]), .S0(n27271), .S1(n26796), .ZN(n24912) );
  MUX41 U12698 ( .I0(ram[4734]), .I1(ram[4726]), .I2(ram[4718]), .I3(
        ram[4710]), .S0(n27271), .S1(n26796), .ZN(n24909) );
  MUX41 U12699 ( .I0(n25165), .I1(n25166), .I2(n25167), .I3(n25168), .S0(
        n26259), .S1(n26377), .ZN(n25164) );
  MUX41 U12700 ( .I0(ram[10814]), .I1(ram[10806]), .I2(ram[10798]), .I3(
        ram[10790]), .S0(n27286), .S1(n26811), .ZN(n25166) );
  MUX41 U12701 ( .I0(ram[10782]), .I1(ram[10774]), .I2(ram[10766]), .I3(
        ram[10758]), .S0(n27286), .S1(n26811), .ZN(n25168) );
  MUX41 U12702 ( .I0(ram[10878]), .I1(ram[10870]), .I2(ram[10862]), .I3(
        ram[10854]), .S0(n27286), .S1(n26811), .ZN(n25165) );
  MUX41 U12703 ( .I0(n25080), .I1(n25081), .I2(n25082), .I3(n25083), .S0(
        n26258), .S1(n26376), .ZN(n25079) );
  MUX41 U12704 ( .I0(ram[8766]), .I1(ram[8758]), .I2(ram[8750]), .I3(
        ram[8742]), .S0(n27281), .S1(n26806), .ZN(n25081) );
  MUX41 U12705 ( .I0(ram[8734]), .I1(ram[8726]), .I2(ram[8718]), .I3(
        ram[8710]), .S0(n27281), .S1(n26806), .ZN(n25083) );
  MUX41 U12706 ( .I0(ram[8830]), .I1(ram[8822]), .I2(ram[8814]), .I3(
        ram[8806]), .S0(n27281), .S1(n26806), .ZN(n25080) );
  MUX41 U12707 ( .I0(n25573), .I1(n25574), .I2(n25575), .I3(n25576), .S0(
        n26265), .S1(n26383), .ZN(n25572) );
  MUX41 U12708 ( .I0(ram[4159]), .I1(ram[4151]), .I2(ram[4143]), .I3(
        ram[4135]), .S0(n27309), .S1(n26834), .ZN(n25574) );
  MUX41 U12709 ( .I0(ram[4127]), .I1(ram[4119]), .I2(ram[4111]), .I3(
        ram[4103]), .S0(n27309), .S1(n26834), .ZN(n25576) );
  MUX41 U12710 ( .I0(ram[4223]), .I1(ram[4215]), .I2(ram[4207]), .I3(
        ram[4199]), .S0(n27309), .S1(n26834), .ZN(n25573) );
  MUX41 U12711 ( .I0(n25593), .I1(n25594), .I2(n25595), .I3(n25596), .S0(
        n26265), .S1(n26383), .ZN(n25592) );
  MUX41 U12712 ( .I0(ram[4671]), .I1(ram[4663]), .I2(ram[4655]), .I3(
        ram[4647]), .S0(n27310), .S1(n26835), .ZN(n25594) );
  MUX41 U12713 ( .I0(ram[4639]), .I1(ram[4631]), .I2(ram[4623]), .I3(
        ram[4615]), .S0(n27310), .S1(n26835), .ZN(n25596) );
  MUX41 U12714 ( .I0(ram[4735]), .I1(ram[4727]), .I2(ram[4719]), .I3(
        ram[4711]), .S0(n27310), .S1(n26835), .ZN(n25593) );
  MUX41 U12715 ( .I0(n25849), .I1(n25850), .I2(n25851), .I3(n25852), .S0(
        n26269), .S1(n26387), .ZN(n25848) );
  MUX41 U12716 ( .I0(ram[10815]), .I1(ram[10807]), .I2(ram[10799]), .I3(
        ram[10791]), .S0(n27325), .S1(n26850), .ZN(n25850) );
  MUX41 U12717 ( .I0(ram[10783]), .I1(ram[10775]), .I2(ram[10767]), .I3(
        ram[10759]), .S0(n27325), .S1(n26850), .ZN(n25852) );
  MUX41 U12718 ( .I0(ram[10879]), .I1(ram[10871]), .I2(ram[10863]), .I3(
        ram[10855]), .S0(n27325), .S1(n26850), .ZN(n25849) );
  MUX41 U12719 ( .I0(n25764), .I1(n25765), .I2(n25766), .I3(n25767), .S0(
        n26268), .S1(n26386), .ZN(n25763) );
  MUX41 U12720 ( .I0(ram[8767]), .I1(ram[8759]), .I2(ram[8751]), .I3(
        ram[8743]), .S0(n27320), .S1(n26845), .ZN(n25765) );
  MUX41 U12721 ( .I0(ram[8735]), .I1(ram[8727]), .I2(ram[8719]), .I3(
        ram[8711]), .S0(n27320), .S1(n26845), .ZN(n25767) );
  MUX41 U12722 ( .I0(ram[8831]), .I1(ram[8823]), .I2(ram[8815]), .I3(
        ram[8807]), .S0(n27320), .S1(n26845), .ZN(n25764) );
  MUX41 U12723 ( .I0(ram[24]), .I1(ram[16]), .I2(ram[8]), .I3(ram[0]), 
        .S0(n27168), .S1(n26624), .ZN(n3194) );
  MUX41 U12724 ( .I0(n20639), .I1(n20640), .I2(n20641), .I3(n20642), .S0(
        n26194), .S1(n26312), .ZN(n20638) );
  MUX41 U12725 ( .I0(ram[696]), .I1(ram[688]), .I2(ram[680]), .I3(
        ram[672]), .S0(n27025), .S1(n26550), .ZN(n20640) );
  MUX41 U12726 ( .I0(ram[664]), .I1(ram[656]), .I2(ram[648]), .I3(
        ram[640]), .S0(n27025), .S1(n26550), .ZN(n20642) );
  MUX41 U12727 ( .I0(ram[760]), .I1(ram[752]), .I2(ram[744]), .I3(
        ram[736]), .S0(n27025), .S1(n26550), .ZN(n20639) );
  MUX41 U12728 ( .I0(ram[4024]), .I1(ram[4016]), .I2(ram[4008]), .I3(
        ram[4000]), .S0(n27033), .S1(n26558), .ZN(n20775) );
  MUX41 U12729 ( .I0(ram[3768]), .I1(ram[3760]), .I2(ram[3752]), .I3(
        ram[3744]), .S0(n27032), .S1(n26557), .ZN(n20765) );
  MUX41 U12730 ( .I0(ram[3640]), .I1(ram[3632]), .I2(ram[3624]), .I3(
        ram[3616]), .S0(n27032), .S1(n26557), .ZN(n20760) );
  MUX41 U12731 ( .I0(ram[2488]), .I1(ram[2480]), .I2(ram[2472]), .I3(
        ram[2464]), .S0(n27029), .S1(n26554), .ZN(n20715) );
  MUX41 U12732 ( .I0(ram[2232]), .I1(ram[2224]), .I2(ram[2216]), .I3(
        ram[2208]), .S0(n27029), .S1(n26554), .ZN(n20705) );
  MUX41 U12733 ( .I0(ram[2104]), .I1(ram[2096]), .I2(ram[2088]), .I3(
        ram[2080]), .S0(n27028), .S1(n26553), .ZN(n20700) );
  MUX41 U12734 ( .I0(ram[3000]), .I1(ram[2992]), .I2(ram[2984]), .I3(
        ram[2976]), .S0(n27031), .S1(n26556), .ZN(n20735) );
  MUX41 U12735 ( .I0(ram[2744]), .I1(ram[2736]), .I2(ram[2728]), .I3(
        ram[2720]), .S0(n27030), .S1(n26555), .ZN(n20725) );
  MUX41 U12736 ( .I0(ram[2616]), .I1(ram[2608]), .I2(ram[2600]), .I3(
        ram[2592]), .S0(n27030), .S1(n26555), .ZN(n20720) );
  MUX41 U12737 ( .I0(ram[1080]), .I1(ram[1072]), .I2(ram[1064]), .I3(
        ram[1056]), .S0(n27026), .S1(n26551), .ZN(n20655) );
  MUX41 U12738 ( .I0(ram[1976]), .I1(ram[1968]), .I2(ram[1960]), .I3(
        ram[1952]), .S0(n27028), .S1(n26553), .ZN(n20690) );
  MUX41 U12739 ( .I0(ram[1720]), .I1(ram[1712]), .I2(ram[1704]), .I3(
        ram[1696]), .S0(n27028), .S1(n26553), .ZN(n20680) );
  MUX41 U12740 ( .I0(ram[1592]), .I1(ram[1584]), .I2(ram[1576]), .I3(
        ram[1568]), .S0(n27027), .S1(n26552), .ZN(n20675) );
  MUX41 U12741 ( .I0(ram[440]), .I1(ram[432]), .I2(ram[424]), .I3(
        ram[416]), .S0(n27024), .S1(n26549), .ZN(n20630) );
  MUX41 U12742 ( .I0(ram[184]), .I1(ram[176]), .I2(ram[168]), .I3(
        ram[160]), .S0(n27024), .S1(n26549), .ZN(n3582) );
  MUX41 U12743 ( .I0(ram[56]), .I1(ram[48]), .I2(ram[40]), .I3(ram[32]), 
        .S0(n27024), .S1(n26549), .ZN(n2936) );
  MUX41 U12744 ( .I0(ram[4025]), .I1(ram[4017]), .I2(ram[4009]), .I3(
        ram[4001]), .S0(n27072), .S1(n26597), .ZN(n21459) );
  MUX41 U12745 ( .I0(ram[3769]), .I1(ram[3761]), .I2(ram[3753]), .I3(
        ram[3745]), .S0(n27072), .S1(n26597), .ZN(n21449) );
  MUX41 U12746 ( .I0(ram[3641]), .I1(ram[3633]), .I2(ram[3625]), .I3(
        ram[3617]), .S0(n27072), .S1(n26597), .ZN(n21444) );
  MUX41 U12747 ( .I0(ram[2489]), .I1(ram[2481]), .I2(ram[2473]), .I3(
        ram[2465]), .S0(n27069), .S1(n26594), .ZN(n21399) );
  MUX41 U12748 ( .I0(ram[2233]), .I1(ram[2225]), .I2(ram[2217]), .I3(
        ram[2209]), .S0(n27068), .S1(n26593), .ZN(n21389) );
  MUX41 U12749 ( .I0(ram[2105]), .I1(ram[2097]), .I2(ram[2089]), .I3(
        ram[2081]), .S0(n27068), .S1(n26593), .ZN(n21384) );
  MUX41 U12750 ( .I0(ram[3001]), .I1(ram[2993]), .I2(ram[2985]), .I3(
        ram[2977]), .S0(n27070), .S1(n26595), .ZN(n21419) );
  MUX41 U12751 ( .I0(ram[2745]), .I1(ram[2737]), .I2(ram[2729]), .I3(
        ram[2721]), .S0(n27069), .S1(n26594), .ZN(n21409) );
  MUX41 U12752 ( .I0(ram[2617]), .I1(ram[2609]), .I2(ram[2601]), .I3(
        ram[2593]), .S0(n27069), .S1(n26594), .ZN(n21404) );
  MUX41 U12753 ( .I0(ram[1081]), .I1(ram[1073]), .I2(ram[1065]), .I3(
        ram[1057]), .S0(n27065), .S1(n26590), .ZN(n21339) );
  MUX41 U12754 ( .I0(ram[1977]), .I1(ram[1969]), .I2(ram[1961]), .I3(
        ram[1953]), .S0(n27068), .S1(n26593), .ZN(n21374) );
  MUX41 U12755 ( .I0(ram[1721]), .I1(ram[1713]), .I2(ram[1705]), .I3(
        ram[1697]), .S0(n27067), .S1(n26592), .ZN(n21364) );
  MUX41 U12756 ( .I0(ram[1593]), .I1(ram[1585]), .I2(ram[1577]), .I3(
        ram[1569]), .S0(n27067), .S1(n26592), .ZN(n21359) );
  MUX41 U12757 ( .I0(ram[441]), .I1(ram[433]), .I2(ram[425]), .I3(
        ram[417]), .S0(n27064), .S1(n26589), .ZN(n21314) );
  MUX41 U12758 ( .I0(ram[185]), .I1(ram[177]), .I2(ram[169]), .I3(
        ram[161]), .S0(n27063), .S1(n26588), .ZN(n21304) );
  MUX41 U12759 ( .I0(ram[57]), .I1(ram[49]), .I2(ram[41]), .I3(ram[33]), 
        .S0(n27063), .S1(n26588), .ZN(n21299) );
  MUX41 U12760 ( .I0(ram[4026]), .I1(ram[4018]), .I2(ram[4010]), .I3(
        ram[4002]), .S0(n27112), .S1(n26637), .ZN(n22143) );
  MUX41 U12761 ( .I0(ram[3770]), .I1(ram[3762]), .I2(ram[3754]), .I3(
        ram[3746]), .S0(n27111), .S1(n26636), .ZN(n22133) );
  MUX41 U12762 ( .I0(ram[3642]), .I1(ram[3634]), .I2(ram[3626]), .I3(
        ram[3618]), .S0(n27111), .S1(n26636), .ZN(n22128) );
  MUX41 U12763 ( .I0(ram[2490]), .I1(ram[2482]), .I2(ram[2474]), .I3(
        ram[2466]), .S0(n27108), .S1(n26633), .ZN(n22083) );
  MUX41 U12764 ( .I0(ram[2234]), .I1(ram[2226]), .I2(ram[2218]), .I3(
        ram[2210]), .S0(n27108), .S1(n26633), .ZN(n22073) );
  MUX41 U12765 ( .I0(ram[2106]), .I1(ram[2098]), .I2(ram[2090]), .I3(
        ram[2082]), .S0(n27107), .S1(n26632), .ZN(n22068) );
  MUX41 U12766 ( .I0(ram[3002]), .I1(ram[2994]), .I2(ram[2986]), .I3(
        ram[2978]), .S0(n27109), .S1(n26634), .ZN(n22103) );
  MUX41 U12767 ( .I0(ram[2746]), .I1(ram[2738]), .I2(ram[2730]), .I3(
        ram[2722]), .S0(n27109), .S1(n26634), .ZN(n22093) );
  MUX41 U12768 ( .I0(ram[2618]), .I1(ram[2610]), .I2(ram[2602]), .I3(
        ram[2594]), .S0(n27108), .S1(n26633), .ZN(n22088) );
  MUX41 U12769 ( .I0(ram[1978]), .I1(ram[1970]), .I2(ram[1962]), .I3(
        ram[1954]), .S0(n27107), .S1(n26632), .ZN(n22058) );
  MUX41 U12770 ( .I0(ram[1722]), .I1(ram[1714]), .I2(ram[1706]), .I3(
        ram[1698]), .S0(n27106), .S1(n26631), .ZN(n22048) );
  MUX41 U12771 ( .I0(ram[1594]), .I1(ram[1586]), .I2(ram[1578]), .I3(
        ram[1570]), .S0(n27106), .S1(n26631), .ZN(n22043) );
  MUX41 U12772 ( .I0(ram[442]), .I1(ram[434]), .I2(ram[426]), .I3(
        ram[418]), .S0(n27103), .S1(n26628), .ZN(n21998) );
  MUX41 U12773 ( .I0(ram[186]), .I1(ram[178]), .I2(ram[170]), .I3(
        ram[162]), .S0(n27103), .S1(n26628), .ZN(n21988) );
  MUX41 U12774 ( .I0(ram[58]), .I1(ram[50]), .I2(ram[42]), .I3(ram[34]), 
        .S0(n27102), .S1(n26627), .ZN(n21983) );
  MUX41 U12775 ( .I0(ram[4027]), .I1(ram[4019]), .I2(ram[4011]), .I3(
        ram[4003]), .S0(n27151), .S1(n26676), .ZN(n22827) );
  MUX41 U12776 ( .I0(ram[3771]), .I1(ram[3763]), .I2(ram[3755]), .I3(
        ram[3747]), .S0(n27151), .S1(n26676), .ZN(n22817) );
  MUX41 U12777 ( .I0(ram[3643]), .I1(ram[3635]), .I2(ram[3627]), .I3(
        ram[3619]), .S0(n27150), .S1(n26675), .ZN(n22812) );
  MUX41 U12778 ( .I0(ram[2491]), .I1(ram[2483]), .I2(ram[2475]), .I3(
        ram[2467]), .S0(n27148), .S1(n26673), .ZN(n22767) );
  MUX41 U12779 ( .I0(ram[2235]), .I1(ram[2227]), .I2(ram[2219]), .I3(
        ram[2211]), .S0(n27147), .S1(n26672), .ZN(n22757) );
  MUX41 U12780 ( .I0(ram[2107]), .I1(ram[2099]), .I2(ram[2091]), .I3(
        ram[2083]), .S0(n27147), .S1(n26672), .ZN(n22752) );
  MUX41 U12781 ( .I0(ram[3003]), .I1(ram[2995]), .I2(ram[2987]), .I3(
        ram[2979]), .S0(n27149), .S1(n26674), .ZN(n22787) );
  MUX41 U12782 ( .I0(ram[2747]), .I1(ram[2739]), .I2(ram[2731]), .I3(
        ram[2723]), .S0(n27148), .S1(n26673), .ZN(n22777) );
  MUX41 U12783 ( .I0(ram[2619]), .I1(ram[2611]), .I2(ram[2603]), .I3(
        ram[2595]), .S0(n27148), .S1(n26673), .ZN(n22772) );
  MUX41 U12784 ( .I0(ram[1979]), .I1(ram[1971]), .I2(ram[1963]), .I3(
        ram[1955]), .S0(n27146), .S1(n26671), .ZN(n22742) );
  MUX41 U12785 ( .I0(ram[1723]), .I1(ram[1715]), .I2(ram[1707]), .I3(
        ram[1699]), .S0(n27146), .S1(n26671), .ZN(n22732) );
  MUX41 U12786 ( .I0(ram[1595]), .I1(ram[1587]), .I2(ram[1579]), .I3(
        ram[1571]), .S0(n27145), .S1(n26670), .ZN(n22727) );
  MUX41 U12787 ( .I0(ram[443]), .I1(ram[435]), .I2(ram[427]), .I3(
        ram[419]), .S0(n27143), .S1(n26668), .ZN(n22682) );
  MUX41 U12788 ( .I0(ram[187]), .I1(ram[179]), .I2(ram[171]), .I3(
        ram[163]), .S0(n27142), .S1(n26667), .ZN(n22672) );
  MUX41 U12789 ( .I0(ram[59]), .I1(ram[51]), .I2(ram[43]), .I3(ram[35]), 
        .S0(n27142), .S1(n26667), .ZN(n22667) );
  MUX41 U12790 ( .I0(ram[4028]), .I1(ram[4020]), .I2(ram[4012]), .I3(
        ram[4004]), .S0(n27191), .S1(n26716), .ZN(n23511) );
  MUX41 U12791 ( .I0(ram[3772]), .I1(ram[3764]), .I2(ram[3756]), .I3(
        ram[3748]), .S0(n27190), .S1(n26715), .ZN(n23501) );
  MUX41 U12792 ( .I0(ram[3644]), .I1(ram[3636]), .I2(ram[3628]), .I3(
        ram[3620]), .S0(n27190), .S1(n26715), .ZN(n23496) );
  MUX41 U12793 ( .I0(ram[2492]), .I1(ram[2484]), .I2(ram[2476]), .I3(
        ram[2468]), .S0(n27187), .S1(n26712), .ZN(n23451) );
  MUX41 U12794 ( .I0(ram[2236]), .I1(ram[2228]), .I2(ram[2220]), .I3(
        ram[2212]), .S0(n27186), .S1(n26711), .ZN(n23441) );
  MUX41 U12795 ( .I0(ram[2108]), .I1(ram[2100]), .I2(ram[2092]), .I3(
        ram[2084]), .S0(n27186), .S1(n26711), .ZN(n23436) );
  MUX41 U12796 ( .I0(ram[3004]), .I1(ram[2996]), .I2(ram[2988]), .I3(
        ram[2980]), .S0(n27188), .S1(n26713), .ZN(n23471) );
  MUX41 U12797 ( .I0(ram[2748]), .I1(ram[2740]), .I2(ram[2732]), .I3(
        ram[2724]), .S0(n27188), .S1(n26713), .ZN(n23461) );
  MUX41 U12798 ( .I0(ram[2620]), .I1(ram[2612]), .I2(ram[2604]), .I3(
        ram[2596]), .S0(n27187), .S1(n26712), .ZN(n23456) );
  MUX41 U12799 ( .I0(ram[1980]), .I1(ram[1972]), .I2(ram[1964]), .I3(
        ram[1956]), .S0(n27186), .S1(n26711), .ZN(n23426) );
  MUX41 U12800 ( .I0(ram[1724]), .I1(ram[1716]), .I2(ram[1708]), .I3(
        ram[1700]), .S0(n27185), .S1(n26710), .ZN(n23416) );
  MUX41 U12801 ( .I0(ram[1596]), .I1(ram[1588]), .I2(ram[1580]), .I3(
        ram[1572]), .S0(n27185), .S1(n26710), .ZN(n23411) );
  MUX41 U12802 ( .I0(ram[444]), .I1(ram[436]), .I2(ram[428]), .I3(
        ram[420]), .S0(n27182), .S1(n26707), .ZN(n23366) );
  MUX41 U12803 ( .I0(ram[188]), .I1(ram[180]), .I2(ram[172]), .I3(
        ram[164]), .S0(n27181), .S1(n26706), .ZN(n23356) );
  MUX41 U12804 ( .I0(ram[60]), .I1(ram[52]), .I2(ram[44]), .I3(ram[36]), 
        .S0(n27181), .S1(n26706), .ZN(n23351) );
  MUX41 U12805 ( .I0(ram[4029]), .I1(ram[4021]), .I2(ram[4013]), .I3(
        ram[4005]), .S0(n27230), .S1(n26755), .ZN(n24195) );
  MUX41 U12806 ( .I0(ram[3773]), .I1(ram[3765]), .I2(ram[3757]), .I3(
        ram[3749]), .S0(n27229), .S1(n26754), .ZN(n24185) );
  MUX41 U12807 ( .I0(ram[3645]), .I1(ram[3637]), .I2(ram[3629]), .I3(
        ram[3621]), .S0(n27229), .S1(n26754), .ZN(n24180) );
  MUX41 U12808 ( .I0(ram[2493]), .I1(ram[2485]), .I2(ram[2477]), .I3(
        ram[2469]), .S0(n27226), .S1(n26751), .ZN(n24135) );
  MUX41 U12809 ( .I0(ram[2237]), .I1(ram[2229]), .I2(ram[2221]), .I3(
        ram[2213]), .S0(n27226), .S1(n26751), .ZN(n24125) );
  MUX41 U12810 ( .I0(ram[2109]), .I1(ram[2101]), .I2(ram[2093]), .I3(
        ram[2085]), .S0(n27225), .S1(n26750), .ZN(n24120) );
  MUX41 U12811 ( .I0(ram[3005]), .I1(ram[2997]), .I2(ram[2989]), .I3(
        ram[2981]), .S0(n27228), .S1(n26753), .ZN(n24155) );
  MUX41 U12812 ( .I0(ram[2749]), .I1(ram[2741]), .I2(ram[2733]), .I3(
        ram[2725]), .S0(n27227), .S1(n26752), .ZN(n24145) );
  MUX41 U12813 ( .I0(ram[2621]), .I1(ram[2613]), .I2(ram[2605]), .I3(
        ram[2597]), .S0(n27227), .S1(n26752), .ZN(n24140) );
  MUX41 U12814 ( .I0(ram[1981]), .I1(ram[1973]), .I2(ram[1965]), .I3(
        ram[1957]), .S0(n27225), .S1(n26750), .ZN(n24110) );
  MUX41 U12815 ( .I0(ram[1725]), .I1(ram[1717]), .I2(ram[1709]), .I3(
        ram[1701]), .S0(n27224), .S1(n26749), .ZN(n24100) );
  MUX41 U12816 ( .I0(ram[1597]), .I1(ram[1589]), .I2(ram[1581]), .I3(
        ram[1573]), .S0(n27224), .S1(n26749), .ZN(n24095) );
  MUX41 U12817 ( .I0(ram[445]), .I1(ram[437]), .I2(ram[429]), .I3(
        ram[421]), .S0(n27221), .S1(n26746), .ZN(n24050) );
  MUX41 U12818 ( .I0(ram[189]), .I1(ram[181]), .I2(ram[173]), .I3(
        ram[165]), .S0(n27221), .S1(n26746), .ZN(n24040) );
  MUX41 U12819 ( .I0(ram[61]), .I1(ram[53]), .I2(ram[45]), .I3(ram[37]), 
        .S0(n27220), .S1(n26745), .ZN(n24035) );
  MUX41 U12820 ( .I0(ram[4030]), .I1(ram[4022]), .I2(ram[4014]), .I3(
        ram[4006]), .S0(n27269), .S1(n26794), .ZN(n24879) );
  MUX41 U12821 ( .I0(ram[3774]), .I1(ram[3766]), .I2(ram[3758]), .I3(
        ram[3750]), .S0(n27269), .S1(n26794), .ZN(n24869) );
  MUX41 U12822 ( .I0(ram[3646]), .I1(ram[3638]), .I2(ram[3630]), .I3(
        ram[3622]), .S0(n27268), .S1(n26793), .ZN(n24864) );
  MUX41 U12823 ( .I0(ram[2494]), .I1(ram[2486]), .I2(ram[2478]), .I3(
        ram[2470]), .S0(n27266), .S1(n26791), .ZN(n24819) );
  MUX41 U12824 ( .I0(ram[2238]), .I1(ram[2230]), .I2(ram[2222]), .I3(
        ram[2214]), .S0(n27265), .S1(n26790), .ZN(n24809) );
  MUX41 U12825 ( .I0(ram[2110]), .I1(ram[2102]), .I2(ram[2094]), .I3(
        ram[2086]), .S0(n27265), .S1(n26790), .ZN(n24804) );
  MUX41 U12826 ( .I0(ram[3006]), .I1(ram[2998]), .I2(ram[2990]), .I3(
        ram[2982]), .S0(n27267), .S1(n26792), .ZN(n24839) );
  MUX41 U12827 ( .I0(ram[2750]), .I1(ram[2742]), .I2(ram[2734]), .I3(
        ram[2726]), .S0(n27266), .S1(n26791), .ZN(n24829) );
  MUX41 U12828 ( .I0(ram[2622]), .I1(ram[2614]), .I2(ram[2606]), .I3(
        ram[2598]), .S0(n27266), .S1(n26791), .ZN(n24824) );
  MUX41 U12829 ( .I0(ram[1982]), .I1(ram[1974]), .I2(ram[1966]), .I3(
        ram[1958]), .S0(n27264), .S1(n26789), .ZN(n24794) );
  MUX41 U12830 ( .I0(ram[1726]), .I1(ram[1718]), .I2(ram[1710]), .I3(
        ram[1702]), .S0(n27264), .S1(n26789), .ZN(n24784) );
  MUX41 U12831 ( .I0(ram[1598]), .I1(ram[1590]), .I2(ram[1582]), .I3(
        ram[1574]), .S0(n27264), .S1(n26789), .ZN(n24779) );
  MUX41 U12832 ( .I0(ram[446]), .I1(ram[438]), .I2(ram[430]), .I3(
        ram[422]), .S0(n27261), .S1(n26786), .ZN(n24734) );
  MUX41 U12833 ( .I0(ram[190]), .I1(ram[182]), .I2(ram[174]), .I3(
        ram[166]), .S0(n27260), .S1(n26785), .ZN(n24724) );
  MUX41 U12834 ( .I0(ram[62]), .I1(ram[54]), .I2(ram[46]), .I3(ram[38]), 
        .S0(n27260), .S1(n26785), .ZN(n24719) );
  MUX41 U12835 ( .I0(ram[4031]), .I1(ram[4023]), .I2(ram[4015]), .I3(
        ram[4007]), .S0(n27309), .S1(n26834), .ZN(n25563) );
  MUX41 U12836 ( .I0(ram[3775]), .I1(ram[3767]), .I2(ram[3759]), .I3(
        ram[3751]), .S0(n27308), .S1(n26833), .ZN(n25553) );
  MUX41 U12837 ( .I0(ram[3647]), .I1(ram[3639]), .I2(ram[3631]), .I3(
        ram[3623]), .S0(n27308), .S1(n26833), .ZN(n25548) );
  MUX41 U12838 ( .I0(ram[2495]), .I1(ram[2487]), .I2(ram[2479]), .I3(
        ram[2471]), .S0(n27305), .S1(n26830), .ZN(n25503) );
  MUX41 U12839 ( .I0(ram[2239]), .I1(ram[2231]), .I2(ram[2223]), .I3(
        ram[2215]), .S0(n27304), .S1(n26829), .ZN(n25493) );
  MUX41 U12840 ( .I0(ram[2111]), .I1(ram[2103]), .I2(ram[2095]), .I3(
        ram[2087]), .S0(n27304), .S1(n26829), .ZN(n25488) );
  MUX41 U12841 ( .I0(ram[3007]), .I1(ram[2999]), .I2(ram[2991]), .I3(
        ram[2983]), .S0(n27306), .S1(n26831), .ZN(n25523) );
  MUX41 U12842 ( .I0(ram[2751]), .I1(ram[2743]), .I2(ram[2735]), .I3(
        ram[2727]), .S0(n27306), .S1(n26831), .ZN(n25513) );
  MUX41 U12843 ( .I0(ram[2623]), .I1(ram[2615]), .I2(ram[2607]), .I3(
        ram[2599]), .S0(n27305), .S1(n26830), .ZN(n25508) );
  MUX41 U12844 ( .I0(ram[1983]), .I1(ram[1975]), .I2(ram[1967]), .I3(
        ram[1959]), .S0(n27304), .S1(n26829), .ZN(n25478) );
  MUX41 U12845 ( .I0(ram[1727]), .I1(ram[1719]), .I2(ram[1711]), .I3(
        ram[1703]), .S0(n27303), .S1(n26828), .ZN(n25468) );
  MUX41 U12846 ( .I0(ram[1599]), .I1(ram[1591]), .I2(ram[1583]), .I3(
        ram[1575]), .S0(n27303), .S1(n26828), .ZN(n25463) );
  MUX41 U12847 ( .I0(ram[447]), .I1(ram[439]), .I2(ram[431]), .I3(
        ram[423]), .S0(n27300), .S1(n26825), .ZN(n25418) );
  MUX41 U12848 ( .I0(ram[191]), .I1(ram[183]), .I2(ram[175]), .I3(
        ram[167]), .S0(n27300), .S1(n26825), .ZN(n25408) );
  MUX41 U12849 ( .I0(ram[63]), .I1(ram[55]), .I2(ram[47]), .I3(ram[39]), 
        .S0(n27299), .S1(n26824), .ZN(n25403) );
  MUX41 U12850 ( .I0(ram[7224]), .I1(ram[7216]), .I2(ram[7208]), .I3(
        ram[7200]), .S0(n27041), .S1(n26566), .ZN(n20911) );
  MUX41 U12851 ( .I0(ram[5560]), .I1(ram[5552]), .I2(ram[5544]), .I3(
        ram[5536]), .S0(n27037), .S1(n26562), .ZN(n20841) );
  MUX41 U12852 ( .I0(ram[5304]), .I1(ram[5296]), .I2(ram[5288]), .I3(
        ram[5280]), .S0(n27036), .S1(n26561), .ZN(n20831) );
  MUX41 U12853 ( .I0(ram[5176]), .I1(ram[5168]), .I2(ram[5160]), .I3(
        ram[5152]), .S0(n27036), .S1(n26561), .ZN(n20826) );
  MUX41 U12854 ( .I0(ram[11448]), .I1(ram[11440]), .I2(ram[11432]), .I3(
        ram[11424]), .S0(n27051), .S1(n26576), .ZN(n21087) );
  MUX41 U12855 ( .I0(ram[11320]), .I1(ram[11312]), .I2(ram[11304]), .I3(
        ram[11296]), .S0(n27051), .S1(n26576), .ZN(n21082) );
  MUX41 U12856 ( .I0(ram[9400]), .I1(ram[9392]), .I2(ram[9384]), .I3(
        ram[9376]), .S0(n27046), .S1(n26571), .ZN(n21002) );
  MUX41 U12857 ( .I0(ram[9272]), .I1(ram[9264]), .I2(ram[9256]), .I3(
        ram[9248]), .S0(n27046), .S1(n26571), .ZN(n20997) );
  MUX41 U12858 ( .I0(ram[7225]), .I1(ram[7217]), .I2(ram[7209]), .I3(
        ram[7201]), .S0(n27080), .S1(n26605), .ZN(n21595) );
  MUX41 U12859 ( .I0(ram[5561]), .I1(ram[5553]), .I2(ram[5545]), .I3(
        ram[5537]), .S0(n27076), .S1(n26601), .ZN(n21525) );
  MUX41 U12860 ( .I0(ram[5305]), .I1(ram[5297]), .I2(ram[5289]), .I3(
        ram[5281]), .S0(n27076), .S1(n26601), .ZN(n21515) );
  MUX41 U12861 ( .I0(ram[5177]), .I1(ram[5169]), .I2(ram[5161]), .I3(
        ram[5153]), .S0(n27075), .S1(n26600), .ZN(n21510) );
  MUX41 U12862 ( .I0(ram[11449]), .I1(ram[11441]), .I2(ram[11433]), .I3(
        ram[11425]), .S0(n27090), .S1(n26615), .ZN(n21771) );
  MUX41 U12863 ( .I0(ram[11321]), .I1(ram[11313]), .I2(ram[11305]), .I3(
        ram[11297]), .S0(n27090), .S1(n26615), .ZN(n21766) );
  MUX41 U12864 ( .I0(ram[9401]), .I1(ram[9393]), .I2(ram[9385]), .I3(
        ram[9377]), .S0(n27085), .S1(n26610), .ZN(n21686) );
  MUX41 U12865 ( .I0(ram[9273]), .I1(ram[9265]), .I2(ram[9257]), .I3(
        ram[9249]), .S0(n27085), .S1(n26610), .ZN(n21681) );
  MUX41 U12866 ( .I0(ram[5562]), .I1(ram[5554]), .I2(ram[5546]), .I3(
        ram[5538]), .S0(n27116), .S1(n26641), .ZN(n22209) );
  MUX41 U12867 ( .I0(ram[5306]), .I1(ram[5298]), .I2(ram[5290]), .I3(
        ram[5282]), .S0(n27115), .S1(n26640), .ZN(n22199) );
  MUX41 U12868 ( .I0(ram[5178]), .I1(ram[5170]), .I2(ram[5162]), .I3(
        ram[5154]), .S0(n27115), .S1(n26640), .ZN(n22194) );
  MUX41 U12869 ( .I0(ram[11322]), .I1(ram[11314]), .I2(ram[11306]), .I3(
        ram[11298]), .S0(n27129), .S1(n26654), .ZN(n22450) );
  MUX41 U12870 ( .I0(ram[9402]), .I1(ram[9394]), .I2(ram[9386]), .I3(
        ram[9378]), .S0(n27125), .S1(n26650), .ZN(n22370) );
  MUX41 U12871 ( .I0(ram[9274]), .I1(ram[9266]), .I2(ram[9258]), .I3(
        ram[9250]), .S0(n27124), .S1(n26649), .ZN(n22365) );
  MUX41 U12872 ( .I0(ram[5563]), .I1(ram[5555]), .I2(ram[5547]), .I3(
        ram[5539]), .S0(n27155), .S1(n26680), .ZN(n22893) );
  MUX41 U12873 ( .I0(ram[5307]), .I1(ram[5299]), .I2(ram[5291]), .I3(
        ram[5283]), .S0(n27154), .S1(n26679), .ZN(n22883) );
  MUX41 U12874 ( .I0(ram[5179]), .I1(ram[5171]), .I2(ram[5163]), .I3(
        ram[5155]), .S0(n27154), .S1(n26679), .ZN(n22878) );
  MUX41 U12875 ( .I0(ram[11323]), .I1(ram[11315]), .I2(ram[11307]), .I3(
        ram[11299]), .S0(n27169), .S1(n26694), .ZN(n23134) );
  MUX41 U12876 ( .I0(ram[9403]), .I1(ram[9395]), .I2(ram[9387]), .I3(
        ram[9379]), .S0(n27164), .S1(n26689), .ZN(n23054) );
  MUX41 U12877 ( .I0(ram[9275]), .I1(ram[9267]), .I2(ram[9259]), .I3(
        ram[9251]), .S0(n27164), .S1(n26689), .ZN(n23049) );
  MUX41 U12878 ( .I0(ram[5564]), .I1(ram[5556]), .I2(ram[5548]), .I3(
        ram[5540]), .S0(n27194), .S1(n26719), .ZN(n23577) );
  MUX41 U12879 ( .I0(ram[5308]), .I1(ram[5300]), .I2(ram[5292]), .I3(
        ram[5284]), .S0(n27194), .S1(n26719), .ZN(n23567) );
  MUX41 U12880 ( .I0(ram[5180]), .I1(ram[5172]), .I2(ram[5164]), .I3(
        ram[5156]), .S0(n27193), .S1(n26718), .ZN(n23562) );
  MUX41 U12881 ( .I0(ram[11324]), .I1(ram[11316]), .I2(ram[11308]), .I3(
        ram[11300]), .S0(n27208), .S1(n26733), .ZN(n23818) );
  MUX41 U12882 ( .I0(ram[9404]), .I1(ram[9396]), .I2(ram[9388]), .I3(
        ram[9380]), .S0(n27204), .S1(n26729), .ZN(n23738) );
  MUX41 U12883 ( .I0(ram[9276]), .I1(ram[9268]), .I2(ram[9260]), .I3(
        ram[9252]), .S0(n27203), .S1(n26728), .ZN(n23733) );
  MUX41 U12884 ( .I0(ram[5565]), .I1(ram[5557]), .I2(ram[5549]), .I3(
        ram[5541]), .S0(n27234), .S1(n26759), .ZN(n24261) );
  MUX41 U12885 ( .I0(ram[5309]), .I1(ram[5301]), .I2(ram[5293]), .I3(
        ram[5285]), .S0(n27233), .S1(n26758), .ZN(n24251) );
  MUX41 U12886 ( .I0(ram[5181]), .I1(ram[5173]), .I2(ram[5165]), .I3(
        ram[5157]), .S0(n27233), .S1(n26758), .ZN(n24246) );
  MUX41 U12887 ( .I0(ram[11325]), .I1(ram[11317]), .I2(ram[11309]), .I3(
        ram[11301]), .S0(n27248), .S1(n26773), .ZN(n24502) );
  MUX41 U12888 ( .I0(ram[9405]), .I1(ram[9397]), .I2(ram[9389]), .I3(
        ram[9381]), .S0(n27243), .S1(n26768), .ZN(n24422) );
  MUX41 U12889 ( .I0(ram[9277]), .I1(ram[9269]), .I2(ram[9261]), .I3(
        ram[9253]), .S0(n27243), .S1(n26768), .ZN(n24417) );
  MUX41 U12890 ( .I0(ram[5566]), .I1(ram[5558]), .I2(ram[5550]), .I3(
        ram[5542]), .S0(n27273), .S1(n26798), .ZN(n24945) );
  MUX41 U12891 ( .I0(ram[5310]), .I1(ram[5302]), .I2(ram[5294]), .I3(
        ram[5286]), .S0(n27272), .S1(n26797), .ZN(n24935) );
  MUX41 U12892 ( .I0(ram[5182]), .I1(ram[5174]), .I2(ram[5166]), .I3(
        ram[5158]), .S0(n27272), .S1(n26797), .ZN(n24930) );
  MUX41 U12893 ( .I0(ram[11326]), .I1(ram[11318]), .I2(ram[11310]), .I3(
        ram[11302]), .S0(n27287), .S1(n26812), .ZN(n25186) );
  MUX41 U12894 ( .I0(ram[9406]), .I1(ram[9398]), .I2(ram[9390]), .I3(
        ram[9382]), .S0(n27282), .S1(n26807), .ZN(n25106) );
  MUX41 U12895 ( .I0(ram[9278]), .I1(ram[9270]), .I2(ram[9262]), .I3(
        ram[9254]), .S0(n27282), .S1(n26807), .ZN(n25101) );
  MUX41 U12896 ( .I0(ram[5567]), .I1(ram[5559]), .I2(ram[5551]), .I3(
        ram[5543]), .S0(n27312), .S1(n26837), .ZN(n25629) );
  MUX41 U12897 ( .I0(ram[5311]), .I1(ram[5303]), .I2(ram[5295]), .I3(
        ram[5287]), .S0(n27312), .S1(n26837), .ZN(n25619) );
  MUX41 U12898 ( .I0(ram[5183]), .I1(ram[5175]), .I2(ram[5167]), .I3(
        ram[5159]), .S0(n27312), .S1(n26837), .ZN(n25614) );
  MUX41 U12899 ( .I0(ram[11327]), .I1(ram[11319]), .I2(ram[11311]), .I3(
        ram[11303]), .S0(n27326), .S1(n26851), .ZN(n25870) );
  MUX41 U12900 ( .I0(ram[9407]), .I1(ram[9399]), .I2(ram[9391]), .I3(
        ram[9383]), .S0(n27322), .S1(n26847), .ZN(n25790) );
  MUX41 U12901 ( .I0(ram[9279]), .I1(ram[9271]), .I2(ram[9263]), .I3(
        ram[9255]), .S0(n27321), .S1(n26846), .ZN(n25785) );
  MUX41 U12902 ( .I0(n20790), .I1(n20791), .I2(n20792), .I3(n20793), .S0(
        n26196), .S1(n26314), .ZN(n20789) );
  MUX41 U12903 ( .I0(ram[4280]), .I1(ram[4272]), .I2(ram[4264]), .I3(
        ram[4256]), .S0(n27034), .S1(n26559), .ZN(n20791) );
  MUX41 U12904 ( .I0(ram[4248]), .I1(ram[4240]), .I2(ram[4232]), .I3(
        ram[4224]), .S0(n27034), .S1(n26559), .ZN(n20793) );
  MUX41 U12905 ( .I0(ram[4344]), .I1(ram[4336]), .I2(ram[4328]), .I3(
        ram[4320]), .S0(n27034), .S1(n26559), .ZN(n20790) );
  MUX41 U12906 ( .I0(n20810), .I1(n20811), .I2(n20812), .I3(n20813), .S0(
        n26197), .S1(n26315), .ZN(n20809) );
  MUX41 U12907 ( .I0(ram[4792]), .I1(ram[4784]), .I2(ram[4776]), .I3(
        ram[4768]), .S0(n27035), .S1(n26560), .ZN(n20811) );
  MUX41 U12908 ( .I0(ram[4760]), .I1(ram[4752]), .I2(ram[4744]), .I3(
        ram[4736]), .S0(n27035), .S1(n26560), .ZN(n20813) );
  MUX41 U12909 ( .I0(ram[4856]), .I1(ram[4848]), .I2(ram[4840]), .I3(
        ram[4832]), .S0(n27035), .S1(n26560), .ZN(n20810) );
  MUX41 U12910 ( .I0(n21066), .I1(n21067), .I2(n21068), .I3(n21069), .S0(
        n26200), .S1(n26318), .ZN(n21065) );
  MUX41 U12911 ( .I0(ram[10936]), .I1(ram[10928]), .I2(ram[10920]), .I3(
        ram[10912]), .S0(n27050), .S1(n26575), .ZN(n21067) );
  MUX41 U12912 ( .I0(ram[10904]), .I1(ram[10896]), .I2(ram[10888]), .I3(
        ram[10880]), .S0(n27050), .S1(n26575), .ZN(n21069) );
  MUX41 U12913 ( .I0(ram[11000]), .I1(ram[10992]), .I2(ram[10984]), .I3(
        ram[10976]), .S0(n27050), .S1(n26575), .ZN(n21066) );
  MUX41 U12914 ( .I0(n20981), .I1(n20982), .I2(n20983), .I3(n20984), .S0(
        n26199), .S1(n26317), .ZN(n20980) );
  MUX41 U12915 ( .I0(ram[8888]), .I1(ram[8880]), .I2(ram[8872]), .I3(
        ram[8864]), .S0(n27045), .S1(n26570), .ZN(n20982) );
  MUX41 U12916 ( .I0(ram[8856]), .I1(ram[8848]), .I2(ram[8840]), .I3(
        ram[8832]), .S0(n27045), .S1(n26570), .ZN(n20984) );
  MUX41 U12917 ( .I0(ram[8952]), .I1(ram[8944]), .I2(ram[8936]), .I3(
        ram[8928]), .S0(n27045), .S1(n26570), .ZN(n20981) );
  MUX41 U12918 ( .I0(n21474), .I1(n21475), .I2(n21476), .I3(n21477), .S0(
        n26206), .S1(n26324), .ZN(n21473) );
  MUX41 U12919 ( .I0(ram[4281]), .I1(ram[4273]), .I2(ram[4265]), .I3(
        ram[4257]), .S0(n27073), .S1(n26598), .ZN(n21475) );
  MUX41 U12920 ( .I0(ram[4249]), .I1(ram[4241]), .I2(ram[4233]), .I3(
        ram[4225]), .S0(n27073), .S1(n26598), .ZN(n21477) );
  MUX41 U12921 ( .I0(ram[4345]), .I1(ram[4337]), .I2(ram[4329]), .I3(
        ram[4321]), .S0(n27073), .S1(n26598), .ZN(n21474) );
  MUX41 U12922 ( .I0(n21494), .I1(n21495), .I2(n21496), .I3(n21497), .S0(
        n26206), .S1(n26324), .ZN(n21493) );
  MUX41 U12923 ( .I0(ram[4793]), .I1(ram[4785]), .I2(ram[4777]), .I3(
        ram[4769]), .S0(n27074), .S1(n26599), .ZN(n21495) );
  MUX41 U12924 ( .I0(ram[4761]), .I1(ram[4753]), .I2(ram[4745]), .I3(
        ram[4737]), .S0(n27074), .S1(n26599), .ZN(n21497) );
  MUX41 U12925 ( .I0(ram[4857]), .I1(ram[4849]), .I2(ram[4841]), .I3(
        ram[4833]), .S0(n27074), .S1(n26599), .ZN(n21494) );
  MUX41 U12926 ( .I0(n21750), .I1(n21751), .I2(n21752), .I3(n21753), .S0(
        n26210), .S1(n26328), .ZN(n21749) );
  MUX41 U12927 ( .I0(ram[10937]), .I1(ram[10929]), .I2(ram[10921]), .I3(
        ram[10913]), .S0(n27089), .S1(n26614), .ZN(n21751) );
  MUX41 U12928 ( .I0(ram[10905]), .I1(ram[10897]), .I2(ram[10889]), .I3(
        ram[10881]), .S0(n27089), .S1(n26614), .ZN(n21753) );
  MUX41 U12929 ( .I0(ram[11001]), .I1(ram[10993]), .I2(ram[10985]), .I3(
        ram[10977]), .S0(n27089), .S1(n26614), .ZN(n21750) );
  MUX41 U12930 ( .I0(n21665), .I1(n21666), .I2(n21667), .I3(n21668), .S0(
        n26209), .S1(n26327), .ZN(n21664) );
  MUX41 U12931 ( .I0(ram[8889]), .I1(ram[8881]), .I2(ram[8873]), .I3(
        ram[8865]), .S0(n27084), .S1(n26609), .ZN(n21666) );
  MUX41 U12932 ( .I0(ram[8857]), .I1(ram[8849]), .I2(ram[8841]), .I3(
        ram[8833]), .S0(n27084), .S1(n26609), .ZN(n21668) );
  MUX41 U12933 ( .I0(ram[8953]), .I1(ram[8945]), .I2(ram[8937]), .I3(
        ram[8929]), .S0(n27084), .S1(n26609), .ZN(n21665) );
  MUX41 U12934 ( .I0(n22158), .I1(n22159), .I2(n22160), .I3(n22161), .S0(
        n26216), .S1(n26334), .ZN(n22157) );
  MUX41 U12935 ( .I0(ram[4282]), .I1(ram[4274]), .I2(ram[4266]), .I3(
        ram[4258]), .S0(n27112), .S1(n26637), .ZN(n22159) );
  MUX41 U12936 ( .I0(ram[4250]), .I1(ram[4242]), .I2(ram[4234]), .I3(
        ram[4226]), .S0(n27112), .S1(n26637), .ZN(n22161) );
  MUX41 U12937 ( .I0(ram[4346]), .I1(ram[4338]), .I2(ram[4330]), .I3(
        ram[4322]), .S0(n27113), .S1(n26638), .ZN(n22158) );
  MUX41 U12938 ( .I0(n22178), .I1(n22179), .I2(n22180), .I3(n22181), .S0(
        n26216), .S1(n26334), .ZN(n22177) );
  MUX41 U12939 ( .I0(ram[4794]), .I1(ram[4786]), .I2(ram[4778]), .I3(
        ram[4770]), .S0(n27114), .S1(n26639), .ZN(n22179) );
  MUX41 U12940 ( .I0(ram[4762]), .I1(ram[4754]), .I2(ram[4746]), .I3(
        ram[4738]), .S0(n27114), .S1(n26639), .ZN(n22181) );
  MUX41 U12941 ( .I0(ram[4858]), .I1(ram[4850]), .I2(ram[4842]), .I3(
        ram[4834]), .S0(n27114), .S1(n26639), .ZN(n22178) );
  MUX41 U12942 ( .I0(n22349), .I1(n22350), .I2(n22351), .I3(n22352), .S0(
        n26219), .S1(n26337), .ZN(n22348) );
  MUX41 U12943 ( .I0(ram[8890]), .I1(ram[8882]), .I2(ram[8874]), .I3(
        ram[8866]), .S0(n27124), .S1(n26649), .ZN(n22350) );
  MUX41 U12944 ( .I0(ram[8858]), .I1(ram[8850]), .I2(ram[8842]), .I3(
        ram[8834]), .S0(n27123), .S1(n26648), .ZN(n22352) );
  MUX41 U12945 ( .I0(ram[8954]), .I1(ram[8946]), .I2(ram[8938]), .I3(
        ram[8930]), .S0(n27124), .S1(n26649), .ZN(n22349) );
  MUX41 U12946 ( .I0(n22842), .I1(n22843), .I2(n22844), .I3(n22845), .S0(
        n26226), .S1(n26344), .ZN(n22841) );
  MUX41 U12947 ( .I0(ram[4283]), .I1(ram[4275]), .I2(ram[4267]), .I3(
        ram[4259]), .S0(n27152), .S1(n26677), .ZN(n22843) );
  MUX41 U12948 ( .I0(ram[4251]), .I1(ram[4243]), .I2(ram[4235]), .I3(
        ram[4227]), .S0(n27152), .S1(n26677), .ZN(n22845) );
  MUX41 U12949 ( .I0(ram[4347]), .I1(ram[4339]), .I2(ram[4331]), .I3(
        ram[4323]), .S0(n27152), .S1(n26677), .ZN(n22842) );
  MUX41 U12950 ( .I0(n22862), .I1(n22863), .I2(n22864), .I3(n22865), .S0(
        n26226), .S1(n26344), .ZN(n22861) );
  MUX41 U12951 ( .I0(ram[4795]), .I1(ram[4787]), .I2(ram[4779]), .I3(
        ram[4771]), .S0(n27153), .S1(n26678), .ZN(n22863) );
  MUX41 U12952 ( .I0(ram[4763]), .I1(ram[4755]), .I2(ram[4747]), .I3(
        ram[4739]), .S0(n27153), .S1(n26678), .ZN(n22865) );
  MUX41 U12953 ( .I0(ram[4859]), .I1(ram[4851]), .I2(ram[4843]), .I3(
        ram[4835]), .S0(n27153), .S1(n26678), .ZN(n22862) );
  MUX41 U12954 ( .I0(n23033), .I1(n23034), .I2(n23035), .I3(n23036), .S0(
        n26229), .S1(n26347), .ZN(n23032) );
  MUX41 U12955 ( .I0(ram[8891]), .I1(ram[8883]), .I2(ram[8875]), .I3(
        ram[8867]), .S0(n27163), .S1(n26688), .ZN(n23034) );
  MUX41 U12956 ( .I0(ram[8859]), .I1(ram[8851]), .I2(ram[8843]), .I3(
        ram[8835]), .S0(n27163), .S1(n26688), .ZN(n23036) );
  MUX41 U12957 ( .I0(ram[8955]), .I1(ram[8947]), .I2(ram[8939]), .I3(
        ram[8931]), .S0(n27163), .S1(n26688), .ZN(n23033) );
  MUX41 U12958 ( .I0(n23526), .I1(n23527), .I2(n23528), .I3(n23529), .S0(
        n26236), .S1(n26354), .ZN(n23525) );
  MUX41 U12959 ( .I0(ram[4284]), .I1(ram[4276]), .I2(ram[4268]), .I3(
        ram[4260]), .S0(n27191), .S1(n26716), .ZN(n23527) );
  MUX41 U12960 ( .I0(ram[4252]), .I1(ram[4244]), .I2(ram[4236]), .I3(
        ram[4228]), .S0(n27191), .S1(n26716), .ZN(n23529) );
  MUX41 U12961 ( .I0(ram[4348]), .I1(ram[4340]), .I2(ram[4332]), .I3(
        ram[4324]), .S0(n27191), .S1(n26716), .ZN(n23526) );
  MUX41 U12962 ( .I0(n23546), .I1(n23547), .I2(n23548), .I3(n23549), .S0(
        n26236), .S1(n26354), .ZN(n23545) );
  MUX41 U12963 ( .I0(ram[4796]), .I1(ram[4788]), .I2(ram[4780]), .I3(
        ram[4772]), .S0(n27192), .S1(n26717), .ZN(n23547) );
  MUX41 U12964 ( .I0(ram[4764]), .I1(ram[4756]), .I2(ram[4748]), .I3(
        ram[4740]), .S0(n27192), .S1(n26717), .ZN(n23549) );
  MUX41 U12965 ( .I0(ram[4860]), .I1(ram[4852]), .I2(ram[4844]), .I3(
        ram[4836]), .S0(n27193), .S1(n26718), .ZN(n23546) );
  MUX41 U12966 ( .I0(n23717), .I1(n23718), .I2(n23719), .I3(n23720), .S0(
        n26238), .S1(n26356), .ZN(n23716) );
  MUX41 U12967 ( .I0(ram[8892]), .I1(ram[8884]), .I2(ram[8876]), .I3(
        ram[8868]), .S0(n27202), .S1(n26727), .ZN(n23718) );
  MUX41 U12968 ( .I0(ram[8860]), .I1(ram[8852]), .I2(ram[8844]), .I3(
        ram[8836]), .S0(n27202), .S1(n26727), .ZN(n23720) );
  MUX41 U12969 ( .I0(ram[8956]), .I1(ram[8948]), .I2(ram[8940]), .I3(
        ram[8932]), .S0(n27202), .S1(n26727), .ZN(n23717) );
  MUX41 U12970 ( .I0(n24210), .I1(n24211), .I2(n24212), .I3(n24213), .S0(
        n26246), .S1(n26364), .ZN(n24209) );
  MUX41 U12971 ( .I0(ram[4285]), .I1(ram[4277]), .I2(ram[4269]), .I3(
        ram[4261]), .S0(n27231), .S1(n26756), .ZN(n24211) );
  MUX41 U12972 ( .I0(ram[4253]), .I1(ram[4245]), .I2(ram[4237]), .I3(
        ram[4229]), .S0(n27231), .S1(n26756), .ZN(n24213) );
  MUX41 U12973 ( .I0(ram[4349]), .I1(ram[4341]), .I2(ram[4333]), .I3(
        ram[4325]), .S0(n27231), .S1(n26756), .ZN(n24210) );
  MUX41 U12974 ( .I0(n24230), .I1(n24231), .I2(n24232), .I3(n24233), .S0(
        n26246), .S1(n26364), .ZN(n24229) );
  MUX41 U12975 ( .I0(ram[4797]), .I1(ram[4789]), .I2(ram[4781]), .I3(
        ram[4773]), .S0(n27232), .S1(n26757), .ZN(n24231) );
  MUX41 U12976 ( .I0(ram[4765]), .I1(ram[4757]), .I2(ram[4749]), .I3(
        ram[4741]), .S0(n27232), .S1(n26757), .ZN(n24233) );
  MUX41 U12977 ( .I0(ram[4861]), .I1(ram[4853]), .I2(ram[4845]), .I3(
        ram[4837]), .S0(n27232), .S1(n26757), .ZN(n24230) );
  MUX41 U12978 ( .I0(n24401), .I1(n24402), .I2(n24403), .I3(n24404), .S0(
        n26248), .S1(n26366), .ZN(n24400) );
  MUX41 U12979 ( .I0(ram[8893]), .I1(ram[8885]), .I2(ram[8877]), .I3(
        ram[8869]), .S0(n27242), .S1(n26767), .ZN(n24402) );
  MUX41 U12980 ( .I0(ram[8861]), .I1(ram[8853]), .I2(ram[8845]), .I3(
        ram[8837]), .S0(n27242), .S1(n26767), .ZN(n24404) );
  MUX41 U12981 ( .I0(ram[8957]), .I1(ram[8949]), .I2(ram[8941]), .I3(
        ram[8933]), .S0(n27242), .S1(n26767), .ZN(n24401) );
  MUX41 U12982 ( .I0(n24894), .I1(n24895), .I2(n24896), .I3(n24897), .S0(
        n26255), .S1(n26373), .ZN(n24893) );
  MUX41 U12983 ( .I0(ram[4286]), .I1(ram[4278]), .I2(ram[4270]), .I3(
        ram[4262]), .S0(n27270), .S1(n26795), .ZN(n24895) );
  MUX41 U12984 ( .I0(ram[4254]), .I1(ram[4246]), .I2(ram[4238]), .I3(
        ram[4230]), .S0(n27270), .S1(n26795), .ZN(n24897) );
  MUX41 U12985 ( .I0(ram[4350]), .I1(ram[4342]), .I2(ram[4334]), .I3(
        ram[4326]), .S0(n27270), .S1(n26795), .ZN(n24894) );
  MUX41 U12986 ( .I0(n24914), .I1(n24915), .I2(n24916), .I3(n24917), .S0(
        n26256), .S1(n26374), .ZN(n24913) );
  MUX41 U12987 ( .I0(ram[4798]), .I1(ram[4790]), .I2(ram[4782]), .I3(
        ram[4774]), .S0(n27271), .S1(n26796), .ZN(n24915) );
  MUX41 U12988 ( .I0(ram[4766]), .I1(ram[4758]), .I2(ram[4750]), .I3(
        ram[4742]), .S0(n27271), .S1(n26796), .ZN(n24917) );
  MUX41 U12989 ( .I0(ram[4862]), .I1(ram[4854]), .I2(ram[4846]), .I3(
        ram[4838]), .S0(n27271), .S1(n26796), .ZN(n24914) );
  MUX41 U12990 ( .I0(n25085), .I1(n25086), .I2(n25087), .I3(n25088), .S0(
        n26258), .S1(n26376), .ZN(n25084) );
  MUX41 U12991 ( .I0(ram[8894]), .I1(ram[8886]), .I2(ram[8878]), .I3(
        ram[8870]), .S0(n27281), .S1(n26806), .ZN(n25086) );
  MUX41 U12992 ( .I0(ram[8862]), .I1(ram[8854]), .I2(ram[8846]), .I3(
        ram[8838]), .S0(n27281), .S1(n26806), .ZN(n25088) );
  MUX41 U12993 ( .I0(ram[8958]), .I1(ram[8950]), .I2(ram[8942]), .I3(
        ram[8934]), .S0(n27281), .S1(n26806), .ZN(n25085) );
  MUX41 U12994 ( .I0(n25578), .I1(n25579), .I2(n25580), .I3(n25581), .S0(
        n26265), .S1(n26383), .ZN(n25577) );
  MUX41 U12995 ( .I0(ram[4287]), .I1(ram[4279]), .I2(ram[4271]), .I3(
        ram[4263]), .S0(n27309), .S1(n26834), .ZN(n25579) );
  MUX41 U12996 ( .I0(ram[4255]), .I1(ram[4247]), .I2(ram[4239]), .I3(
        ram[4231]), .S0(n27309), .S1(n26834), .ZN(n25581) );
  MUX41 U12997 ( .I0(ram[4351]), .I1(ram[4343]), .I2(ram[4335]), .I3(
        ram[4327]), .S0(n27310), .S1(n26835), .ZN(n25578) );
  MUX41 U12998 ( .I0(n25598), .I1(n25599), .I2(n25600), .I3(n25601), .S0(
        n26266), .S1(n26384), .ZN(n25597) );
  MUX41 U12999 ( .I0(ram[4799]), .I1(ram[4791]), .I2(ram[4783]), .I3(
        ram[4775]), .S0(n27311), .S1(n26836), .ZN(n25599) );
  MUX41 U13000 ( .I0(ram[4767]), .I1(ram[4759]), .I2(ram[4751]), .I3(
        ram[4743]), .S0(n27311), .S1(n26836), .ZN(n25601) );
  MUX41 U13001 ( .I0(ram[4863]), .I1(ram[4855]), .I2(ram[4847]), .I3(
        ram[4839]), .S0(n27311), .S1(n26836), .ZN(n25598) );
  MUX41 U13002 ( .I0(n25769), .I1(n25770), .I2(n25771), .I3(n25772), .S0(
        n26268), .S1(n26386), .ZN(n25768) );
  MUX41 U13003 ( .I0(ram[8895]), .I1(ram[8887]), .I2(ram[8879]), .I3(
        ram[8871]), .S0(n27320), .S1(n26845), .ZN(n25770) );
  MUX41 U13004 ( .I0(ram[8863]), .I1(ram[8855]), .I2(ram[8847]), .I3(
        ram[8839]), .S0(n27320), .S1(n26845), .ZN(n25772) );
  MUX41 U13005 ( .I0(ram[8959]), .I1(ram[8951]), .I2(ram[8943]), .I3(
        ram[8935]), .S0(n27321), .S1(n26846), .ZN(n25769) );
  MUX41 U13006 ( .I0(ram[728]), .I1(ram[720]), .I2(ram[712]), .I3(
        ram[704]), .S0(n27025), .S1(n26550), .ZN(n20641) );
  MUX41 U13007 ( .I0(ram[600]), .I1(ram[592]), .I2(ram[584]), .I3(
        ram[576]), .S0(n27025), .S1(n26550), .ZN(n20636) );
  MUX41 U13008 ( .I0(ram[601]), .I1(ram[593]), .I2(ram[585]), .I3(
        ram[577]), .S0(n27064), .S1(n26589), .ZN(n21320) );
  MUX41 U13009 ( .I0(ram[6744]), .I1(ram[6736]), .I2(ram[6728]), .I3(
        ram[6720]), .S0(n27040), .S1(n26565), .ZN(n20892) );
  MUX41 U13010 ( .I0(ram[4312]), .I1(ram[4304]), .I2(ram[4296]), .I3(
        ram[4288]), .S0(n27034), .S1(n26559), .ZN(n20792) );
  MUX41 U13011 ( .I0(ram[4184]), .I1(ram[4176]), .I2(ram[4168]), .I3(
        ram[4160]), .S0(n27033), .S1(n26558), .ZN(n20787) );
  MUX41 U13012 ( .I0(ram[5080]), .I1(ram[5072]), .I2(ram[5064]), .I3(
        ram[5056]), .S0(n27036), .S1(n26561), .ZN(n20822) );
  MUX41 U13013 ( .I0(ram[4824]), .I1(ram[4816]), .I2(ram[4808]), .I3(
        ram[4800]), .S0(n27035), .S1(n26560), .ZN(n20812) );
  MUX41 U13014 ( .I0(ram[4696]), .I1(ram[4688]), .I2(ram[4680]), .I3(
        ram[4672]), .S0(n27035), .S1(n26560), .ZN(n20807) );
  MUX41 U13015 ( .I0(ram[10968]), .I1(ram[10960]), .I2(ram[10952]), .I3(
        ram[10944]), .S0(n27050), .S1(n26575), .ZN(n21068) );
  MUX41 U13016 ( .I0(ram[10840]), .I1(ram[10832]), .I2(ram[10824]), .I3(
        ram[10816]), .S0(n27049), .S1(n26574), .ZN(n21063) );
  MUX41 U13017 ( .I0(ram[8280]), .I1(ram[8272]), .I2(ram[8264]), .I3(
        ram[8256]), .S0(n27043), .S1(n26568), .ZN(n20958) );
  MUX41 U13018 ( .I0(ram[8920]), .I1(ram[8912]), .I2(ram[8904]), .I3(
        ram[8896]), .S0(n27045), .S1(n26570), .ZN(n20983) );
  MUX41 U13019 ( .I0(ram[8792]), .I1(ram[8784]), .I2(ram[8776]), .I3(
        ram[8768]), .S0(n27045), .S1(n26570), .ZN(n20978) );
  MUX41 U13020 ( .I0(ram[6745]), .I1(ram[6737]), .I2(ram[6729]), .I3(
        ram[6721]), .S0(n27079), .S1(n26604), .ZN(n21576) );
  MUX41 U13021 ( .I0(ram[4313]), .I1(ram[4305]), .I2(ram[4297]), .I3(
        ram[4289]), .S0(n27073), .S1(n26598), .ZN(n21476) );
  MUX41 U13022 ( .I0(ram[4185]), .I1(ram[4177]), .I2(ram[4169]), .I3(
        ram[4161]), .S0(n27073), .S1(n26598), .ZN(n21471) );
  MUX41 U13023 ( .I0(ram[5081]), .I1(ram[5073]), .I2(ram[5065]), .I3(
        ram[5057]), .S0(n27075), .S1(n26600), .ZN(n21506) );
  MUX41 U13024 ( .I0(ram[4825]), .I1(ram[4817]), .I2(ram[4809]), .I3(
        ram[4801]), .S0(n27074), .S1(n26599), .ZN(n21496) );
  MUX41 U13025 ( .I0(ram[4697]), .I1(ram[4689]), .I2(ram[4681]), .I3(
        ram[4673]), .S0(n27074), .S1(n26599), .ZN(n21491) );
  MUX41 U13026 ( .I0(ram[10969]), .I1(ram[10961]), .I2(ram[10953]), .I3(
        ram[10945]), .S0(n27089), .S1(n26614), .ZN(n21752) );
  MUX41 U13027 ( .I0(ram[10841]), .I1(ram[10833]), .I2(ram[10825]), .I3(
        ram[10817]), .S0(n27089), .S1(n26614), .ZN(n21747) );
  MUX41 U13028 ( .I0(ram[8281]), .I1(ram[8273]), .I2(ram[8265]), .I3(
        ram[8257]), .S0(n27083), .S1(n26608), .ZN(n21642) );
  MUX41 U13029 ( .I0(ram[8921]), .I1(ram[8913]), .I2(ram[8905]), .I3(
        ram[8897]), .S0(n27084), .S1(n26609), .ZN(n21667) );
  MUX41 U13030 ( .I0(ram[8793]), .I1(ram[8785]), .I2(ram[8777]), .I3(
        ram[8769]), .S0(n27084), .S1(n26609), .ZN(n21662) );
  MUX41 U13031 ( .I0(ram[4314]), .I1(ram[4306]), .I2(ram[4298]), .I3(
        ram[4290]), .S0(n27113), .S1(n26638), .ZN(n22160) );
  MUX41 U13032 ( .I0(ram[4186]), .I1(ram[4178]), .I2(ram[4170]), .I3(
        ram[4162]), .S0(n27112), .S1(n26637), .ZN(n22155) );
  MUX41 U13033 ( .I0(ram[5082]), .I1(ram[5074]), .I2(ram[5066]), .I3(
        ram[5058]), .S0(n27114), .S1(n26639), .ZN(n22190) );
  MUX41 U13034 ( .I0(ram[4826]), .I1(ram[4818]), .I2(ram[4810]), .I3(
        ram[4802]), .S0(n27114), .S1(n26639), .ZN(n22180) );
  MUX41 U13035 ( .I0(ram[4698]), .I1(ram[4690]), .I2(ram[4682]), .I3(
        ram[4674]), .S0(n27113), .S1(n26638), .ZN(n22175) );
  MUX41 U13036 ( .I0(ram[10842]), .I1(ram[10834]), .I2(ram[10826]), .I3(
        ram[10818]), .S0(n27128), .S1(n26653), .ZN(n22431) );
  MUX41 U13037 ( .I0(ram[8922]), .I1(ram[8914]), .I2(ram[8906]), .I3(
        ram[8898]), .S0(n27124), .S1(n26649), .ZN(n22351) );
  MUX41 U13038 ( .I0(ram[8794]), .I1(ram[8786]), .I2(ram[8778]), .I3(
        ram[8770]), .S0(n27123), .S1(n26648), .ZN(n22346) );
  MUX41 U13039 ( .I0(ram[4315]), .I1(ram[4307]), .I2(ram[4299]), .I3(
        ram[4291]), .S0(n27152), .S1(n26677), .ZN(n22844) );
  MUX41 U13040 ( .I0(ram[4187]), .I1(ram[4179]), .I2(ram[4171]), .I3(
        ram[4163]), .S0(n27152), .S1(n26677), .ZN(n22839) );
  MUX41 U13041 ( .I0(ram[5083]), .I1(ram[5075]), .I2(ram[5067]), .I3(
        ram[5059]), .S0(n27154), .S1(n26679), .ZN(n22874) );
  MUX41 U13042 ( .I0(ram[4827]), .I1(ram[4819]), .I2(ram[4811]), .I3(
        ram[4803]), .S0(n27153), .S1(n26678), .ZN(n22864) );
  MUX41 U13043 ( .I0(ram[4699]), .I1(ram[4691]), .I2(ram[4683]), .I3(
        ram[4675]), .S0(n27153), .S1(n26678), .ZN(n22859) );
  MUX41 U13044 ( .I0(ram[10843]), .I1(ram[10835]), .I2(ram[10827]), .I3(
        ram[10819]), .S0(n27168), .S1(n26693), .ZN(n23115) );
  MUX41 U13045 ( .I0(ram[8923]), .I1(ram[8915]), .I2(ram[8907]), .I3(
        ram[8899]), .S0(n27163), .S1(n26688), .ZN(n23035) );
  MUX41 U13046 ( .I0(ram[8795]), .I1(ram[8787]), .I2(ram[8779]), .I3(
        ram[8771]), .S0(n27163), .S1(n26688), .ZN(n23030) );
  MUX41 U13047 ( .I0(ram[4316]), .I1(ram[4308]), .I2(ram[4300]), .I3(
        ram[4292]), .S0(n27191), .S1(n26716), .ZN(n23528) );
  MUX41 U13048 ( .I0(ram[4188]), .I1(ram[4180]), .I2(ram[4172]), .I3(
        ram[4164]), .S0(n27191), .S1(n26716), .ZN(n23523) );
  MUX41 U13049 ( .I0(ram[5084]), .I1(ram[5076]), .I2(ram[5068]), .I3(
        ram[5060]), .S0(n27193), .S1(n26718), .ZN(n23558) );
  MUX41 U13050 ( .I0(ram[4828]), .I1(ram[4820]), .I2(ram[4812]), .I3(
        ram[4804]), .S0(n27193), .S1(n26718), .ZN(n23548) );
  MUX41 U13051 ( .I0(ram[4700]), .I1(ram[4692]), .I2(ram[4684]), .I3(
        ram[4676]), .S0(n27192), .S1(n26717), .ZN(n23543) );
  MUX41 U13052 ( .I0(ram[10844]), .I1(ram[10836]), .I2(ram[10828]), .I3(
        ram[10820]), .S0(n27207), .S1(n26732), .ZN(n23799) );
  MUX41 U13053 ( .I0(ram[8924]), .I1(ram[8916]), .I2(ram[8908]), .I3(
        ram[8900]), .S0(n27202), .S1(n26727), .ZN(n23719) );
  MUX41 U13054 ( .I0(ram[8796]), .I1(ram[8788]), .I2(ram[8780]), .I3(
        ram[8772]), .S0(n27202), .S1(n26727), .ZN(n23714) );
  MUX41 U13055 ( .I0(ram[4317]), .I1(ram[4309]), .I2(ram[4301]), .I3(
        ram[4293]), .S0(n27231), .S1(n26756), .ZN(n24212) );
  MUX41 U13056 ( .I0(ram[4189]), .I1(ram[4181]), .I2(ram[4173]), .I3(
        ram[4165]), .S0(n27230), .S1(n26755), .ZN(n24207) );
  MUX41 U13057 ( .I0(ram[5085]), .I1(ram[5077]), .I2(ram[5069]), .I3(
        ram[5061]), .S0(n27233), .S1(n26758), .ZN(n24242) );
  MUX41 U13058 ( .I0(ram[4829]), .I1(ram[4821]), .I2(ram[4813]), .I3(
        ram[4805]), .S0(n27232), .S1(n26757), .ZN(n24232) );
  MUX41 U13059 ( .I0(ram[4701]), .I1(ram[4693]), .I2(ram[4685]), .I3(
        ram[4677]), .S0(n27232), .S1(n26757), .ZN(n24227) );
  MUX41 U13060 ( .I0(ram[10845]), .I1(ram[10837]), .I2(ram[10829]), .I3(
        ram[10821]), .S0(n27246), .S1(n26771), .ZN(n24483) );
  MUX41 U13061 ( .I0(ram[8925]), .I1(ram[8917]), .I2(ram[8909]), .I3(
        ram[8901]), .S0(n27242), .S1(n26767), .ZN(n24403) );
  MUX41 U13062 ( .I0(ram[8797]), .I1(ram[8789]), .I2(ram[8781]), .I3(
        ram[8773]), .S0(n27241), .S1(n26766), .ZN(n24398) );
  MUX41 U13063 ( .I0(ram[4318]), .I1(ram[4310]), .I2(ram[4302]), .I3(
        ram[4294]), .S0(n27270), .S1(n26795), .ZN(n24896) );
  MUX41 U13064 ( .I0(ram[4190]), .I1(ram[4182]), .I2(ram[4174]), .I3(
        ram[4166]), .S0(n27270), .S1(n26795), .ZN(n24891) );
  MUX41 U13065 ( .I0(ram[5086]), .I1(ram[5078]), .I2(ram[5070]), .I3(
        ram[5062]), .S0(n27272), .S1(n26797), .ZN(n24926) );
  MUX41 U13066 ( .I0(ram[4830]), .I1(ram[4822]), .I2(ram[4814]), .I3(
        ram[4806]), .S0(n27271), .S1(n26796), .ZN(n24916) );
  MUX41 U13067 ( .I0(ram[4702]), .I1(ram[4694]), .I2(ram[4686]), .I3(
        ram[4678]), .S0(n27271), .S1(n26796), .ZN(n24911) );
  MUX41 U13068 ( .I0(ram[10846]), .I1(ram[10838]), .I2(ram[10830]), .I3(
        ram[10822]), .S0(n27286), .S1(n26811), .ZN(n25167) );
  MUX41 U13069 ( .I0(ram[8926]), .I1(ram[8918]), .I2(ram[8910]), .I3(
        ram[8902]), .S0(n27281), .S1(n26806), .ZN(n25087) );
  MUX41 U13070 ( .I0(ram[8798]), .I1(ram[8790]), .I2(ram[8782]), .I3(
        ram[8774]), .S0(n27281), .S1(n26806), .ZN(n25082) );
  MUX41 U13071 ( .I0(ram[4319]), .I1(ram[4311]), .I2(ram[4303]), .I3(
        ram[4295]), .S0(n27309), .S1(n26834), .ZN(n25580) );
  MUX41 U13072 ( .I0(ram[4191]), .I1(ram[4183]), .I2(ram[4175]), .I3(
        ram[4167]), .S0(n27309), .S1(n26834), .ZN(n25575) );
  MUX41 U13073 ( .I0(ram[5087]), .I1(ram[5079]), .I2(ram[5071]), .I3(
        ram[5063]), .S0(n27311), .S1(n26836), .ZN(n25610) );
  MUX41 U13074 ( .I0(ram[4831]), .I1(ram[4823]), .I2(ram[4815]), .I3(
        ram[4807]), .S0(n27311), .S1(n26836), .ZN(n25600) );
  MUX41 U13075 ( .I0(ram[4703]), .I1(ram[4695]), .I2(ram[4687]), .I3(
        ram[4679]), .S0(n27310), .S1(n26835), .ZN(n25595) );
  MUX41 U13076 ( .I0(ram[10847]), .I1(ram[10839]), .I2(ram[10831]), .I3(
        ram[10823]), .S0(n27325), .S1(n26850), .ZN(n25851) );
  MUX41 U13077 ( .I0(ram[8927]), .I1(ram[8919]), .I2(ram[8911]), .I3(
        ram[8903]), .S0(n27321), .S1(n26846), .ZN(n25771) );
  MUX41 U13078 ( .I0(ram[8799]), .I1(ram[8791]), .I2(ram[8783]), .I3(
        ram[8775]), .S0(n27320), .S1(n26845), .ZN(n25766) );
  MUX41 U13079 ( .I0(ram[2296]), .I1(ram[2288]), .I2(ram[2280]), .I3(
        ram[2272]), .S0(n27029), .S1(n26554), .ZN(n20704) );
  MUX41 U13080 ( .I0(ram[2168]), .I1(ram[2160]), .I2(ram[2152]), .I3(
        ram[2144]), .S0(n27029), .S1(n26554), .ZN(n20699) );
  MUX41 U13081 ( .I0(ram[3064]), .I1(ram[3056]), .I2(ram[3048]), .I3(
        ram[3040]), .S0(n27031), .S1(n26556), .ZN(n20734) );
  MUX41 U13082 ( .I0(ram[2808]), .I1(ram[2800]), .I2(ram[2792]), .I3(
        ram[2784]), .S0(n27030), .S1(n26555), .ZN(n20724) );
  MUX41 U13083 ( .I0(ram[2680]), .I1(ram[2672]), .I2(ram[2664]), .I3(
        ram[2656]), .S0(n27030), .S1(n26555), .ZN(n20719) );
  MUX41 U13084 ( .I0(ram[504]), .I1(ram[496]), .I2(ram[488]), .I3(
        ram[480]), .S0(n27025), .S1(n26550), .ZN(n20629) );
  MUX41 U13085 ( .I0(ram[248]), .I1(ram[240]), .I2(ram[232]), .I3(
        ram[224]), .S0(n27024), .S1(n26549), .ZN(n3453) );
  MUX41 U13086 ( .I0(ram[120]), .I1(ram[112]), .I2(ram[104]), .I3(ram[96]), .S0(n27024), .S1(n26549), .ZN(n2807) );
  MUX41 U13087 ( .I0(ram[2297]), .I1(ram[2289]), .I2(ram[2281]), .I3(
        ram[2273]), .S0(n27068), .S1(n26593), .ZN(n21388) );
  MUX41 U13088 ( .I0(ram[2169]), .I1(ram[2161]), .I2(ram[2153]), .I3(
        ram[2145]), .S0(n27068), .S1(n26593), .ZN(n21383) );
  MUX41 U13089 ( .I0(ram[3065]), .I1(ram[3057]), .I2(ram[3049]), .I3(
        ram[3041]), .S0(n27070), .S1(n26595), .ZN(n21418) );
  MUX41 U13090 ( .I0(ram[2809]), .I1(ram[2801]), .I2(ram[2793]), .I3(
        ram[2785]), .S0(n27070), .S1(n26595), .ZN(n21408) );
  MUX41 U13091 ( .I0(ram[2681]), .I1(ram[2673]), .I2(ram[2665]), .I3(
        ram[2657]), .S0(n27069), .S1(n26594), .ZN(n21403) );
  MUX41 U13092 ( .I0(ram[249]), .I1(ram[241]), .I2(ram[233]), .I3(
        ram[225]), .S0(n27063), .S1(n26588), .ZN(n21303) );
  MUX41 U13093 ( .I0(ram[121]), .I1(ram[113]), .I2(ram[105]), .I3(ram[97]), .S0(n27063), .S1(n26588), .ZN(n21298) );
  MUX41 U13094 ( .I0(ram[2298]), .I1(ram[2290]), .I2(ram[2282]), .I3(
        ram[2274]), .S0(n27108), .S1(n26633), .ZN(n22072) );
  MUX41 U13095 ( .I0(ram[2170]), .I1(ram[2162]), .I2(ram[2154]), .I3(
        ram[2146]), .S0(n27107), .S1(n26632), .ZN(n22067) );
  MUX41 U13096 ( .I0(ram[3066]), .I1(ram[3058]), .I2(ram[3050]), .I3(
        ram[3042]), .S0(n27110), .S1(n26635), .ZN(n22102) );
  MUX41 U13097 ( .I0(ram[2810]), .I1(ram[2802]), .I2(ram[2794]), .I3(
        ram[2786]), .S0(n27109), .S1(n26634), .ZN(n22092) );
  MUX41 U13098 ( .I0(ram[2682]), .I1(ram[2674]), .I2(ram[2666]), .I3(
        ram[2658]), .S0(n27109), .S1(n26634), .ZN(n22087) );
  MUX41 U13099 ( .I0(ram[250]), .I1(ram[242]), .I2(ram[234]), .I3(
        ram[226]), .S0(n27103), .S1(n26628), .ZN(n21987) );
  MUX41 U13100 ( .I0(ram[122]), .I1(ram[114]), .I2(ram[106]), .I3(ram[98]), .S0(n27102), .S1(n26627), .ZN(n21982) );
  MUX41 U13101 ( .I0(ram[2299]), .I1(ram[2291]), .I2(ram[2283]), .I3(
        ram[2275]), .S0(n27147), .S1(n26672), .ZN(n22756) );
  MUX41 U13102 ( .I0(ram[2171]), .I1(ram[2163]), .I2(ram[2155]), .I3(
        ram[2147]), .S0(n27147), .S1(n26672), .ZN(n22751) );
  MUX41 U13103 ( .I0(ram[3067]), .I1(ram[3059]), .I2(ram[3051]), .I3(
        ram[3043]), .S0(n27149), .S1(n26674), .ZN(n22786) );
  MUX41 U13104 ( .I0(ram[2811]), .I1(ram[2803]), .I2(ram[2795]), .I3(
        ram[2787]), .S0(n27148), .S1(n26673), .ZN(n22776) );
  MUX41 U13105 ( .I0(ram[2683]), .I1(ram[2675]), .I2(ram[2667]), .I3(
        ram[2659]), .S0(n27148), .S1(n26673), .ZN(n22771) );
  MUX41 U13106 ( .I0(ram[251]), .I1(ram[243]), .I2(ram[235]), .I3(
        ram[227]), .S0(n27142), .S1(n26667), .ZN(n22671) );
  MUX41 U13107 ( .I0(ram[123]), .I1(ram[115]), .I2(ram[107]), .I3(ram[99]), .S0(n27142), .S1(n26667), .ZN(n22666) );
  MUX41 U13108 ( .I0(ram[2300]), .I1(ram[2292]), .I2(ram[2284]), .I3(
        ram[2276]), .S0(n27186), .S1(n26711), .ZN(n23440) );
  MUX41 U13109 ( .I0(ram[2172]), .I1(ram[2164]), .I2(ram[2156]), .I3(
        ram[2148]), .S0(n27186), .S1(n26711), .ZN(n23435) );
  MUX41 U13110 ( .I0(ram[3068]), .I1(ram[3060]), .I2(ram[3052]), .I3(
        ram[3044]), .S0(n27188), .S1(n26713), .ZN(n23470) );
  MUX41 U13111 ( .I0(ram[2812]), .I1(ram[2804]), .I2(ram[2796]), .I3(
        ram[2788]), .S0(n27188), .S1(n26713), .ZN(n23460) );
  MUX41 U13112 ( .I0(ram[2684]), .I1(ram[2676]), .I2(ram[2668]), .I3(
        ram[2660]), .S0(n27187), .S1(n26712), .ZN(n23455) );
  MUX41 U13113 ( .I0(ram[252]), .I1(ram[244]), .I2(ram[236]), .I3(
        ram[228]), .S0(n27182), .S1(n26707), .ZN(n23355) );
  MUX41 U13114 ( .I0(ram[124]), .I1(ram[116]), .I2(ram[108]), .I3(
        ram[100]), .S0(n27181), .S1(n26706), .ZN(n23350) );
  MUX41 U13115 ( .I0(ram[2301]), .I1(ram[2293]), .I2(ram[2285]), .I3(
        ram[2277]), .S0(n27226), .S1(n26751), .ZN(n24124) );
  MUX41 U13116 ( .I0(ram[2173]), .I1(ram[2165]), .I2(ram[2157]), .I3(
        ram[2149]), .S0(n27226), .S1(n26751), .ZN(n24119) );
  MUX41 U13117 ( .I0(ram[3069]), .I1(ram[3061]), .I2(ram[3053]), .I3(
        ram[3045]), .S0(n27228), .S1(n26753), .ZN(n24154) );
  MUX41 U13118 ( .I0(ram[2813]), .I1(ram[2805]), .I2(ram[2797]), .I3(
        ram[2789]), .S0(n27227), .S1(n26752), .ZN(n24144) );
  MUX41 U13119 ( .I0(ram[2685]), .I1(ram[2677]), .I2(ram[2669]), .I3(
        ram[2661]), .S0(n27227), .S1(n26752), .ZN(n24139) );
  MUX41 U13120 ( .I0(ram[253]), .I1(ram[245]), .I2(ram[237]), .I3(
        ram[229]), .S0(n27221), .S1(n26746), .ZN(n24039) );
  MUX41 U13121 ( .I0(ram[125]), .I1(ram[117]), .I2(ram[109]), .I3(
        ram[101]), .S0(n27221), .S1(n26746), .ZN(n24034) );
  MUX41 U13122 ( .I0(ram[2302]), .I1(ram[2294]), .I2(ram[2286]), .I3(
        ram[2278]), .S0(n27265), .S1(n26790), .ZN(n24808) );
  MUX41 U13123 ( .I0(ram[2174]), .I1(ram[2166]), .I2(ram[2158]), .I3(
        ram[2150]), .S0(n27265), .S1(n26790), .ZN(n24803) );
  MUX41 U13124 ( .I0(ram[3070]), .I1(ram[3062]), .I2(ram[3054]), .I3(
        ram[3046]), .S0(n27267), .S1(n26792), .ZN(n24838) );
  MUX41 U13125 ( .I0(ram[2814]), .I1(ram[2806]), .I2(ram[2798]), .I3(
        ram[2790]), .S0(n27266), .S1(n26791), .ZN(n24828) );
  MUX41 U13126 ( .I0(ram[2686]), .I1(ram[2678]), .I2(ram[2670]), .I3(
        ram[2662]), .S0(n27266), .S1(n26791), .ZN(n24823) );
  MUX41 U13127 ( .I0(ram[254]), .I1(ram[246]), .I2(ram[238]), .I3(
        ram[230]), .S0(n27260), .S1(n26785), .ZN(n24723) );
  MUX41 U13128 ( .I0(ram[126]), .I1(ram[118]), .I2(ram[110]), .I3(
        ram[102]), .S0(n27260), .S1(n26785), .ZN(n24718) );
  MUX41 U13129 ( .I0(ram[2303]), .I1(ram[2295]), .I2(ram[2287]), .I3(
        ram[2279]), .S0(n27305), .S1(n26830), .ZN(n25492) );
  MUX41 U13130 ( .I0(ram[2175]), .I1(ram[2167]), .I2(ram[2159]), .I3(
        ram[2151]), .S0(n27304), .S1(n26829), .ZN(n25487) );
  MUX41 U13131 ( .I0(ram[3071]), .I1(ram[3063]), .I2(ram[3055]), .I3(
        ram[3047]), .S0(n27306), .S1(n26831), .ZN(n25522) );
  MUX41 U13132 ( .I0(ram[2815]), .I1(ram[2807]), .I2(ram[2799]), .I3(
        ram[2791]), .S0(n27306), .S1(n26831), .ZN(n25512) );
  MUX41 U13133 ( .I0(ram[2687]), .I1(ram[2679]), .I2(ram[2671]), .I3(
        ram[2663]), .S0(n27306), .S1(n26831), .ZN(n25507) );
  MUX41 U13134 ( .I0(ram[255]), .I1(ram[247]), .I2(ram[239]), .I3(
        ram[231]), .S0(n27300), .S1(n26825), .ZN(n25407) );
  MUX41 U13135 ( .I0(ram[127]), .I1(ram[119]), .I2(ram[111]), .I3(
        ram[103]), .S0(n27299), .S1(n26824), .ZN(n25402) );
  MUX41 U13136 ( .I0(n20820), .I1(n20821), .I2(n20822), .I3(n20823), .S0(
        n26197), .S1(n26315), .ZN(n20819) );
  MUX41 U13137 ( .I0(ram[5048]), .I1(ram[5040]), .I2(ram[5032]), .I3(
        ram[5024]), .S0(n27036), .S1(n26561), .ZN(n20821) );
  MUX41 U13138 ( .I0(ram[5016]), .I1(ram[5008]), .I2(ram[5000]), .I3(
        ram[4992]), .S0(n27035), .S1(n26560), .ZN(n20823) );
  MUX41 U13139 ( .I0(ram[5112]), .I1(ram[5104]), .I2(ram[5096]), .I3(
        ram[5088]), .S0(n27036), .S1(n26561), .ZN(n20820) );
  MUX41 U13140 ( .I0(n21504), .I1(n21505), .I2(n21506), .I3(n21507), .S0(
        n26207), .S1(n26325), .ZN(n21503) );
  MUX41 U13141 ( .I0(ram[5049]), .I1(ram[5041]), .I2(ram[5033]), .I3(
        ram[5025]), .S0(n27075), .S1(n26600), .ZN(n21505) );
  MUX41 U13142 ( .I0(ram[5017]), .I1(ram[5009]), .I2(ram[5001]), .I3(
        ram[4993]), .S0(n27075), .S1(n26600), .ZN(n21507) );
  MUX41 U13143 ( .I0(ram[5113]), .I1(ram[5105]), .I2(ram[5097]), .I3(
        ram[5089]), .S0(n27075), .S1(n26600), .ZN(n21504) );
  MUX41 U13144 ( .I0(n22188), .I1(n22189), .I2(n22190), .I3(n22191), .S0(
        n26216), .S1(n26334), .ZN(n22187) );
  MUX41 U13145 ( .I0(ram[5050]), .I1(ram[5042]), .I2(ram[5034]), .I3(
        ram[5026]), .S0(n27114), .S1(n26639), .ZN(n22189) );
  MUX41 U13146 ( .I0(ram[5018]), .I1(ram[5010]), .I2(ram[5002]), .I3(
        ram[4994]), .S0(n27114), .S1(n26639), .ZN(n22191) );
  MUX41 U13147 ( .I0(ram[5114]), .I1(ram[5106]), .I2(ram[5098]), .I3(
        ram[5090]), .S0(n27114), .S1(n26639), .ZN(n22188) );
  MUX41 U13148 ( .I0(n22872), .I1(n22873), .I2(n22874), .I3(n22875), .S0(
        n26226), .S1(n26344), .ZN(n22871) );
  MUX41 U13149 ( .I0(ram[5051]), .I1(ram[5043]), .I2(ram[5035]), .I3(
        ram[5027]), .S0(n27154), .S1(n26679), .ZN(n22873) );
  MUX41 U13150 ( .I0(ram[5019]), .I1(ram[5011]), .I2(ram[5003]), .I3(
        ram[4995]), .S0(n27154), .S1(n26679), .ZN(n22875) );
  MUX41 U13151 ( .I0(ram[5115]), .I1(ram[5107]), .I2(ram[5099]), .I3(
        ram[5091]), .S0(n27154), .S1(n26679), .ZN(n22872) );
  MUX41 U13152 ( .I0(n23556), .I1(n23557), .I2(n23558), .I3(n23559), .S0(
        n26236), .S1(n26354), .ZN(n23555) );
  MUX41 U13153 ( .I0(ram[5052]), .I1(ram[5044]), .I2(ram[5036]), .I3(
        ram[5028]), .S0(n27193), .S1(n26718), .ZN(n23557) );
  MUX41 U13154 ( .I0(ram[5020]), .I1(ram[5012]), .I2(ram[5004]), .I3(
        ram[4996]), .S0(n27193), .S1(n26718), .ZN(n23559) );
  MUX41 U13155 ( .I0(ram[5116]), .I1(ram[5108]), .I2(ram[5100]), .I3(
        ram[5092]), .S0(n27193), .S1(n26718), .ZN(n23556) );
  MUX41 U13156 ( .I0(n24240), .I1(n24241), .I2(n24242), .I3(n24243), .S0(
        n26246), .S1(n26364), .ZN(n24239) );
  MUX41 U13157 ( .I0(ram[5053]), .I1(ram[5045]), .I2(ram[5037]), .I3(
        ram[5029]), .S0(n27232), .S1(n26757), .ZN(n24241) );
  MUX41 U13158 ( .I0(ram[5021]), .I1(ram[5013]), .I2(ram[5005]), .I3(
        ram[4997]), .S0(n27232), .S1(n26757), .ZN(n24243) );
  MUX41 U13159 ( .I0(ram[5117]), .I1(ram[5109]), .I2(ram[5101]), .I3(
        ram[5093]), .S0(n27233), .S1(n26758), .ZN(n24240) );
  MUX41 U13160 ( .I0(n24924), .I1(n24925), .I2(n24926), .I3(n24927), .S0(
        n26256), .S1(n26374), .ZN(n24923) );
  MUX41 U13161 ( .I0(ram[5054]), .I1(ram[5046]), .I2(ram[5038]), .I3(
        ram[5030]), .S0(n27272), .S1(n26797), .ZN(n24925) );
  MUX41 U13162 ( .I0(ram[5022]), .I1(ram[5014]), .I2(ram[5006]), .I3(
        ram[4998]), .S0(n27272), .S1(n26797), .ZN(n24927) );
  MUX41 U13163 ( .I0(ram[5118]), .I1(ram[5110]), .I2(ram[5102]), .I3(
        ram[5094]), .S0(n27272), .S1(n26797), .ZN(n24924) );
  MUX41 U13164 ( .I0(n25608), .I1(n25609), .I2(n25610), .I3(n25611), .S0(
        n26266), .S1(n26384), .ZN(n25607) );
  MUX41 U13165 ( .I0(ram[5055]), .I1(ram[5047]), .I2(ram[5039]), .I3(
        ram[5031]), .S0(n27311), .S1(n26836), .ZN(n25609) );
  MUX41 U13166 ( .I0(ram[5023]), .I1(ram[5015]), .I2(ram[5007]), .I3(
        ram[4999]), .S0(n27311), .S1(n26836), .ZN(n25611) );
  MUX41 U13167 ( .I0(ram[5119]), .I1(ram[5111]), .I2(ram[5103]), .I3(
        ram[5095]), .S0(n27311), .S1(n26836), .ZN(n25608) );
  BUF U13168 ( .I(raddr[3]), .Z(n29318) );
  BUF U13169 ( .I(raddr[2]), .Z(n29317) );
  MOAI22 U13170 ( .A1(n13), .A2(n29088), .B1(ram[0]), .B2(n15), .ZN(n4241) );
  MOAI22 U13171 ( .A1(n13), .A2(n28853), .B1(ram[1]), .B2(n15), .ZN(n4242) );
  MOAI22 U13172 ( .A1(n13), .A2(n28618), .B1(ram[2]), .B2(n15), .ZN(n4243) );
  MOAI22 U13173 ( .A1(n13), .A2(n28383), .B1(ram[3]), .B2(n15), .ZN(n4244) );
  MOAI22 U13174 ( .A1(n13), .A2(n28148), .B1(ram[4]), .B2(n15), .ZN(n4245) );
  MOAI22 U13175 ( .A1(n13), .A2(n27913), .B1(ram[5]), .B2(n15), .ZN(n4246) );
  MOAI22 U13176 ( .A1(n13), .A2(n27678), .B1(ram[6]), .B2(n15), .ZN(n4247) );
  MOAI22 U13177 ( .A1(n13), .A2(n27443), .B1(ram[7]), .B2(n15), .ZN(n4248) );
  MOAI22 U13178 ( .A1(n29088), .A2(n25), .B1(ram[8]), .B2(n26), .ZN(n4249) );
  MOAI22 U13179 ( .A1(n28853), .A2(n25), .B1(ram[9]), .B2(n26), .ZN(n4250) );
  MOAI22 U13180 ( .A1(n28618), .A2(n25), .B1(ram[10]), .B2(n26), .ZN(
        n4251) );
  MOAI22 U13181 ( .A1(n28383), .A2(n25), .B1(ram[11]), .B2(n26), .ZN(
        n4252) );
  MOAI22 U13182 ( .A1(n28148), .A2(n25), .B1(ram[12]), .B2(n26), .ZN(
        n4253) );
  MOAI22 U13183 ( .A1(n27913), .A2(n25), .B1(ram[13]), .B2(n26), .ZN(
        n4254) );
  MOAI22 U13184 ( .A1(n27678), .A2(n25), .B1(ram[14]), .B2(n26), .ZN(
        n4255) );
  MOAI22 U13185 ( .A1(n27443), .A2(n25), .B1(ram[15]), .B2(n26), .ZN(
        n4256) );
  MOAI22 U13186 ( .A1(n29088), .A2(n28), .B1(ram[16]), .B2(n29), .ZN(
        n4257) );
  MOAI22 U13187 ( .A1(n28853), .A2(n28), .B1(ram[17]), .B2(n29), .ZN(
        n4258) );
  MOAI22 U13188 ( .A1(n28618), .A2(n28), .B1(ram[18]), .B2(n29), .ZN(
        n4259) );
  MOAI22 U13189 ( .A1(n28383), .A2(n28), .B1(ram[19]), .B2(n29), .ZN(
        n4260) );
  MOAI22 U13190 ( .A1(n28148), .A2(n28), .B1(ram[20]), .B2(n29), .ZN(
        n4261) );
  MOAI22 U13191 ( .A1(n27913), .A2(n28), .B1(ram[21]), .B2(n29), .ZN(
        n4262) );
  MOAI22 U13192 ( .A1(n27678), .A2(n28), .B1(ram[22]), .B2(n29), .ZN(
        n4263) );
  MOAI22 U13193 ( .A1(n27443), .A2(n28), .B1(ram[23]), .B2(n29), .ZN(
        n4264) );
  MOAI22 U13194 ( .A1(n29088), .A2(n31), .B1(ram[24]), .B2(n32), .ZN(
        n4265) );
  MOAI22 U13195 ( .A1(n28853), .A2(n31), .B1(ram[25]), .B2(n32), .ZN(
        n4266) );
  MOAI22 U13196 ( .A1(n28618), .A2(n31), .B1(ram[26]), .B2(n32), .ZN(
        n4267) );
  MOAI22 U13197 ( .A1(n28383), .A2(n31), .B1(ram[27]), .B2(n32), .ZN(
        n4268) );
  MOAI22 U13198 ( .A1(n28148), .A2(n31), .B1(ram[28]), .B2(n32), .ZN(
        n4269) );
  MOAI22 U13199 ( .A1(n27913), .A2(n31), .B1(ram[29]), .B2(n32), .ZN(
        n4270) );
  MOAI22 U13200 ( .A1(n27678), .A2(n31), .B1(ram[30]), .B2(n32), .ZN(
        n4271) );
  MOAI22 U13201 ( .A1(n27443), .A2(n31), .B1(ram[31]), .B2(n32), .ZN(
        n4272) );
  MOAI22 U13202 ( .A1(n29088), .A2(n34), .B1(ram[32]), .B2(n35), .ZN(
        n4273) );
  MOAI22 U13203 ( .A1(n28853), .A2(n34), .B1(ram[33]), .B2(n35), .ZN(
        n4274) );
  MOAI22 U13204 ( .A1(n28618), .A2(n34), .B1(ram[34]), .B2(n35), .ZN(
        n4275) );
  MOAI22 U13205 ( .A1(n28383), .A2(n34), .B1(ram[35]), .B2(n35), .ZN(
        n4276) );
  MOAI22 U13206 ( .A1(n28148), .A2(n34), .B1(ram[36]), .B2(n35), .ZN(
        n4277) );
  MOAI22 U13207 ( .A1(n27913), .A2(n34), .B1(ram[37]), .B2(n35), .ZN(
        n4278) );
  MOAI22 U13208 ( .A1(n27678), .A2(n34), .B1(ram[38]), .B2(n35), .ZN(
        n4279) );
  MOAI22 U13209 ( .A1(n27443), .A2(n34), .B1(ram[39]), .B2(n35), .ZN(
        n4280) );
  MOAI22 U13210 ( .A1(n29088), .A2(n37), .B1(ram[40]), .B2(n38), .ZN(
        n4281) );
  MOAI22 U13211 ( .A1(n28853), .A2(n37), .B1(ram[41]), .B2(n38), .ZN(
        n4282) );
  MOAI22 U13212 ( .A1(n28618), .A2(n37), .B1(ram[42]), .B2(n38), .ZN(
        n4283) );
  MOAI22 U13213 ( .A1(n28383), .A2(n37), .B1(ram[43]), .B2(n38), .ZN(
        n4284) );
  MOAI22 U13214 ( .A1(n28148), .A2(n37), .B1(ram[44]), .B2(n38), .ZN(
        n4285) );
  MOAI22 U13215 ( .A1(n27913), .A2(n37), .B1(ram[45]), .B2(n38), .ZN(
        n4286) );
  MOAI22 U13216 ( .A1(n27678), .A2(n37), .B1(ram[46]), .B2(n38), .ZN(
        n4287) );
  MOAI22 U13217 ( .A1(n27443), .A2(n37), .B1(ram[47]), .B2(n38), .ZN(
        n4288) );
  MOAI22 U13218 ( .A1(n29088), .A2(n40), .B1(ram[48]), .B2(n41), .ZN(
        n4289) );
  MOAI22 U13219 ( .A1(n28853), .A2(n40), .B1(ram[49]), .B2(n41), .ZN(
        n4290) );
  MOAI22 U13220 ( .A1(n28618), .A2(n40), .B1(ram[50]), .B2(n41), .ZN(
        n4291) );
  MOAI22 U13221 ( .A1(n28383), .A2(n40), .B1(ram[51]), .B2(n41), .ZN(
        n4292) );
  MOAI22 U13222 ( .A1(n28148), .A2(n40), .B1(ram[52]), .B2(n41), .ZN(
        n4293) );
  MOAI22 U13223 ( .A1(n27913), .A2(n40), .B1(ram[53]), .B2(n41), .ZN(
        n4294) );
  MOAI22 U13224 ( .A1(n27678), .A2(n40), .B1(ram[54]), .B2(n41), .ZN(
        n4295) );
  MOAI22 U13225 ( .A1(n27443), .A2(n40), .B1(ram[55]), .B2(n41), .ZN(
        n4296) );
  MOAI22 U13226 ( .A1(n29088), .A2(n43), .B1(ram[56]), .B2(n44), .ZN(
        n4297) );
  MOAI22 U13227 ( .A1(n28853), .A2(n43), .B1(ram[57]), .B2(n44), .ZN(
        n4298) );
  MOAI22 U13228 ( .A1(n28618), .A2(n43), .B1(ram[58]), .B2(n44), .ZN(
        n4299) );
  MOAI22 U13229 ( .A1(n28383), .A2(n43), .B1(ram[59]), .B2(n44), .ZN(
        n4300) );
  MOAI22 U13230 ( .A1(n28148), .A2(n43), .B1(ram[60]), .B2(n44), .ZN(
        n4301) );
  MOAI22 U13231 ( .A1(n27913), .A2(n43), .B1(ram[61]), .B2(n44), .ZN(
        n4302) );
  MOAI22 U13232 ( .A1(n27678), .A2(n43), .B1(ram[62]), .B2(n44), .ZN(
        n4303) );
  MOAI22 U13233 ( .A1(n27443), .A2(n43), .B1(ram[63]), .B2(n44), .ZN(
        n4304) );
  MOAI22 U13234 ( .A1(n29088), .A2(n46), .B1(ram[64]), .B2(n47), .ZN(
        n4305) );
  MOAI22 U13235 ( .A1(n28853), .A2(n46), .B1(ram[65]), .B2(n47), .ZN(
        n4306) );
  MOAI22 U13236 ( .A1(n28618), .A2(n46), .B1(ram[66]), .B2(n47), .ZN(
        n4307) );
  MOAI22 U13237 ( .A1(n28383), .A2(n46), .B1(ram[67]), .B2(n47), .ZN(
        n4308) );
  MOAI22 U13238 ( .A1(n28148), .A2(n46), .B1(ram[68]), .B2(n47), .ZN(
        n4309) );
  MOAI22 U13239 ( .A1(n27913), .A2(n46), .B1(ram[69]), .B2(n47), .ZN(
        n4310) );
  MOAI22 U13240 ( .A1(n27678), .A2(n46), .B1(ram[70]), .B2(n47), .ZN(
        n4311) );
  MOAI22 U13241 ( .A1(n27443), .A2(n46), .B1(ram[71]), .B2(n47), .ZN(
        n4312) );
  MOAI22 U13242 ( .A1(n29088), .A2(n49), .B1(ram[72]), .B2(n50), .ZN(
        n4313) );
  MOAI22 U13243 ( .A1(n28853), .A2(n49), .B1(ram[73]), .B2(n50), .ZN(
        n4314) );
  MOAI22 U13244 ( .A1(n28618), .A2(n49), .B1(ram[74]), .B2(n50), .ZN(
        n4315) );
  MOAI22 U13245 ( .A1(n28383), .A2(n49), .B1(ram[75]), .B2(n50), .ZN(
        n4316) );
  MOAI22 U13246 ( .A1(n28148), .A2(n49), .B1(ram[76]), .B2(n50), .ZN(
        n4317) );
  MOAI22 U13247 ( .A1(n27913), .A2(n49), .B1(ram[77]), .B2(n50), .ZN(
        n4318) );
  MOAI22 U13248 ( .A1(n27678), .A2(n49), .B1(ram[78]), .B2(n50), .ZN(
        n4319) );
  MOAI22 U13249 ( .A1(n27443), .A2(n49), .B1(ram[79]), .B2(n50), .ZN(
        n4320) );
  MOAI22 U13250 ( .A1(n29088), .A2(n52), .B1(ram[80]), .B2(n53), .ZN(
        n4321) );
  MOAI22 U13251 ( .A1(n28853), .A2(n52), .B1(ram[81]), .B2(n53), .ZN(
        n4322) );
  MOAI22 U13252 ( .A1(n28618), .A2(n52), .B1(ram[82]), .B2(n53), .ZN(
        n4323) );
  MOAI22 U13253 ( .A1(n28383), .A2(n52), .B1(ram[83]), .B2(n53), .ZN(
        n4324) );
  MOAI22 U13254 ( .A1(n28148), .A2(n52), .B1(ram[84]), .B2(n53), .ZN(
        n4325) );
  MOAI22 U13255 ( .A1(n27913), .A2(n52), .B1(ram[85]), .B2(n53), .ZN(
        n4326) );
  MOAI22 U13256 ( .A1(n27678), .A2(n52), .B1(ram[86]), .B2(n53), .ZN(
        n4327) );
  MOAI22 U13257 ( .A1(n27443), .A2(n52), .B1(ram[87]), .B2(n53), .ZN(
        n4328) );
  MOAI22 U13258 ( .A1(n29088), .A2(n55), .B1(ram[88]), .B2(n56), .ZN(
        n4329) );
  MOAI22 U13259 ( .A1(n28853), .A2(n55), .B1(ram[89]), .B2(n56), .ZN(
        n4330) );
  MOAI22 U13260 ( .A1(n28618), .A2(n55), .B1(ram[90]), .B2(n56), .ZN(
        n4331) );
  MOAI22 U13261 ( .A1(n28383), .A2(n55), .B1(ram[91]), .B2(n56), .ZN(
        n4332) );
  MOAI22 U13262 ( .A1(n28148), .A2(n55), .B1(ram[92]), .B2(n56), .ZN(
        n4333) );
  MOAI22 U13263 ( .A1(n27913), .A2(n55), .B1(ram[93]), .B2(n56), .ZN(
        n4334) );
  MOAI22 U13264 ( .A1(n27678), .A2(n55), .B1(ram[94]), .B2(n56), .ZN(
        n4335) );
  MOAI22 U13265 ( .A1(n27443), .A2(n55), .B1(ram[95]), .B2(n56), .ZN(
        n4336) );
  MOAI22 U13266 ( .A1(n29088), .A2(n58), .B1(ram[96]), .B2(n59), .ZN(
        n4337) );
  MOAI22 U13267 ( .A1(n28853), .A2(n58), .B1(ram[97]), .B2(n59), .ZN(
        n4338) );
  MOAI22 U13268 ( .A1(n28618), .A2(n58), .B1(ram[98]), .B2(n59), .ZN(
        n4339) );
  MOAI22 U13269 ( .A1(n28383), .A2(n58), .B1(ram[99]), .B2(n59), .ZN(
        n4340) );
  MOAI22 U13270 ( .A1(n28148), .A2(n58), .B1(ram[100]), .B2(n59), .ZN(
        n4341) );
  MOAI22 U13271 ( .A1(n27913), .A2(n58), .B1(ram[101]), .B2(n59), .ZN(
        n4342) );
  MOAI22 U13272 ( .A1(n27678), .A2(n58), .B1(ram[102]), .B2(n59), .ZN(
        n4343) );
  MOAI22 U13273 ( .A1(n27443), .A2(n58), .B1(ram[103]), .B2(n59), .ZN(
        n4344) );
  MOAI22 U13274 ( .A1(n29089), .A2(n61), .B1(ram[104]), .B2(n62), .ZN(
        n4345) );
  MOAI22 U13275 ( .A1(n28854), .A2(n61), .B1(ram[105]), .B2(n62), .ZN(
        n4346) );
  MOAI22 U13276 ( .A1(n28619), .A2(n61), .B1(ram[106]), .B2(n62), .ZN(
        n4347) );
  MOAI22 U13277 ( .A1(n28384), .A2(n61), .B1(ram[107]), .B2(n62), .ZN(
        n4348) );
  MOAI22 U13278 ( .A1(n28149), .A2(n61), .B1(ram[108]), .B2(n62), .ZN(
        n4349) );
  MOAI22 U13279 ( .A1(n27914), .A2(n61), .B1(ram[109]), .B2(n62), .ZN(
        n4350) );
  MOAI22 U13280 ( .A1(n27679), .A2(n61), .B1(ram[110]), .B2(n62), .ZN(
        n4351) );
  MOAI22 U13281 ( .A1(n27444), .A2(n61), .B1(ram[111]), .B2(n62), .ZN(
        n4352) );
  MOAI22 U13282 ( .A1(n29089), .A2(n64), .B1(ram[112]), .B2(n65), .ZN(
        n4353) );
  MOAI22 U13283 ( .A1(n28854), .A2(n64), .B1(ram[113]), .B2(n65), .ZN(
        n4354) );
  MOAI22 U13284 ( .A1(n28619), .A2(n64), .B1(ram[114]), .B2(n65), .ZN(
        n4355) );
  MOAI22 U13285 ( .A1(n28384), .A2(n64), .B1(ram[115]), .B2(n65), .ZN(
        n4356) );
  MOAI22 U13286 ( .A1(n28149), .A2(n64), .B1(ram[116]), .B2(n65), .ZN(
        n4357) );
  MOAI22 U13287 ( .A1(n27914), .A2(n64), .B1(ram[117]), .B2(n65), .ZN(
        n4358) );
  MOAI22 U13288 ( .A1(n27679), .A2(n64), .B1(ram[118]), .B2(n65), .ZN(
        n4359) );
  MOAI22 U13289 ( .A1(n27444), .A2(n64), .B1(ram[119]), .B2(n65), .ZN(
        n4360) );
  MOAI22 U13290 ( .A1(n29089), .A2(n67), .B1(ram[120]), .B2(n68), .ZN(
        n4361) );
  MOAI22 U13291 ( .A1(n28854), .A2(n67), .B1(ram[121]), .B2(n68), .ZN(
        n4362) );
  MOAI22 U13292 ( .A1(n28619), .A2(n67), .B1(ram[122]), .B2(n68), .ZN(
        n4363) );
  MOAI22 U13293 ( .A1(n28384), .A2(n67), .B1(ram[123]), .B2(n68), .ZN(
        n4364) );
  MOAI22 U13294 ( .A1(n28149), .A2(n67), .B1(ram[124]), .B2(n68), .ZN(
        n4365) );
  MOAI22 U13295 ( .A1(n27914), .A2(n67), .B1(ram[125]), .B2(n68), .ZN(
        n4366) );
  MOAI22 U13296 ( .A1(n27679), .A2(n67), .B1(ram[126]), .B2(n68), .ZN(
        n4367) );
  MOAI22 U13297 ( .A1(n27444), .A2(n67), .B1(ram[127]), .B2(n68), .ZN(
        n4368) );
  MOAI22 U13298 ( .A1(n29089), .A2(n70), .B1(ram[128]), .B2(n71), .ZN(
        n4369) );
  MOAI22 U13299 ( .A1(n28854), .A2(n70), .B1(ram[129]), .B2(n71), .ZN(
        n4370) );
  MOAI22 U13300 ( .A1(n28619), .A2(n70), .B1(ram[130]), .B2(n71), .ZN(
        n4371) );
  MOAI22 U13301 ( .A1(n28384), .A2(n70), .B1(ram[131]), .B2(n71), .ZN(
        n4372) );
  MOAI22 U13302 ( .A1(n28149), .A2(n70), .B1(ram[132]), .B2(n71), .ZN(
        n4373) );
  MOAI22 U13303 ( .A1(n27914), .A2(n70), .B1(ram[133]), .B2(n71), .ZN(
        n4374) );
  MOAI22 U13304 ( .A1(n27679), .A2(n70), .B1(ram[134]), .B2(n71), .ZN(
        n4375) );
  MOAI22 U13305 ( .A1(n27444), .A2(n70), .B1(ram[135]), .B2(n71), .ZN(
        n4376) );
  MOAI22 U13306 ( .A1(n29089), .A2(n73), .B1(ram[136]), .B2(n74), .ZN(
        n4377) );
  MOAI22 U13307 ( .A1(n28854), .A2(n73), .B1(ram[137]), .B2(n74), .ZN(
        n4378) );
  MOAI22 U13308 ( .A1(n28619), .A2(n73), .B1(ram[138]), .B2(n74), .ZN(
        n4379) );
  MOAI22 U13309 ( .A1(n28384), .A2(n73), .B1(ram[139]), .B2(n74), .ZN(
        n4380) );
  MOAI22 U13310 ( .A1(n28149), .A2(n73), .B1(ram[140]), .B2(n74), .ZN(
        n4381) );
  MOAI22 U13311 ( .A1(n27914), .A2(n73), .B1(ram[141]), .B2(n74), .ZN(
        n4382) );
  MOAI22 U13312 ( .A1(n27679), .A2(n73), .B1(ram[142]), .B2(n74), .ZN(
        n4383) );
  MOAI22 U13313 ( .A1(n27444), .A2(n73), .B1(ram[143]), .B2(n74), .ZN(
        n4384) );
  MOAI22 U13314 ( .A1(n29089), .A2(n76), .B1(ram[144]), .B2(n77), .ZN(
        n4385) );
  MOAI22 U13315 ( .A1(n28854), .A2(n76), .B1(ram[145]), .B2(n77), .ZN(
        n4386) );
  MOAI22 U13316 ( .A1(n28619), .A2(n76), .B1(ram[146]), .B2(n77), .ZN(
        n4387) );
  MOAI22 U13317 ( .A1(n28384), .A2(n76), .B1(ram[147]), .B2(n77), .ZN(
        n4388) );
  MOAI22 U13318 ( .A1(n28149), .A2(n76), .B1(ram[148]), .B2(n77), .ZN(
        n4389) );
  MOAI22 U13319 ( .A1(n27914), .A2(n76), .B1(ram[149]), .B2(n77), .ZN(
        n4390) );
  MOAI22 U13320 ( .A1(n27679), .A2(n76), .B1(ram[150]), .B2(n77), .ZN(
        n4391) );
  MOAI22 U13321 ( .A1(n27444), .A2(n76), .B1(ram[151]), .B2(n77), .ZN(
        n4392) );
  MOAI22 U13322 ( .A1(n29089), .A2(n79), .B1(ram[152]), .B2(n80), .ZN(
        n4393) );
  MOAI22 U13323 ( .A1(n28854), .A2(n79), .B1(ram[153]), .B2(n80), .ZN(
        n4394) );
  MOAI22 U13324 ( .A1(n28619), .A2(n79), .B1(ram[154]), .B2(n80), .ZN(
        n4395) );
  MOAI22 U13325 ( .A1(n28384), .A2(n79), .B1(ram[155]), .B2(n80), .ZN(
        n4396) );
  MOAI22 U13326 ( .A1(n28149), .A2(n79), .B1(ram[156]), .B2(n80), .ZN(
        n4397) );
  MOAI22 U13327 ( .A1(n27914), .A2(n79), .B1(ram[157]), .B2(n80), .ZN(
        n4398) );
  MOAI22 U13328 ( .A1(n27679), .A2(n79), .B1(ram[158]), .B2(n80), .ZN(
        n4399) );
  MOAI22 U13329 ( .A1(n27444), .A2(n79), .B1(ram[159]), .B2(n80), .ZN(
        n4400) );
  MOAI22 U13330 ( .A1(n29089), .A2(n82), .B1(ram[160]), .B2(n83), .ZN(
        n4401) );
  MOAI22 U13331 ( .A1(n28854), .A2(n82), .B1(ram[161]), .B2(n83), .ZN(
        n4402) );
  MOAI22 U13332 ( .A1(n28619), .A2(n82), .B1(ram[162]), .B2(n83), .ZN(
        n4403) );
  MOAI22 U13333 ( .A1(n28384), .A2(n82), .B1(ram[163]), .B2(n83), .ZN(
        n4404) );
  MOAI22 U13334 ( .A1(n28149), .A2(n82), .B1(ram[164]), .B2(n83), .ZN(
        n4405) );
  MOAI22 U13335 ( .A1(n27914), .A2(n82), .B1(ram[165]), .B2(n83), .ZN(
        n4406) );
  MOAI22 U13336 ( .A1(n27679), .A2(n82), .B1(ram[166]), .B2(n83), .ZN(
        n4407) );
  MOAI22 U13337 ( .A1(n27444), .A2(n82), .B1(ram[167]), .B2(n83), .ZN(
        n4408) );
  MOAI22 U13338 ( .A1(n29089), .A2(n85), .B1(ram[168]), .B2(n86), .ZN(
        n4409) );
  MOAI22 U13339 ( .A1(n28854), .A2(n85), .B1(ram[169]), .B2(n86), .ZN(
        n4410) );
  MOAI22 U13340 ( .A1(n28619), .A2(n85), .B1(ram[170]), .B2(n86), .ZN(
        n4411) );
  MOAI22 U13341 ( .A1(n28384), .A2(n85), .B1(ram[171]), .B2(n86), .ZN(
        n4412) );
  MOAI22 U13342 ( .A1(n28149), .A2(n85), .B1(ram[172]), .B2(n86), .ZN(
        n4413) );
  MOAI22 U13343 ( .A1(n27914), .A2(n85), .B1(ram[173]), .B2(n86), .ZN(
        n4414) );
  MOAI22 U13344 ( .A1(n27679), .A2(n85), .B1(ram[174]), .B2(n86), .ZN(
        n4415) );
  MOAI22 U13345 ( .A1(n27444), .A2(n85), .B1(ram[175]), .B2(n86), .ZN(
        n4416) );
  MOAI22 U13346 ( .A1(n29089), .A2(n88), .B1(ram[176]), .B2(n89), .ZN(
        n4417) );
  MOAI22 U13347 ( .A1(n28854), .A2(n88), .B1(ram[177]), .B2(n89), .ZN(
        n4418) );
  MOAI22 U13348 ( .A1(n28619), .A2(n88), .B1(ram[178]), .B2(n89), .ZN(
        n4419) );
  MOAI22 U13349 ( .A1(n28384), .A2(n88), .B1(ram[179]), .B2(n89), .ZN(
        n4420) );
  MOAI22 U13350 ( .A1(n28149), .A2(n88), .B1(ram[180]), .B2(n89), .ZN(
        n4421) );
  MOAI22 U13351 ( .A1(n27914), .A2(n88), .B1(ram[181]), .B2(n89), .ZN(
        n4422) );
  MOAI22 U13352 ( .A1(n27679), .A2(n88), .B1(ram[182]), .B2(n89), .ZN(
        n4423) );
  MOAI22 U13353 ( .A1(n27444), .A2(n88), .B1(ram[183]), .B2(n89), .ZN(
        n4424) );
  MOAI22 U13354 ( .A1(n29089), .A2(n91), .B1(ram[184]), .B2(n92), .ZN(
        n4425) );
  MOAI22 U13355 ( .A1(n28854), .A2(n91), .B1(ram[185]), .B2(n92), .ZN(
        n4426) );
  MOAI22 U13356 ( .A1(n28619), .A2(n91), .B1(ram[186]), .B2(n92), .ZN(
        n4427) );
  MOAI22 U13357 ( .A1(n28384), .A2(n91), .B1(ram[187]), .B2(n92), .ZN(
        n4428) );
  MOAI22 U13358 ( .A1(n28149), .A2(n91), .B1(ram[188]), .B2(n92), .ZN(
        n4429) );
  MOAI22 U13359 ( .A1(n27914), .A2(n91), .B1(ram[189]), .B2(n92), .ZN(
        n4430) );
  MOAI22 U13360 ( .A1(n27679), .A2(n91), .B1(ram[190]), .B2(n92), .ZN(
        n4431) );
  MOAI22 U13361 ( .A1(n27444), .A2(n91), .B1(ram[191]), .B2(n92), .ZN(
        n4432) );
  MOAI22 U13362 ( .A1(n29089), .A2(n94), .B1(ram[192]), .B2(n95), .ZN(
        n4433) );
  MOAI22 U13363 ( .A1(n28854), .A2(n94), .B1(ram[193]), .B2(n95), .ZN(
        n4434) );
  MOAI22 U13364 ( .A1(n28619), .A2(n94), .B1(ram[194]), .B2(n95), .ZN(
        n4435) );
  MOAI22 U13365 ( .A1(n28384), .A2(n94), .B1(ram[195]), .B2(n95), .ZN(
        n4436) );
  MOAI22 U13366 ( .A1(n28149), .A2(n94), .B1(ram[196]), .B2(n95), .ZN(
        n4437) );
  MOAI22 U13367 ( .A1(n27914), .A2(n94), .B1(ram[197]), .B2(n95), .ZN(
        n4438) );
  MOAI22 U13368 ( .A1(n27679), .A2(n94), .B1(ram[198]), .B2(n95), .ZN(
        n4439) );
  MOAI22 U13369 ( .A1(n27444), .A2(n94), .B1(ram[199]), .B2(n95), .ZN(
        n4440) );
  MOAI22 U13370 ( .A1(n29089), .A2(n97), .B1(ram[200]), .B2(n98), .ZN(
        n4441) );
  MOAI22 U13371 ( .A1(n28854), .A2(n97), .B1(ram[201]), .B2(n98), .ZN(
        n4442) );
  MOAI22 U13372 ( .A1(n28619), .A2(n97), .B1(ram[202]), .B2(n98), .ZN(
        n4443) );
  MOAI22 U13373 ( .A1(n28384), .A2(n97), .B1(ram[203]), .B2(n98), .ZN(
        n4444) );
  MOAI22 U13374 ( .A1(n28149), .A2(n97), .B1(ram[204]), .B2(n98), .ZN(
        n4445) );
  MOAI22 U13375 ( .A1(n27914), .A2(n97), .B1(ram[205]), .B2(n98), .ZN(
        n4446) );
  MOAI22 U13376 ( .A1(n27679), .A2(n97), .B1(ram[206]), .B2(n98), .ZN(
        n4447) );
  MOAI22 U13377 ( .A1(n27444), .A2(n97), .B1(ram[207]), .B2(n98), .ZN(
        n4448) );
  MOAI22 U13378 ( .A1(n29090), .A2(n100), .B1(ram[208]), .B2(n101), .ZN(
        n4449) );
  MOAI22 U13379 ( .A1(n28855), .A2(n100), .B1(ram[209]), .B2(n101), .ZN(
        n4450) );
  MOAI22 U13380 ( .A1(n28620), .A2(n100), .B1(ram[210]), .B2(n101), .ZN(
        n4451) );
  MOAI22 U13381 ( .A1(n28385), .A2(n100), .B1(ram[211]), .B2(n101), .ZN(
        n4452) );
  MOAI22 U13382 ( .A1(n28150), .A2(n100), .B1(ram[212]), .B2(n101), .ZN(
        n4453) );
  MOAI22 U13383 ( .A1(n27915), .A2(n100), .B1(ram[213]), .B2(n101), .ZN(
        n4454) );
  MOAI22 U13384 ( .A1(n27680), .A2(n100), .B1(ram[214]), .B2(n101), .ZN(
        n4455) );
  MOAI22 U13385 ( .A1(n27445), .A2(n100), .B1(ram[215]), .B2(n101), .ZN(
        n4456) );
  MOAI22 U13386 ( .A1(n29090), .A2(n103), .B1(ram[216]), .B2(n104), .ZN(
        n4457) );
  MOAI22 U13387 ( .A1(n28855), .A2(n103), .B1(ram[217]), .B2(n104), .ZN(
        n4458) );
  MOAI22 U13388 ( .A1(n28620), .A2(n103), .B1(ram[218]), .B2(n104), .ZN(
        n4459) );
  MOAI22 U13389 ( .A1(n28385), .A2(n103), .B1(ram[219]), .B2(n104), .ZN(
        n4460) );
  MOAI22 U13390 ( .A1(n28150), .A2(n103), .B1(ram[220]), .B2(n104), .ZN(
        n4461) );
  MOAI22 U13391 ( .A1(n27915), .A2(n103), .B1(ram[221]), .B2(n104), .ZN(
        n4462) );
  MOAI22 U13392 ( .A1(n27680), .A2(n103), .B1(ram[222]), .B2(n104), .ZN(
        n4463) );
  MOAI22 U13393 ( .A1(n27445), .A2(n103), .B1(ram[223]), .B2(n104), .ZN(
        n4464) );
  MOAI22 U13394 ( .A1(n29090), .A2(n106), .B1(ram[224]), .B2(n107), .ZN(
        n4465) );
  MOAI22 U13395 ( .A1(n28855), .A2(n106), .B1(ram[225]), .B2(n107), .ZN(
        n4466) );
  MOAI22 U13396 ( .A1(n28620), .A2(n106), .B1(ram[226]), .B2(n107), .ZN(
        n4467) );
  MOAI22 U13397 ( .A1(n28385), .A2(n106), .B1(ram[227]), .B2(n107), .ZN(
        n4468) );
  MOAI22 U13398 ( .A1(n28150), .A2(n106), .B1(ram[228]), .B2(n107), .ZN(
        n4469) );
  MOAI22 U13399 ( .A1(n27915), .A2(n106), .B1(ram[229]), .B2(n107), .ZN(
        n4470) );
  MOAI22 U13400 ( .A1(n27680), .A2(n106), .B1(ram[230]), .B2(n107), .ZN(
        n4471) );
  MOAI22 U13401 ( .A1(n27445), .A2(n106), .B1(ram[231]), .B2(n107), .ZN(
        n4472) );
  MOAI22 U13402 ( .A1(n29090), .A2(n109), .B1(ram[232]), .B2(n110), .ZN(
        n4473) );
  MOAI22 U13403 ( .A1(n28855), .A2(n109), .B1(ram[233]), .B2(n110), .ZN(
        n4474) );
  MOAI22 U13404 ( .A1(n28620), .A2(n109), .B1(ram[234]), .B2(n110), .ZN(
        n4475) );
  MOAI22 U13405 ( .A1(n28385), .A2(n109), .B1(ram[235]), .B2(n110), .ZN(
        n4476) );
  MOAI22 U13406 ( .A1(n28150), .A2(n109), .B1(ram[236]), .B2(n110), .ZN(
        n4477) );
  MOAI22 U13407 ( .A1(n27915), .A2(n109), .B1(ram[237]), .B2(n110), .ZN(
        n4478) );
  MOAI22 U13408 ( .A1(n27680), .A2(n109), .B1(ram[238]), .B2(n110), .ZN(
        n4479) );
  MOAI22 U13409 ( .A1(n27445), .A2(n109), .B1(ram[239]), .B2(n110), .ZN(
        n4480) );
  MOAI22 U13410 ( .A1(n29090), .A2(n112), .B1(ram[240]), .B2(n113), .ZN(
        n4481) );
  MOAI22 U13411 ( .A1(n28855), .A2(n112), .B1(ram[241]), .B2(n113), .ZN(
        n4482) );
  MOAI22 U13412 ( .A1(n28620), .A2(n112), .B1(ram[242]), .B2(n113), .ZN(
        n4483) );
  MOAI22 U13413 ( .A1(n28385), .A2(n112), .B1(ram[243]), .B2(n113), .ZN(
        n4484) );
  MOAI22 U13414 ( .A1(n28150), .A2(n112), .B1(ram[244]), .B2(n113), .ZN(
        n4485) );
  MOAI22 U13415 ( .A1(n27915), .A2(n112), .B1(ram[245]), .B2(n113), .ZN(
        n4486) );
  MOAI22 U13416 ( .A1(n27680), .A2(n112), .B1(ram[246]), .B2(n113), .ZN(
        n4487) );
  MOAI22 U13417 ( .A1(n27445), .A2(n112), .B1(ram[247]), .B2(n113), .ZN(
        n4488) );
  MOAI22 U13418 ( .A1(n29090), .A2(n115), .B1(ram[248]), .B2(n116), .ZN(
        n4489) );
  MOAI22 U13419 ( .A1(n28855), .A2(n115), .B1(ram[249]), .B2(n116), .ZN(
        n4490) );
  MOAI22 U13420 ( .A1(n28620), .A2(n115), .B1(ram[250]), .B2(n116), .ZN(
        n4491) );
  MOAI22 U13421 ( .A1(n28385), .A2(n115), .B1(ram[251]), .B2(n116), .ZN(
        n4492) );
  MOAI22 U13422 ( .A1(n28150), .A2(n115), .B1(ram[252]), .B2(n116), .ZN(
        n4493) );
  MOAI22 U13423 ( .A1(n27915), .A2(n115), .B1(ram[253]), .B2(n116), .ZN(
        n4494) );
  MOAI22 U13424 ( .A1(n27680), .A2(n115), .B1(ram[254]), .B2(n116), .ZN(
        n4495) );
  MOAI22 U13425 ( .A1(n27445), .A2(n115), .B1(ram[255]), .B2(n116), .ZN(
        n4496) );
  MOAI22 U13426 ( .A1(n29090), .A2(n118), .B1(ram[256]), .B2(n119), .ZN(
        n4497) );
  MOAI22 U13427 ( .A1(n28855), .A2(n118), .B1(ram[257]), .B2(n119), .ZN(
        n4498) );
  MOAI22 U13428 ( .A1(n28620), .A2(n118), .B1(ram[258]), .B2(n119), .ZN(
        n4499) );
  MOAI22 U13429 ( .A1(n28385), .A2(n118), .B1(ram[259]), .B2(n119), .ZN(
        n4500) );
  MOAI22 U13430 ( .A1(n28150), .A2(n118), .B1(ram[260]), .B2(n119), .ZN(
        n4501) );
  MOAI22 U13431 ( .A1(n27915), .A2(n118), .B1(ram[261]), .B2(n119), .ZN(
        n4502) );
  MOAI22 U13432 ( .A1(n27680), .A2(n118), .B1(ram[262]), .B2(n119), .ZN(
        n4503) );
  MOAI22 U13433 ( .A1(n27445), .A2(n118), .B1(ram[263]), .B2(n119), .ZN(
        n4504) );
  MOAI22 U13434 ( .A1(n29090), .A2(n121), .B1(ram[264]), .B2(n122), .ZN(
        n4505) );
  MOAI22 U13435 ( .A1(n28855), .A2(n121), .B1(ram[265]), .B2(n122), .ZN(
        n4506) );
  MOAI22 U13436 ( .A1(n28620), .A2(n121), .B1(ram[266]), .B2(n122), .ZN(
        n4507) );
  MOAI22 U13437 ( .A1(n28385), .A2(n121), .B1(ram[267]), .B2(n122), .ZN(
        n4508) );
  MOAI22 U13438 ( .A1(n28150), .A2(n121), .B1(ram[268]), .B2(n122), .ZN(
        n4509) );
  MOAI22 U13439 ( .A1(n27915), .A2(n121), .B1(ram[269]), .B2(n122), .ZN(
        n4510) );
  MOAI22 U13440 ( .A1(n27680), .A2(n121), .B1(ram[270]), .B2(n122), .ZN(
        n4511) );
  MOAI22 U13441 ( .A1(n27445), .A2(n121), .B1(ram[271]), .B2(n122), .ZN(
        n4512) );
  MOAI22 U13442 ( .A1(n29090), .A2(n124), .B1(ram[272]), .B2(n125), .ZN(
        n4513) );
  MOAI22 U13443 ( .A1(n28855), .A2(n124), .B1(ram[273]), .B2(n125), .ZN(
        n4514) );
  MOAI22 U13444 ( .A1(n28620), .A2(n124), .B1(ram[274]), .B2(n125), .ZN(
        n4515) );
  MOAI22 U13445 ( .A1(n28385), .A2(n124), .B1(ram[275]), .B2(n125), .ZN(
        n4516) );
  MOAI22 U13446 ( .A1(n28150), .A2(n124), .B1(ram[276]), .B2(n125), .ZN(
        n4517) );
  MOAI22 U13447 ( .A1(n27915), .A2(n124), .B1(ram[277]), .B2(n125), .ZN(
        n4518) );
  MOAI22 U13448 ( .A1(n27680), .A2(n124), .B1(ram[278]), .B2(n125), .ZN(
        n4519) );
  MOAI22 U13449 ( .A1(n27445), .A2(n124), .B1(ram[279]), .B2(n125), .ZN(
        n4520) );
  MOAI22 U13450 ( .A1(n29090), .A2(n127), .B1(ram[280]), .B2(n128), .ZN(
        n4521) );
  MOAI22 U13451 ( .A1(n28855), .A2(n127), .B1(ram[281]), .B2(n128), .ZN(
        n4522) );
  MOAI22 U13452 ( .A1(n28620), .A2(n127), .B1(ram[282]), .B2(n128), .ZN(
        n4523) );
  MOAI22 U13453 ( .A1(n28385), .A2(n127), .B1(ram[283]), .B2(n128), .ZN(
        n4524) );
  MOAI22 U13454 ( .A1(n28150), .A2(n127), .B1(ram[284]), .B2(n128), .ZN(
        n4525) );
  MOAI22 U13455 ( .A1(n27915), .A2(n127), .B1(ram[285]), .B2(n128), .ZN(
        n4526) );
  MOAI22 U13456 ( .A1(n27680), .A2(n127), .B1(ram[286]), .B2(n128), .ZN(
        n4527) );
  MOAI22 U13457 ( .A1(n27445), .A2(n127), .B1(ram[287]), .B2(n128), .ZN(
        n4528) );
  MOAI22 U13458 ( .A1(n29090), .A2(n130), .B1(ram[288]), .B2(n131), .ZN(
        n4529) );
  MOAI22 U13459 ( .A1(n28855), .A2(n130), .B1(ram[289]), .B2(n131), .ZN(
        n4530) );
  MOAI22 U13460 ( .A1(n28620), .A2(n130), .B1(ram[290]), .B2(n131), .ZN(
        n4531) );
  MOAI22 U13461 ( .A1(n28385), .A2(n130), .B1(ram[291]), .B2(n131), .ZN(
        n4532) );
  MOAI22 U13462 ( .A1(n28150), .A2(n130), .B1(ram[292]), .B2(n131), .ZN(
        n4533) );
  MOAI22 U13463 ( .A1(n27915), .A2(n130), .B1(ram[293]), .B2(n131), .ZN(
        n4534) );
  MOAI22 U13464 ( .A1(n27680), .A2(n130), .B1(ram[294]), .B2(n131), .ZN(
        n4535) );
  MOAI22 U13465 ( .A1(n27445), .A2(n130), .B1(ram[295]), .B2(n131), .ZN(
        n4536) );
  MOAI22 U13466 ( .A1(n29090), .A2(n133), .B1(ram[296]), .B2(n134), .ZN(
        n4537) );
  MOAI22 U13467 ( .A1(n28855), .A2(n133), .B1(ram[297]), .B2(n134), .ZN(
        n4538) );
  MOAI22 U13468 ( .A1(n28620), .A2(n133), .B1(ram[298]), .B2(n134), .ZN(
        n4539) );
  MOAI22 U13469 ( .A1(n28385), .A2(n133), .B1(ram[299]), .B2(n134), .ZN(
        n4540) );
  MOAI22 U13470 ( .A1(n28150), .A2(n133), .B1(ram[300]), .B2(n134), .ZN(
        n4541) );
  MOAI22 U13471 ( .A1(n27915), .A2(n133), .B1(ram[301]), .B2(n134), .ZN(
        n4542) );
  MOAI22 U13472 ( .A1(n27680), .A2(n133), .B1(ram[302]), .B2(n134), .ZN(
        n4543) );
  MOAI22 U13473 ( .A1(n27445), .A2(n133), .B1(ram[303]), .B2(n134), .ZN(
        n4544) );
  MOAI22 U13474 ( .A1(n29090), .A2(n136), .B1(ram[304]), .B2(n137), .ZN(
        n4545) );
  MOAI22 U13475 ( .A1(n28855), .A2(n136), .B1(ram[305]), .B2(n137), .ZN(
        n4546) );
  MOAI22 U13476 ( .A1(n28620), .A2(n136), .B1(ram[306]), .B2(n137), .ZN(
        n4547) );
  MOAI22 U13477 ( .A1(n28385), .A2(n136), .B1(ram[307]), .B2(n137), .ZN(
        n4548) );
  MOAI22 U13478 ( .A1(n28150), .A2(n136), .B1(ram[308]), .B2(n137), .ZN(
        n4549) );
  MOAI22 U13479 ( .A1(n27915), .A2(n136), .B1(ram[309]), .B2(n137), .ZN(
        n4550) );
  MOAI22 U13480 ( .A1(n27680), .A2(n136), .B1(ram[310]), .B2(n137), .ZN(
        n4551) );
  MOAI22 U13481 ( .A1(n27445), .A2(n136), .B1(ram[311]), .B2(n137), .ZN(
        n4552) );
  MOAI22 U13482 ( .A1(n29091), .A2(n139), .B1(ram[312]), .B2(n140), .ZN(
        n4553) );
  MOAI22 U13483 ( .A1(n28856), .A2(n139), .B1(ram[313]), .B2(n140), .ZN(
        n4554) );
  MOAI22 U13484 ( .A1(n28621), .A2(n139), .B1(ram[314]), .B2(n140), .ZN(
        n4555) );
  MOAI22 U13485 ( .A1(n28386), .A2(n139), .B1(ram[315]), .B2(n140), .ZN(
        n4556) );
  MOAI22 U13486 ( .A1(n28151), .A2(n139), .B1(ram[316]), .B2(n140), .ZN(
        n4557) );
  MOAI22 U13487 ( .A1(n27916), .A2(n139), .B1(ram[317]), .B2(n140), .ZN(
        n4558) );
  MOAI22 U13488 ( .A1(n27681), .A2(n139), .B1(ram[318]), .B2(n140), .ZN(
        n4559) );
  MOAI22 U13489 ( .A1(n27446), .A2(n139), .B1(ram[319]), .B2(n140), .ZN(
        n4560) );
  MOAI22 U13490 ( .A1(n29091), .A2(n142), .B1(ram[320]), .B2(n143), .ZN(
        n4561) );
  MOAI22 U13491 ( .A1(n28856), .A2(n142), .B1(ram[321]), .B2(n143), .ZN(
        n4562) );
  MOAI22 U13492 ( .A1(n28621), .A2(n142), .B1(ram[322]), .B2(n143), .ZN(
        n4563) );
  MOAI22 U13493 ( .A1(n28386), .A2(n142), .B1(ram[323]), .B2(n143), .ZN(
        n4564) );
  MOAI22 U13494 ( .A1(n28151), .A2(n142), .B1(ram[324]), .B2(n143), .ZN(
        n4565) );
  MOAI22 U13495 ( .A1(n27916), .A2(n142), .B1(ram[325]), .B2(n143), .ZN(
        n4566) );
  MOAI22 U13496 ( .A1(n27681), .A2(n142), .B1(ram[326]), .B2(n143), .ZN(
        n4567) );
  MOAI22 U13497 ( .A1(n27446), .A2(n142), .B1(ram[327]), .B2(n143), .ZN(
        n4568) );
  MOAI22 U13498 ( .A1(n29091), .A2(n145), .B1(ram[328]), .B2(n146), .ZN(
        n4569) );
  MOAI22 U13499 ( .A1(n28856), .A2(n145), .B1(ram[329]), .B2(n146), .ZN(
        n4570) );
  MOAI22 U13500 ( .A1(n28621), .A2(n145), .B1(ram[330]), .B2(n146), .ZN(
        n4571) );
  MOAI22 U13501 ( .A1(n28386), .A2(n145), .B1(ram[331]), .B2(n146), .ZN(
        n4572) );
  MOAI22 U13502 ( .A1(n28151), .A2(n145), .B1(ram[332]), .B2(n146), .ZN(
        n4573) );
  MOAI22 U13503 ( .A1(n27916), .A2(n145), .B1(ram[333]), .B2(n146), .ZN(
        n4574) );
  MOAI22 U13504 ( .A1(n27681), .A2(n145), .B1(ram[334]), .B2(n146), .ZN(
        n4575) );
  MOAI22 U13505 ( .A1(n27446), .A2(n145), .B1(ram[335]), .B2(n146), .ZN(
        n4576) );
  MOAI22 U13506 ( .A1(n29091), .A2(n148), .B1(ram[336]), .B2(n149), .ZN(
        n4577) );
  MOAI22 U13507 ( .A1(n28856), .A2(n148), .B1(ram[337]), .B2(n149), .ZN(
        n4578) );
  MOAI22 U13508 ( .A1(n28621), .A2(n148), .B1(ram[338]), .B2(n149), .ZN(
        n4579) );
  MOAI22 U13509 ( .A1(n28386), .A2(n148), .B1(ram[339]), .B2(n149), .ZN(
        n4580) );
  MOAI22 U13510 ( .A1(n28151), .A2(n148), .B1(ram[340]), .B2(n149), .ZN(
        n4581) );
  MOAI22 U13511 ( .A1(n27916), .A2(n148), .B1(ram[341]), .B2(n149), .ZN(
        n4582) );
  MOAI22 U13512 ( .A1(n27681), .A2(n148), .B1(ram[342]), .B2(n149), .ZN(
        n4583) );
  MOAI22 U13513 ( .A1(n27446), .A2(n148), .B1(ram[343]), .B2(n149), .ZN(
        n4584) );
  MOAI22 U13514 ( .A1(n29091), .A2(n151), .B1(ram[344]), .B2(n152), .ZN(
        n4585) );
  MOAI22 U13515 ( .A1(n28856), .A2(n151), .B1(ram[345]), .B2(n152), .ZN(
        n4586) );
  MOAI22 U13516 ( .A1(n28621), .A2(n151), .B1(ram[346]), .B2(n152), .ZN(
        n4587) );
  MOAI22 U13517 ( .A1(n28386), .A2(n151), .B1(ram[347]), .B2(n152), .ZN(
        n4588) );
  MOAI22 U13518 ( .A1(n28151), .A2(n151), .B1(ram[348]), .B2(n152), .ZN(
        n4589) );
  MOAI22 U13519 ( .A1(n27916), .A2(n151), .B1(ram[349]), .B2(n152), .ZN(
        n4590) );
  MOAI22 U13520 ( .A1(n27681), .A2(n151), .B1(ram[350]), .B2(n152), .ZN(
        n4591) );
  MOAI22 U13521 ( .A1(n27446), .A2(n151), .B1(ram[351]), .B2(n152), .ZN(
        n4592) );
  MOAI22 U13522 ( .A1(n29091), .A2(n154), .B1(ram[352]), .B2(n155), .ZN(
        n4593) );
  MOAI22 U13523 ( .A1(n28856), .A2(n154), .B1(ram[353]), .B2(n155), .ZN(
        n4594) );
  MOAI22 U13524 ( .A1(n28621), .A2(n154), .B1(ram[354]), .B2(n155), .ZN(
        n4595) );
  MOAI22 U13525 ( .A1(n28386), .A2(n154), .B1(ram[355]), .B2(n155), .ZN(
        n4596) );
  MOAI22 U13526 ( .A1(n28151), .A2(n154), .B1(ram[356]), .B2(n155), .ZN(
        n4597) );
  MOAI22 U13527 ( .A1(n27916), .A2(n154), .B1(ram[357]), .B2(n155), .ZN(
        n4598) );
  MOAI22 U13528 ( .A1(n27681), .A2(n154), .B1(ram[358]), .B2(n155), .ZN(
        n4599) );
  MOAI22 U13529 ( .A1(n27446), .A2(n154), .B1(ram[359]), .B2(n155), .ZN(
        n4600) );
  MOAI22 U13530 ( .A1(n29091), .A2(n157), .B1(ram[360]), .B2(n158), .ZN(
        n4601) );
  MOAI22 U13531 ( .A1(n28856), .A2(n157), .B1(ram[361]), .B2(n158), .ZN(
        n4602) );
  MOAI22 U13532 ( .A1(n28621), .A2(n157), .B1(ram[362]), .B2(n158), .ZN(
        n4603) );
  MOAI22 U13533 ( .A1(n28386), .A2(n157), .B1(ram[363]), .B2(n158), .ZN(
        n4604) );
  MOAI22 U13534 ( .A1(n28151), .A2(n157), .B1(ram[364]), .B2(n158), .ZN(
        n4605) );
  MOAI22 U13535 ( .A1(n27916), .A2(n157), .B1(ram[365]), .B2(n158), .ZN(
        n4606) );
  MOAI22 U13536 ( .A1(n27681), .A2(n157), .B1(ram[366]), .B2(n158), .ZN(
        n4607) );
  MOAI22 U13537 ( .A1(n27446), .A2(n157), .B1(ram[367]), .B2(n158), .ZN(
        n4608) );
  MOAI22 U13538 ( .A1(n29091), .A2(n160), .B1(ram[368]), .B2(n161), .ZN(
        n4609) );
  MOAI22 U13539 ( .A1(n28856), .A2(n160), .B1(ram[369]), .B2(n161), .ZN(
        n4610) );
  MOAI22 U13540 ( .A1(n28621), .A2(n160), .B1(ram[370]), .B2(n161), .ZN(
        n4611) );
  MOAI22 U13541 ( .A1(n28386), .A2(n160), .B1(ram[371]), .B2(n161), .ZN(
        n4612) );
  MOAI22 U13542 ( .A1(n28151), .A2(n160), .B1(ram[372]), .B2(n161), .ZN(
        n4613) );
  MOAI22 U13543 ( .A1(n27916), .A2(n160), .B1(ram[373]), .B2(n161), .ZN(
        n4614) );
  MOAI22 U13544 ( .A1(n27681), .A2(n160), .B1(ram[374]), .B2(n161), .ZN(
        n4615) );
  MOAI22 U13545 ( .A1(n27446), .A2(n160), .B1(ram[375]), .B2(n161), .ZN(
        n4616) );
  MOAI22 U13546 ( .A1(n29091), .A2(n163), .B1(ram[376]), .B2(n164), .ZN(
        n4617) );
  MOAI22 U13547 ( .A1(n28856), .A2(n163), .B1(ram[377]), .B2(n164), .ZN(
        n4618) );
  MOAI22 U13548 ( .A1(n28621), .A2(n163), .B1(ram[378]), .B2(n164), .ZN(
        n4619) );
  MOAI22 U13549 ( .A1(n28386), .A2(n163), .B1(ram[379]), .B2(n164), .ZN(
        n4620) );
  MOAI22 U13550 ( .A1(n28151), .A2(n163), .B1(ram[380]), .B2(n164), .ZN(
        n4621) );
  MOAI22 U13551 ( .A1(n27916), .A2(n163), .B1(ram[381]), .B2(n164), .ZN(
        n4622) );
  MOAI22 U13552 ( .A1(n27681), .A2(n163), .B1(ram[382]), .B2(n164), .ZN(
        n4623) );
  MOAI22 U13553 ( .A1(n27446), .A2(n163), .B1(ram[383]), .B2(n164), .ZN(
        n4624) );
  MOAI22 U13554 ( .A1(n29091), .A2(n166), .B1(ram[384]), .B2(n167), .ZN(
        n4625) );
  MOAI22 U13555 ( .A1(n28856), .A2(n166), .B1(ram[385]), .B2(n167), .ZN(
        n4626) );
  MOAI22 U13556 ( .A1(n28621), .A2(n166), .B1(ram[386]), .B2(n167), .ZN(
        n4627) );
  MOAI22 U13557 ( .A1(n28386), .A2(n166), .B1(ram[387]), .B2(n167), .ZN(
        n4628) );
  MOAI22 U13558 ( .A1(n28151), .A2(n166), .B1(ram[388]), .B2(n167), .ZN(
        n4629) );
  MOAI22 U13559 ( .A1(n27916), .A2(n166), .B1(ram[389]), .B2(n167), .ZN(
        n4630) );
  MOAI22 U13560 ( .A1(n27681), .A2(n166), .B1(ram[390]), .B2(n167), .ZN(
        n4631) );
  MOAI22 U13561 ( .A1(n27446), .A2(n166), .B1(ram[391]), .B2(n167), .ZN(
        n4632) );
  MOAI22 U13562 ( .A1(n29091), .A2(n169), .B1(ram[392]), .B2(n170), .ZN(
        n4633) );
  MOAI22 U13563 ( .A1(n28856), .A2(n169), .B1(ram[393]), .B2(n170), .ZN(
        n4634) );
  MOAI22 U13564 ( .A1(n28621), .A2(n169), .B1(ram[394]), .B2(n170), .ZN(
        n4635) );
  MOAI22 U13565 ( .A1(n28386), .A2(n169), .B1(ram[395]), .B2(n170), .ZN(
        n4636) );
  MOAI22 U13566 ( .A1(n28151), .A2(n169), .B1(ram[396]), .B2(n170), .ZN(
        n4637) );
  MOAI22 U13567 ( .A1(n27916), .A2(n169), .B1(ram[397]), .B2(n170), .ZN(
        n4638) );
  MOAI22 U13568 ( .A1(n27681), .A2(n169), .B1(ram[398]), .B2(n170), .ZN(
        n4639) );
  MOAI22 U13569 ( .A1(n27446), .A2(n169), .B1(ram[399]), .B2(n170), .ZN(
        n4640) );
  MOAI22 U13570 ( .A1(n29091), .A2(n172), .B1(ram[400]), .B2(n173), .ZN(
        n4641) );
  MOAI22 U13571 ( .A1(n28856), .A2(n172), .B1(ram[401]), .B2(n173), .ZN(
        n4642) );
  MOAI22 U13572 ( .A1(n28621), .A2(n172), .B1(ram[402]), .B2(n173), .ZN(
        n4643) );
  MOAI22 U13573 ( .A1(n28386), .A2(n172), .B1(ram[403]), .B2(n173), .ZN(
        n4644) );
  MOAI22 U13574 ( .A1(n28151), .A2(n172), .B1(ram[404]), .B2(n173), .ZN(
        n4645) );
  MOAI22 U13575 ( .A1(n27916), .A2(n172), .B1(ram[405]), .B2(n173), .ZN(
        n4646) );
  MOAI22 U13576 ( .A1(n27681), .A2(n172), .B1(ram[406]), .B2(n173), .ZN(
        n4647) );
  MOAI22 U13577 ( .A1(n27446), .A2(n172), .B1(ram[407]), .B2(n173), .ZN(
        n4648) );
  MOAI22 U13578 ( .A1(n29091), .A2(n175), .B1(ram[408]), .B2(n176), .ZN(
        n4649) );
  MOAI22 U13579 ( .A1(n28856), .A2(n175), .B1(ram[409]), .B2(n176), .ZN(
        n4650) );
  MOAI22 U13580 ( .A1(n28621), .A2(n175), .B1(ram[410]), .B2(n176), .ZN(
        n4651) );
  MOAI22 U13581 ( .A1(n28386), .A2(n175), .B1(ram[411]), .B2(n176), .ZN(
        n4652) );
  MOAI22 U13582 ( .A1(n28151), .A2(n175), .B1(ram[412]), .B2(n176), .ZN(
        n4653) );
  MOAI22 U13583 ( .A1(n27916), .A2(n175), .B1(ram[413]), .B2(n176), .ZN(
        n4654) );
  MOAI22 U13584 ( .A1(n27681), .A2(n175), .B1(ram[414]), .B2(n176), .ZN(
        n4655) );
  MOAI22 U13585 ( .A1(n27446), .A2(n175), .B1(ram[415]), .B2(n176), .ZN(
        n4656) );
  MOAI22 U13586 ( .A1(n29092), .A2(n178), .B1(ram[416]), .B2(n179), .ZN(
        n4657) );
  MOAI22 U13587 ( .A1(n28857), .A2(n178), .B1(ram[417]), .B2(n179), .ZN(
        n4658) );
  MOAI22 U13588 ( .A1(n28622), .A2(n178), .B1(ram[418]), .B2(n179), .ZN(
        n4659) );
  MOAI22 U13589 ( .A1(n28387), .A2(n178), .B1(ram[419]), .B2(n179), .ZN(
        n4660) );
  MOAI22 U13590 ( .A1(n28152), .A2(n178), .B1(ram[420]), .B2(n179), .ZN(
        n4661) );
  MOAI22 U13591 ( .A1(n27917), .A2(n178), .B1(ram[421]), .B2(n179), .ZN(
        n4662) );
  MOAI22 U13592 ( .A1(n27682), .A2(n178), .B1(ram[422]), .B2(n179), .ZN(
        n4663) );
  MOAI22 U13593 ( .A1(n27447), .A2(n178), .B1(ram[423]), .B2(n179), .ZN(
        n4664) );
  MOAI22 U13594 ( .A1(n29092), .A2(n181), .B1(ram[424]), .B2(n182), .ZN(
        n4665) );
  MOAI22 U13595 ( .A1(n28857), .A2(n181), .B1(ram[425]), .B2(n182), .ZN(
        n4666) );
  MOAI22 U13596 ( .A1(n28622), .A2(n181), .B1(ram[426]), .B2(n182), .ZN(
        n4667) );
  MOAI22 U13597 ( .A1(n28387), .A2(n181), .B1(ram[427]), .B2(n182), .ZN(
        n4668) );
  MOAI22 U13598 ( .A1(n28152), .A2(n181), .B1(ram[428]), .B2(n182), .ZN(
        n4669) );
  MOAI22 U13599 ( .A1(n27917), .A2(n181), .B1(ram[429]), .B2(n182), .ZN(
        n4670) );
  MOAI22 U13600 ( .A1(n27682), .A2(n181), .B1(ram[430]), .B2(n182), .ZN(
        n4671) );
  MOAI22 U13601 ( .A1(n27447), .A2(n181), .B1(ram[431]), .B2(n182), .ZN(
        n4672) );
  MOAI22 U13602 ( .A1(n29092), .A2(n184), .B1(ram[432]), .B2(n185), .ZN(
        n4673) );
  MOAI22 U13603 ( .A1(n28857), .A2(n184), .B1(ram[433]), .B2(n185), .ZN(
        n4674) );
  MOAI22 U13604 ( .A1(n28622), .A2(n184), .B1(ram[434]), .B2(n185), .ZN(
        n4675) );
  MOAI22 U13605 ( .A1(n28387), .A2(n184), .B1(ram[435]), .B2(n185), .ZN(
        n4676) );
  MOAI22 U13606 ( .A1(n28152), .A2(n184), .B1(ram[436]), .B2(n185), .ZN(
        n4677) );
  MOAI22 U13607 ( .A1(n27917), .A2(n184), .B1(ram[437]), .B2(n185), .ZN(
        n4678) );
  MOAI22 U13608 ( .A1(n27682), .A2(n184), .B1(ram[438]), .B2(n185), .ZN(
        n4679) );
  MOAI22 U13609 ( .A1(n27447), .A2(n184), .B1(ram[439]), .B2(n185), .ZN(
        n4680) );
  MOAI22 U13610 ( .A1(n29092), .A2(n187), .B1(ram[440]), .B2(n188), .ZN(
        n4681) );
  MOAI22 U13611 ( .A1(n28857), .A2(n187), .B1(ram[441]), .B2(n188), .ZN(
        n4682) );
  MOAI22 U13612 ( .A1(n28622), .A2(n187), .B1(ram[442]), .B2(n188), .ZN(
        n4683) );
  MOAI22 U13613 ( .A1(n28387), .A2(n187), .B1(ram[443]), .B2(n188), .ZN(
        n4684) );
  MOAI22 U13614 ( .A1(n28152), .A2(n187), .B1(ram[444]), .B2(n188), .ZN(
        n4685) );
  MOAI22 U13615 ( .A1(n27917), .A2(n187), .B1(ram[445]), .B2(n188), .ZN(
        n4686) );
  MOAI22 U13616 ( .A1(n27682), .A2(n187), .B1(ram[446]), .B2(n188), .ZN(
        n4687) );
  MOAI22 U13617 ( .A1(n27447), .A2(n187), .B1(ram[447]), .B2(n188), .ZN(
        n4688) );
  MOAI22 U13618 ( .A1(n29092), .A2(n190), .B1(ram[448]), .B2(n191), .ZN(
        n4689) );
  MOAI22 U13619 ( .A1(n28857), .A2(n190), .B1(ram[449]), .B2(n191), .ZN(
        n4690) );
  MOAI22 U13620 ( .A1(n28622), .A2(n190), .B1(ram[450]), .B2(n191), .ZN(
        n4691) );
  MOAI22 U13621 ( .A1(n28387), .A2(n190), .B1(ram[451]), .B2(n191), .ZN(
        n4692) );
  MOAI22 U13622 ( .A1(n28152), .A2(n190), .B1(ram[452]), .B2(n191), .ZN(
        n4693) );
  MOAI22 U13623 ( .A1(n27917), .A2(n190), .B1(ram[453]), .B2(n191), .ZN(
        n4694) );
  MOAI22 U13624 ( .A1(n27682), .A2(n190), .B1(ram[454]), .B2(n191), .ZN(
        n4695) );
  MOAI22 U13625 ( .A1(n27447), .A2(n190), .B1(ram[455]), .B2(n191), .ZN(
        n4696) );
  MOAI22 U13626 ( .A1(n29092), .A2(n193), .B1(ram[456]), .B2(n194), .ZN(
        n4697) );
  MOAI22 U13627 ( .A1(n28857), .A2(n193), .B1(ram[457]), .B2(n194), .ZN(
        n4698) );
  MOAI22 U13628 ( .A1(n28622), .A2(n193), .B1(ram[458]), .B2(n194), .ZN(
        n4699) );
  MOAI22 U13629 ( .A1(n28387), .A2(n193), .B1(ram[459]), .B2(n194), .ZN(
        n4700) );
  MOAI22 U13630 ( .A1(n28152), .A2(n193), .B1(ram[460]), .B2(n194), .ZN(
        n4701) );
  MOAI22 U13631 ( .A1(n27917), .A2(n193), .B1(ram[461]), .B2(n194), .ZN(
        n4702) );
  MOAI22 U13632 ( .A1(n27682), .A2(n193), .B1(ram[462]), .B2(n194), .ZN(
        n4703) );
  MOAI22 U13633 ( .A1(n27447), .A2(n193), .B1(ram[463]), .B2(n194), .ZN(
        n4704) );
  MOAI22 U13634 ( .A1(n29092), .A2(n196), .B1(ram[464]), .B2(n197), .ZN(
        n4705) );
  MOAI22 U13635 ( .A1(n28857), .A2(n196), .B1(ram[465]), .B2(n197), .ZN(
        n4706) );
  MOAI22 U13636 ( .A1(n28622), .A2(n196), .B1(ram[466]), .B2(n197), .ZN(
        n4707) );
  MOAI22 U13637 ( .A1(n28387), .A2(n196), .B1(ram[467]), .B2(n197), .ZN(
        n4708) );
  MOAI22 U13638 ( .A1(n28152), .A2(n196), .B1(ram[468]), .B2(n197), .ZN(
        n4709) );
  MOAI22 U13639 ( .A1(n27917), .A2(n196), .B1(ram[469]), .B2(n197), .ZN(
        n4710) );
  MOAI22 U13640 ( .A1(n27682), .A2(n196), .B1(ram[470]), .B2(n197), .ZN(
        n4711) );
  MOAI22 U13641 ( .A1(n27447), .A2(n196), .B1(ram[471]), .B2(n197), .ZN(
        n4712) );
  MOAI22 U13642 ( .A1(n29092), .A2(n199), .B1(ram[472]), .B2(n200), .ZN(
        n4713) );
  MOAI22 U13643 ( .A1(n28857), .A2(n199), .B1(ram[473]), .B2(n200), .ZN(
        n4714) );
  MOAI22 U13644 ( .A1(n28622), .A2(n199), .B1(ram[474]), .B2(n200), .ZN(
        n4715) );
  MOAI22 U13645 ( .A1(n28387), .A2(n199), .B1(ram[475]), .B2(n200), .ZN(
        n4716) );
  MOAI22 U13646 ( .A1(n28152), .A2(n199), .B1(ram[476]), .B2(n200), .ZN(
        n4717) );
  MOAI22 U13647 ( .A1(n27917), .A2(n199), .B1(ram[477]), .B2(n200), .ZN(
        n4718) );
  MOAI22 U13648 ( .A1(n27682), .A2(n199), .B1(ram[478]), .B2(n200), .ZN(
        n4719) );
  MOAI22 U13649 ( .A1(n27447), .A2(n199), .B1(ram[479]), .B2(n200), .ZN(
        n4720) );
  MOAI22 U13650 ( .A1(n29092), .A2(n202), .B1(ram[480]), .B2(n203), .ZN(
        n4721) );
  MOAI22 U13651 ( .A1(n28857), .A2(n202), .B1(ram[481]), .B2(n203), .ZN(
        n4722) );
  MOAI22 U13652 ( .A1(n28622), .A2(n202), .B1(ram[482]), .B2(n203), .ZN(
        n4723) );
  MOAI22 U13653 ( .A1(n28387), .A2(n202), .B1(ram[483]), .B2(n203), .ZN(
        n4724) );
  MOAI22 U13654 ( .A1(n28152), .A2(n202), .B1(ram[484]), .B2(n203), .ZN(
        n4725) );
  MOAI22 U13655 ( .A1(n27917), .A2(n202), .B1(ram[485]), .B2(n203), .ZN(
        n4726) );
  MOAI22 U13656 ( .A1(n27682), .A2(n202), .B1(ram[486]), .B2(n203), .ZN(
        n4727) );
  MOAI22 U13657 ( .A1(n27447), .A2(n202), .B1(ram[487]), .B2(n203), .ZN(
        n4728) );
  MOAI22 U13658 ( .A1(n29092), .A2(n205), .B1(ram[488]), .B2(n206), .ZN(
        n4729) );
  MOAI22 U13659 ( .A1(n28857), .A2(n205), .B1(ram[489]), .B2(n206), .ZN(
        n4730) );
  MOAI22 U13660 ( .A1(n28622), .A2(n205), .B1(ram[490]), .B2(n206), .ZN(
        n4731) );
  MOAI22 U13661 ( .A1(n28387), .A2(n205), .B1(ram[491]), .B2(n206), .ZN(
        n4732) );
  MOAI22 U13662 ( .A1(n28152), .A2(n205), .B1(ram[492]), .B2(n206), .ZN(
        n4733) );
  MOAI22 U13663 ( .A1(n27917), .A2(n205), .B1(ram[493]), .B2(n206), .ZN(
        n4734) );
  MOAI22 U13664 ( .A1(n27682), .A2(n205), .B1(ram[494]), .B2(n206), .ZN(
        n4735) );
  MOAI22 U13665 ( .A1(n27447), .A2(n205), .B1(ram[495]), .B2(n206), .ZN(
        n4736) );
  MOAI22 U13666 ( .A1(n29092), .A2(n208), .B1(ram[496]), .B2(n209), .ZN(
        n4737) );
  MOAI22 U13667 ( .A1(n28857), .A2(n208), .B1(ram[497]), .B2(n209), .ZN(
        n4738) );
  MOAI22 U13668 ( .A1(n28622), .A2(n208), .B1(ram[498]), .B2(n209), .ZN(
        n4739) );
  MOAI22 U13669 ( .A1(n28387), .A2(n208), .B1(ram[499]), .B2(n209), .ZN(
        n4740) );
  MOAI22 U13670 ( .A1(n28152), .A2(n208), .B1(ram[500]), .B2(n209), .ZN(
        n4741) );
  MOAI22 U13671 ( .A1(n27917), .A2(n208), .B1(ram[501]), .B2(n209), .ZN(
        n4742) );
  MOAI22 U13672 ( .A1(n27682), .A2(n208), .B1(ram[502]), .B2(n209), .ZN(
        n4743) );
  MOAI22 U13673 ( .A1(n27447), .A2(n208), .B1(ram[503]), .B2(n209), .ZN(
        n4744) );
  MOAI22 U13674 ( .A1(n29092), .A2(n211), .B1(ram[504]), .B2(n212), .ZN(
        n4745) );
  MOAI22 U13675 ( .A1(n28857), .A2(n211), .B1(ram[505]), .B2(n212), .ZN(
        n4746) );
  MOAI22 U13676 ( .A1(n28622), .A2(n211), .B1(ram[506]), .B2(n212), .ZN(
        n4747) );
  MOAI22 U13677 ( .A1(n28387), .A2(n211), .B1(ram[507]), .B2(n212), .ZN(
        n4748) );
  MOAI22 U13678 ( .A1(n28152), .A2(n211), .B1(ram[508]), .B2(n212), .ZN(
        n4749) );
  MOAI22 U13679 ( .A1(n27917), .A2(n211), .B1(ram[509]), .B2(n212), .ZN(
        n4750) );
  MOAI22 U13680 ( .A1(n27682), .A2(n211), .B1(ram[510]), .B2(n212), .ZN(
        n4751) );
  MOAI22 U13681 ( .A1(n27447), .A2(n211), .B1(ram[511]), .B2(n212), .ZN(
        n4752) );
  MOAI22 U13682 ( .A1(n29092), .A2(n216), .B1(ram[512]), .B2(n217), .ZN(
        n4753) );
  MOAI22 U13683 ( .A1(n28857), .A2(n216), .B1(ram[513]), .B2(n217), .ZN(
        n4754) );
  MOAI22 U13684 ( .A1(n28622), .A2(n216), .B1(ram[514]), .B2(n217), .ZN(
        n4755) );
  MOAI22 U13685 ( .A1(n28387), .A2(n216), .B1(ram[515]), .B2(n217), .ZN(
        n4756) );
  MOAI22 U13686 ( .A1(n28152), .A2(n216), .B1(ram[516]), .B2(n217), .ZN(
        n4757) );
  MOAI22 U13687 ( .A1(n27917), .A2(n216), .B1(ram[517]), .B2(n217), .ZN(
        n4758) );
  MOAI22 U13688 ( .A1(n27682), .A2(n216), .B1(ram[518]), .B2(n217), .ZN(
        n4759) );
  MOAI22 U13689 ( .A1(n27447), .A2(n216), .B1(ram[519]), .B2(n217), .ZN(
        n4760) );
  MOAI22 U13690 ( .A1(n29093), .A2(n219), .B1(ram[520]), .B2(n220), .ZN(
        n4761) );
  MOAI22 U13691 ( .A1(n28858), .A2(n219), .B1(ram[521]), .B2(n220), .ZN(
        n4762) );
  MOAI22 U13692 ( .A1(n28623), .A2(n219), .B1(ram[522]), .B2(n220), .ZN(
        n4763) );
  MOAI22 U13693 ( .A1(n28388), .A2(n219), .B1(ram[523]), .B2(n220), .ZN(
        n4764) );
  MOAI22 U13694 ( .A1(n28153), .A2(n219), .B1(ram[524]), .B2(n220), .ZN(
        n4765) );
  MOAI22 U13695 ( .A1(n27918), .A2(n219), .B1(ram[525]), .B2(n220), .ZN(
        n4766) );
  MOAI22 U13696 ( .A1(n27683), .A2(n219), .B1(ram[526]), .B2(n220), .ZN(
        n4767) );
  MOAI22 U13697 ( .A1(n27448), .A2(n219), .B1(ram[527]), .B2(n220), .ZN(
        n4768) );
  MOAI22 U13698 ( .A1(n29093), .A2(n221), .B1(ram[528]), .B2(n222), .ZN(
        n4769) );
  MOAI22 U13699 ( .A1(n28858), .A2(n221), .B1(ram[529]), .B2(n222), .ZN(
        n4770) );
  MOAI22 U13700 ( .A1(n28623), .A2(n221), .B1(ram[530]), .B2(n222), .ZN(
        n4771) );
  MOAI22 U13701 ( .A1(n28388), .A2(n221), .B1(ram[531]), .B2(n222), .ZN(
        n4772) );
  MOAI22 U13702 ( .A1(n28153), .A2(n221), .B1(ram[532]), .B2(n222), .ZN(
        n4773) );
  MOAI22 U13703 ( .A1(n27918), .A2(n221), .B1(ram[533]), .B2(n222), .ZN(
        n4774) );
  MOAI22 U13704 ( .A1(n27683), .A2(n221), .B1(ram[534]), .B2(n222), .ZN(
        n4775) );
  MOAI22 U13705 ( .A1(n27448), .A2(n221), .B1(ram[535]), .B2(n222), .ZN(
        n4776) );
  MOAI22 U13706 ( .A1(n29093), .A2(n223), .B1(ram[536]), .B2(n224), .ZN(
        n4777) );
  MOAI22 U13707 ( .A1(n28858), .A2(n223), .B1(ram[537]), .B2(n224), .ZN(
        n4778) );
  MOAI22 U13708 ( .A1(n28623), .A2(n223), .B1(ram[538]), .B2(n224), .ZN(
        n4779) );
  MOAI22 U13709 ( .A1(n28388), .A2(n223), .B1(ram[539]), .B2(n224), .ZN(
        n4780) );
  MOAI22 U13710 ( .A1(n28153), .A2(n223), .B1(ram[540]), .B2(n224), .ZN(
        n4781) );
  MOAI22 U13711 ( .A1(n27918), .A2(n223), .B1(ram[541]), .B2(n224), .ZN(
        n4782) );
  MOAI22 U13712 ( .A1(n27683), .A2(n223), .B1(ram[542]), .B2(n224), .ZN(
        n4783) );
  MOAI22 U13713 ( .A1(n27448), .A2(n223), .B1(ram[543]), .B2(n224), .ZN(
        n4784) );
  MOAI22 U13714 ( .A1(n29093), .A2(n225), .B1(ram[544]), .B2(n226), .ZN(
        n4785) );
  MOAI22 U13715 ( .A1(n28858), .A2(n225), .B1(ram[545]), .B2(n226), .ZN(
        n4786) );
  MOAI22 U13716 ( .A1(n28623), .A2(n225), .B1(ram[546]), .B2(n226), .ZN(
        n4787) );
  MOAI22 U13717 ( .A1(n28388), .A2(n225), .B1(ram[547]), .B2(n226), .ZN(
        n4788) );
  MOAI22 U13718 ( .A1(n28153), .A2(n225), .B1(ram[548]), .B2(n226), .ZN(
        n4789) );
  MOAI22 U13719 ( .A1(n27918), .A2(n225), .B1(ram[549]), .B2(n226), .ZN(
        n4790) );
  MOAI22 U13720 ( .A1(n27683), .A2(n225), .B1(ram[550]), .B2(n226), .ZN(
        n4791) );
  MOAI22 U13721 ( .A1(n27448), .A2(n225), .B1(ram[551]), .B2(n226), .ZN(
        n4792) );
  MOAI22 U13722 ( .A1(n29093), .A2(n227), .B1(ram[552]), .B2(n228), .ZN(
        n4793) );
  MOAI22 U13723 ( .A1(n28858), .A2(n227), .B1(ram[553]), .B2(n228), .ZN(
        n4794) );
  MOAI22 U13724 ( .A1(n28623), .A2(n227), .B1(ram[554]), .B2(n228), .ZN(
        n4795) );
  MOAI22 U13725 ( .A1(n28388), .A2(n227), .B1(ram[555]), .B2(n228), .ZN(
        n4796) );
  MOAI22 U13726 ( .A1(n28153), .A2(n227), .B1(ram[556]), .B2(n228), .ZN(
        n4797) );
  MOAI22 U13727 ( .A1(n27918), .A2(n227), .B1(ram[557]), .B2(n228), .ZN(
        n4798) );
  MOAI22 U13728 ( .A1(n27683), .A2(n227), .B1(ram[558]), .B2(n228), .ZN(
        n4799) );
  MOAI22 U13729 ( .A1(n27448), .A2(n227), .B1(ram[559]), .B2(n228), .ZN(
        n4800) );
  MOAI22 U13730 ( .A1(n29093), .A2(n229), .B1(ram[560]), .B2(n230), .ZN(
        n4801) );
  MOAI22 U13731 ( .A1(n28858), .A2(n229), .B1(ram[561]), .B2(n230), .ZN(
        n4802) );
  MOAI22 U13732 ( .A1(n28623), .A2(n229), .B1(ram[562]), .B2(n230), .ZN(
        n4803) );
  MOAI22 U13733 ( .A1(n28388), .A2(n229), .B1(ram[563]), .B2(n230), .ZN(
        n4804) );
  MOAI22 U13734 ( .A1(n28153), .A2(n229), .B1(ram[564]), .B2(n230), .ZN(
        n4805) );
  MOAI22 U13735 ( .A1(n27918), .A2(n229), .B1(ram[565]), .B2(n230), .ZN(
        n4806) );
  MOAI22 U13736 ( .A1(n27683), .A2(n229), .B1(ram[566]), .B2(n230), .ZN(
        n4807) );
  MOAI22 U13737 ( .A1(n27448), .A2(n229), .B1(ram[567]), .B2(n230), .ZN(
        n4808) );
  MOAI22 U13738 ( .A1(n29093), .A2(n231), .B1(ram[568]), .B2(n232), .ZN(
        n4809) );
  MOAI22 U13739 ( .A1(n28858), .A2(n231), .B1(ram[569]), .B2(n232), .ZN(
        n4810) );
  MOAI22 U13740 ( .A1(n28623), .A2(n231), .B1(ram[570]), .B2(n232), .ZN(
        n4811) );
  MOAI22 U13741 ( .A1(n28388), .A2(n231), .B1(ram[571]), .B2(n232), .ZN(
        n4812) );
  MOAI22 U13742 ( .A1(n28153), .A2(n231), .B1(ram[572]), .B2(n232), .ZN(
        n4813) );
  MOAI22 U13743 ( .A1(n27918), .A2(n231), .B1(ram[573]), .B2(n232), .ZN(
        n4814) );
  MOAI22 U13744 ( .A1(n27683), .A2(n231), .B1(ram[574]), .B2(n232), .ZN(
        n4815) );
  MOAI22 U13745 ( .A1(n27448), .A2(n231), .B1(ram[575]), .B2(n232), .ZN(
        n4816) );
  MOAI22 U13746 ( .A1(n29093), .A2(n233), .B1(ram[576]), .B2(n234), .ZN(
        n4817) );
  MOAI22 U13747 ( .A1(n28858), .A2(n233), .B1(ram[577]), .B2(n234), .ZN(
        n4818) );
  MOAI22 U13748 ( .A1(n28623), .A2(n233), .B1(ram[578]), .B2(n234), .ZN(
        n4819) );
  MOAI22 U13749 ( .A1(n28388), .A2(n233), .B1(ram[579]), .B2(n234), .ZN(
        n4820) );
  MOAI22 U13750 ( .A1(n28153), .A2(n233), .B1(ram[580]), .B2(n234), .ZN(
        n4821) );
  MOAI22 U13751 ( .A1(n27918), .A2(n233), .B1(ram[581]), .B2(n234), .ZN(
        n4822) );
  MOAI22 U13752 ( .A1(n27683), .A2(n233), .B1(ram[582]), .B2(n234), .ZN(
        n4823) );
  MOAI22 U13753 ( .A1(n27448), .A2(n233), .B1(ram[583]), .B2(n234), .ZN(
        n4824) );
  MOAI22 U13754 ( .A1(n29093), .A2(n235), .B1(ram[584]), .B2(n236), .ZN(
        n4825) );
  MOAI22 U13755 ( .A1(n28858), .A2(n235), .B1(ram[585]), .B2(n236), .ZN(
        n4826) );
  MOAI22 U13756 ( .A1(n28623), .A2(n235), .B1(ram[586]), .B2(n236), .ZN(
        n4827) );
  MOAI22 U13757 ( .A1(n28388), .A2(n235), .B1(ram[587]), .B2(n236), .ZN(
        n4828) );
  MOAI22 U13758 ( .A1(n28153), .A2(n235), .B1(ram[588]), .B2(n236), .ZN(
        n4829) );
  MOAI22 U13759 ( .A1(n27918), .A2(n235), .B1(ram[589]), .B2(n236), .ZN(
        n4830) );
  MOAI22 U13760 ( .A1(n27683), .A2(n235), .B1(ram[590]), .B2(n236), .ZN(
        n4831) );
  MOAI22 U13761 ( .A1(n27448), .A2(n235), .B1(ram[591]), .B2(n236), .ZN(
        n4832) );
  MOAI22 U13762 ( .A1(n29093), .A2(n237), .B1(ram[592]), .B2(n238), .ZN(
        n4833) );
  MOAI22 U13763 ( .A1(n28858), .A2(n237), .B1(ram[593]), .B2(n238), .ZN(
        n4834) );
  MOAI22 U13764 ( .A1(n28623), .A2(n237), .B1(ram[594]), .B2(n238), .ZN(
        n4835) );
  MOAI22 U13765 ( .A1(n28388), .A2(n237), .B1(ram[595]), .B2(n238), .ZN(
        n4836) );
  MOAI22 U13766 ( .A1(n28153), .A2(n237), .B1(ram[596]), .B2(n238), .ZN(
        n4837) );
  MOAI22 U13767 ( .A1(n27918), .A2(n237), .B1(ram[597]), .B2(n238), .ZN(
        n4838) );
  MOAI22 U13768 ( .A1(n27683), .A2(n237), .B1(ram[598]), .B2(n238), .ZN(
        n4839) );
  MOAI22 U13769 ( .A1(n27448), .A2(n237), .B1(ram[599]), .B2(n238), .ZN(
        n4840) );
  MOAI22 U13770 ( .A1(n29093), .A2(n239), .B1(ram[600]), .B2(n240), .ZN(
        n4841) );
  MOAI22 U13771 ( .A1(n28858), .A2(n239), .B1(ram[601]), .B2(n240), .ZN(
        n4842) );
  MOAI22 U13772 ( .A1(n28623), .A2(n239), .B1(ram[602]), .B2(n240), .ZN(
        n4843) );
  MOAI22 U13773 ( .A1(n28388), .A2(n239), .B1(ram[603]), .B2(n240), .ZN(
        n4844) );
  MOAI22 U13774 ( .A1(n28153), .A2(n239), .B1(ram[604]), .B2(n240), .ZN(
        n4845) );
  MOAI22 U13775 ( .A1(n27918), .A2(n239), .B1(ram[605]), .B2(n240), .ZN(
        n4846) );
  MOAI22 U13776 ( .A1(n27683), .A2(n239), .B1(ram[606]), .B2(n240), .ZN(
        n4847) );
  MOAI22 U13777 ( .A1(n27448), .A2(n239), .B1(ram[607]), .B2(n240), .ZN(
        n4848) );
  MOAI22 U13778 ( .A1(n29093), .A2(n241), .B1(ram[608]), .B2(n242), .ZN(
        n4849) );
  MOAI22 U13779 ( .A1(n28858), .A2(n241), .B1(ram[609]), .B2(n242), .ZN(
        n4850) );
  MOAI22 U13780 ( .A1(n28623), .A2(n241), .B1(ram[610]), .B2(n242), .ZN(
        n4851) );
  MOAI22 U13781 ( .A1(n28388), .A2(n241), .B1(ram[611]), .B2(n242), .ZN(
        n4852) );
  MOAI22 U13782 ( .A1(n28153), .A2(n241), .B1(ram[612]), .B2(n242), .ZN(
        n4853) );
  MOAI22 U13783 ( .A1(n27918), .A2(n241), .B1(ram[613]), .B2(n242), .ZN(
        n4854) );
  MOAI22 U13784 ( .A1(n27683), .A2(n241), .B1(ram[614]), .B2(n242), .ZN(
        n4855) );
  MOAI22 U13785 ( .A1(n27448), .A2(n241), .B1(ram[615]), .B2(n242), .ZN(
        n4856) );
  MOAI22 U13786 ( .A1(n29093), .A2(n243), .B1(ram[616]), .B2(n244), .ZN(
        n4857) );
  MOAI22 U13787 ( .A1(n28858), .A2(n243), .B1(ram[617]), .B2(n244), .ZN(
        n4858) );
  MOAI22 U13788 ( .A1(n28623), .A2(n243), .B1(ram[618]), .B2(n244), .ZN(
        n4859) );
  MOAI22 U13789 ( .A1(n28388), .A2(n243), .B1(ram[619]), .B2(n244), .ZN(
        n4860) );
  MOAI22 U13790 ( .A1(n28153), .A2(n243), .B1(ram[620]), .B2(n244), .ZN(
        n4861) );
  MOAI22 U13791 ( .A1(n27918), .A2(n243), .B1(ram[621]), .B2(n244), .ZN(
        n4862) );
  MOAI22 U13792 ( .A1(n27683), .A2(n243), .B1(ram[622]), .B2(n244), .ZN(
        n4863) );
  MOAI22 U13793 ( .A1(n27448), .A2(n243), .B1(ram[623]), .B2(n244), .ZN(
        n4864) );
  MOAI22 U13794 ( .A1(n29094), .A2(n245), .B1(ram[624]), .B2(n246), .ZN(
        n4865) );
  MOAI22 U13795 ( .A1(n28859), .A2(n245), .B1(ram[625]), .B2(n246), .ZN(
        n4866) );
  MOAI22 U13796 ( .A1(n28624), .A2(n245), .B1(ram[626]), .B2(n246), .ZN(
        n4867) );
  MOAI22 U13797 ( .A1(n28389), .A2(n245), .B1(ram[627]), .B2(n246), .ZN(
        n4868) );
  MOAI22 U13798 ( .A1(n28154), .A2(n245), .B1(ram[628]), .B2(n246), .ZN(
        n4869) );
  MOAI22 U13799 ( .A1(n27919), .A2(n245), .B1(ram[629]), .B2(n246), .ZN(
        n4870) );
  MOAI22 U13800 ( .A1(n27684), .A2(n245), .B1(ram[630]), .B2(n246), .ZN(
        n4871) );
  MOAI22 U13801 ( .A1(n27449), .A2(n245), .B1(ram[631]), .B2(n246), .ZN(
        n4872) );
  MOAI22 U13802 ( .A1(n29094), .A2(n247), .B1(ram[632]), .B2(n248), .ZN(
        n4873) );
  MOAI22 U13803 ( .A1(n28859), .A2(n247), .B1(ram[633]), .B2(n248), .ZN(
        n4874) );
  MOAI22 U13804 ( .A1(n28624), .A2(n247), .B1(ram[634]), .B2(n248), .ZN(
        n4875) );
  MOAI22 U13805 ( .A1(n28389), .A2(n247), .B1(ram[635]), .B2(n248), .ZN(
        n4876) );
  MOAI22 U13806 ( .A1(n28154), .A2(n247), .B1(ram[636]), .B2(n248), .ZN(
        n4877) );
  MOAI22 U13807 ( .A1(n27919), .A2(n247), .B1(ram[637]), .B2(n248), .ZN(
        n4878) );
  MOAI22 U13808 ( .A1(n27684), .A2(n247), .B1(ram[638]), .B2(n248), .ZN(
        n4879) );
  MOAI22 U13809 ( .A1(n27449), .A2(n247), .B1(ram[639]), .B2(n248), .ZN(
        n4880) );
  MOAI22 U13810 ( .A1(n29094), .A2(n249), .B1(ram[640]), .B2(n250), .ZN(
        n4881) );
  MOAI22 U13811 ( .A1(n28859), .A2(n249), .B1(ram[641]), .B2(n250), .ZN(
        n4882) );
  MOAI22 U13812 ( .A1(n28624), .A2(n249), .B1(ram[642]), .B2(n250), .ZN(
        n4883) );
  MOAI22 U13813 ( .A1(n28389), .A2(n249), .B1(ram[643]), .B2(n250), .ZN(
        n4884) );
  MOAI22 U13814 ( .A1(n28154), .A2(n249), .B1(ram[644]), .B2(n250), .ZN(
        n4885) );
  MOAI22 U13815 ( .A1(n27919), .A2(n249), .B1(ram[645]), .B2(n250), .ZN(
        n4886) );
  MOAI22 U13816 ( .A1(n27684), .A2(n249), .B1(ram[646]), .B2(n250), .ZN(
        n4887) );
  MOAI22 U13817 ( .A1(n27449), .A2(n249), .B1(ram[647]), .B2(n250), .ZN(
        n4888) );
  MOAI22 U13818 ( .A1(n29094), .A2(n251), .B1(ram[648]), .B2(n252), .ZN(
        n4889) );
  MOAI22 U13819 ( .A1(n28859), .A2(n251), .B1(ram[649]), .B2(n252), .ZN(
        n4890) );
  MOAI22 U13820 ( .A1(n28624), .A2(n251), .B1(ram[650]), .B2(n252), .ZN(
        n4891) );
  MOAI22 U13821 ( .A1(n28389), .A2(n251), .B1(ram[651]), .B2(n252), .ZN(
        n4892) );
  MOAI22 U13822 ( .A1(n28154), .A2(n251), .B1(ram[652]), .B2(n252), .ZN(
        n4893) );
  MOAI22 U13823 ( .A1(n27919), .A2(n251), .B1(ram[653]), .B2(n252), .ZN(
        n4894) );
  MOAI22 U13824 ( .A1(n27684), .A2(n251), .B1(ram[654]), .B2(n252), .ZN(
        n4895) );
  MOAI22 U13825 ( .A1(n27449), .A2(n251), .B1(ram[655]), .B2(n252), .ZN(
        n4896) );
  MOAI22 U13826 ( .A1(n29094), .A2(n253), .B1(ram[656]), .B2(n254), .ZN(
        n4897) );
  MOAI22 U13827 ( .A1(n28859), .A2(n253), .B1(ram[657]), .B2(n254), .ZN(
        n4898) );
  MOAI22 U13828 ( .A1(n28624), .A2(n253), .B1(ram[658]), .B2(n254), .ZN(
        n4899) );
  MOAI22 U13829 ( .A1(n28389), .A2(n253), .B1(ram[659]), .B2(n254), .ZN(
        n4900) );
  MOAI22 U13830 ( .A1(n28154), .A2(n253), .B1(ram[660]), .B2(n254), .ZN(
        n4901) );
  MOAI22 U13831 ( .A1(n27919), .A2(n253), .B1(ram[661]), .B2(n254), .ZN(
        n4902) );
  MOAI22 U13832 ( .A1(n27684), .A2(n253), .B1(ram[662]), .B2(n254), .ZN(
        n4903) );
  MOAI22 U13833 ( .A1(n27449), .A2(n253), .B1(ram[663]), .B2(n254), .ZN(
        n4904) );
  MOAI22 U13834 ( .A1(n29094), .A2(n255), .B1(ram[664]), .B2(n256), .ZN(
        n4905) );
  MOAI22 U13835 ( .A1(n28859), .A2(n255), .B1(ram[665]), .B2(n256), .ZN(
        n4906) );
  MOAI22 U13836 ( .A1(n28624), .A2(n255), .B1(ram[666]), .B2(n256), .ZN(
        n4907) );
  MOAI22 U13837 ( .A1(n28389), .A2(n255), .B1(ram[667]), .B2(n256), .ZN(
        n4908) );
  MOAI22 U13838 ( .A1(n28154), .A2(n255), .B1(ram[668]), .B2(n256), .ZN(
        n4909) );
  MOAI22 U13839 ( .A1(n27919), .A2(n255), .B1(ram[669]), .B2(n256), .ZN(
        n4910) );
  MOAI22 U13840 ( .A1(n27684), .A2(n255), .B1(ram[670]), .B2(n256), .ZN(
        n4911) );
  MOAI22 U13841 ( .A1(n27449), .A2(n255), .B1(ram[671]), .B2(n256), .ZN(
        n4912) );
  MOAI22 U13842 ( .A1(n29094), .A2(n257), .B1(ram[672]), .B2(n258), .ZN(
        n4913) );
  MOAI22 U13843 ( .A1(n28859), .A2(n257), .B1(ram[673]), .B2(n258), .ZN(
        n4914) );
  MOAI22 U13844 ( .A1(n28624), .A2(n257), .B1(ram[674]), .B2(n258), .ZN(
        n4915) );
  MOAI22 U13845 ( .A1(n28389), .A2(n257), .B1(ram[675]), .B2(n258), .ZN(
        n4916) );
  MOAI22 U13846 ( .A1(n28154), .A2(n257), .B1(ram[676]), .B2(n258), .ZN(
        n4917) );
  MOAI22 U13847 ( .A1(n27919), .A2(n257), .B1(ram[677]), .B2(n258), .ZN(
        n4918) );
  MOAI22 U13848 ( .A1(n27684), .A2(n257), .B1(ram[678]), .B2(n258), .ZN(
        n4919) );
  MOAI22 U13849 ( .A1(n27449), .A2(n257), .B1(ram[679]), .B2(n258), .ZN(
        n4920) );
  MOAI22 U13850 ( .A1(n29094), .A2(n259), .B1(ram[680]), .B2(n260), .ZN(
        n4921) );
  MOAI22 U13851 ( .A1(n28859), .A2(n259), .B1(ram[681]), .B2(n260), .ZN(
        n4922) );
  MOAI22 U13852 ( .A1(n28624), .A2(n259), .B1(ram[682]), .B2(n260), .ZN(
        n4923) );
  MOAI22 U13853 ( .A1(n28389), .A2(n259), .B1(ram[683]), .B2(n260), .ZN(
        n4924) );
  MOAI22 U13854 ( .A1(n28154), .A2(n259), .B1(ram[684]), .B2(n260), .ZN(
        n4925) );
  MOAI22 U13855 ( .A1(n27919), .A2(n259), .B1(ram[685]), .B2(n260), .ZN(
        n4926) );
  MOAI22 U13856 ( .A1(n27684), .A2(n259), .B1(ram[686]), .B2(n260), .ZN(
        n4927) );
  MOAI22 U13857 ( .A1(n27449), .A2(n259), .B1(ram[687]), .B2(n260), .ZN(
        n4928) );
  MOAI22 U13858 ( .A1(n29094), .A2(n261), .B1(ram[688]), .B2(n262), .ZN(
        n4929) );
  MOAI22 U13859 ( .A1(n28859), .A2(n261), .B1(ram[689]), .B2(n262), .ZN(
        n4930) );
  MOAI22 U13860 ( .A1(n28624), .A2(n261), .B1(ram[690]), .B2(n262), .ZN(
        n4931) );
  MOAI22 U13861 ( .A1(n28389), .A2(n261), .B1(ram[691]), .B2(n262), .ZN(
        n4932) );
  MOAI22 U13862 ( .A1(n28154), .A2(n261), .B1(ram[692]), .B2(n262), .ZN(
        n4933) );
  MOAI22 U13863 ( .A1(n27919), .A2(n261), .B1(ram[693]), .B2(n262), .ZN(
        n4934) );
  MOAI22 U13864 ( .A1(n27684), .A2(n261), .B1(ram[694]), .B2(n262), .ZN(
        n4935) );
  MOAI22 U13865 ( .A1(n27449), .A2(n261), .B1(ram[695]), .B2(n262), .ZN(
        n4936) );
  MOAI22 U13866 ( .A1(n29094), .A2(n263), .B1(ram[696]), .B2(n264), .ZN(
        n4937) );
  MOAI22 U13867 ( .A1(n28859), .A2(n263), .B1(ram[697]), .B2(n264), .ZN(
        n4938) );
  MOAI22 U13868 ( .A1(n28624), .A2(n263), .B1(ram[698]), .B2(n264), .ZN(
        n4939) );
  MOAI22 U13869 ( .A1(n28389), .A2(n263), .B1(ram[699]), .B2(n264), .ZN(
        n4940) );
  MOAI22 U13870 ( .A1(n28154), .A2(n263), .B1(ram[700]), .B2(n264), .ZN(
        n4941) );
  MOAI22 U13871 ( .A1(n27919), .A2(n263), .B1(ram[701]), .B2(n264), .ZN(
        n4942) );
  MOAI22 U13872 ( .A1(n27684), .A2(n263), .B1(ram[702]), .B2(n264), .ZN(
        n4943) );
  MOAI22 U13873 ( .A1(n27449), .A2(n263), .B1(ram[703]), .B2(n264), .ZN(
        n4944) );
  MOAI22 U13874 ( .A1(n29094), .A2(n265), .B1(ram[704]), .B2(n266), .ZN(
        n4945) );
  MOAI22 U13875 ( .A1(n28859), .A2(n265), .B1(ram[705]), .B2(n266), .ZN(
        n4946) );
  MOAI22 U13876 ( .A1(n28624), .A2(n265), .B1(ram[706]), .B2(n266), .ZN(
        n4947) );
  MOAI22 U13877 ( .A1(n28389), .A2(n265), .B1(ram[707]), .B2(n266), .ZN(
        n4948) );
  MOAI22 U13878 ( .A1(n28154), .A2(n265), .B1(ram[708]), .B2(n266), .ZN(
        n4949) );
  MOAI22 U13879 ( .A1(n27919), .A2(n265), .B1(ram[709]), .B2(n266), .ZN(
        n4950) );
  MOAI22 U13880 ( .A1(n27684), .A2(n265), .B1(ram[710]), .B2(n266), .ZN(
        n4951) );
  MOAI22 U13881 ( .A1(n27449), .A2(n265), .B1(ram[711]), .B2(n266), .ZN(
        n4952) );
  MOAI22 U13882 ( .A1(n29094), .A2(n267), .B1(ram[712]), .B2(n268), .ZN(
        n4953) );
  MOAI22 U13883 ( .A1(n28859), .A2(n267), .B1(ram[713]), .B2(n268), .ZN(
        n4954) );
  MOAI22 U13884 ( .A1(n28624), .A2(n267), .B1(ram[714]), .B2(n268), .ZN(
        n4955) );
  MOAI22 U13885 ( .A1(n28389), .A2(n267), .B1(ram[715]), .B2(n268), .ZN(
        n4956) );
  MOAI22 U13886 ( .A1(n28154), .A2(n267), .B1(ram[716]), .B2(n268), .ZN(
        n4957) );
  MOAI22 U13887 ( .A1(n27919), .A2(n267), .B1(ram[717]), .B2(n268), .ZN(
        n4958) );
  MOAI22 U13888 ( .A1(n27684), .A2(n267), .B1(ram[718]), .B2(n268), .ZN(
        n4959) );
  MOAI22 U13889 ( .A1(n27449), .A2(n267), .B1(ram[719]), .B2(n268), .ZN(
        n4960) );
  MOAI22 U13890 ( .A1(n29094), .A2(n269), .B1(ram[720]), .B2(n270), .ZN(
        n4961) );
  MOAI22 U13891 ( .A1(n28859), .A2(n269), .B1(ram[721]), .B2(n270), .ZN(
        n4962) );
  MOAI22 U13892 ( .A1(n28624), .A2(n269), .B1(ram[722]), .B2(n270), .ZN(
        n4963) );
  MOAI22 U13893 ( .A1(n28389), .A2(n269), .B1(ram[723]), .B2(n270), .ZN(
        n4964) );
  MOAI22 U13894 ( .A1(n28154), .A2(n269), .B1(ram[724]), .B2(n270), .ZN(
        n4965) );
  MOAI22 U13895 ( .A1(n27919), .A2(n269), .B1(ram[725]), .B2(n270), .ZN(
        n4966) );
  MOAI22 U13896 ( .A1(n27684), .A2(n269), .B1(ram[726]), .B2(n270), .ZN(
        n4967) );
  MOAI22 U13897 ( .A1(n27449), .A2(n269), .B1(ram[727]), .B2(n270), .ZN(
        n4968) );
  MOAI22 U13898 ( .A1(n29095), .A2(n271), .B1(ram[728]), .B2(n272), .ZN(
        n4969) );
  MOAI22 U13899 ( .A1(n28860), .A2(n271), .B1(ram[729]), .B2(n272), .ZN(
        n4970) );
  MOAI22 U13900 ( .A1(n28625), .A2(n271), .B1(ram[730]), .B2(n272), .ZN(
        n4971) );
  MOAI22 U13901 ( .A1(n28390), .A2(n271), .B1(ram[731]), .B2(n272), .ZN(
        n4972) );
  MOAI22 U13902 ( .A1(n28155), .A2(n271), .B1(ram[732]), .B2(n272), .ZN(
        n4973) );
  MOAI22 U13903 ( .A1(n27920), .A2(n271), .B1(ram[733]), .B2(n272), .ZN(
        n4974) );
  MOAI22 U13904 ( .A1(n27685), .A2(n271), .B1(ram[734]), .B2(n272), .ZN(
        n4975) );
  MOAI22 U13905 ( .A1(n27450), .A2(n271), .B1(ram[735]), .B2(n272), .ZN(
        n4976) );
  MOAI22 U13906 ( .A1(n29095), .A2(n273), .B1(ram[736]), .B2(n274), .ZN(
        n4977) );
  MOAI22 U13907 ( .A1(n28860), .A2(n273), .B1(ram[737]), .B2(n274), .ZN(
        n4978) );
  MOAI22 U13908 ( .A1(n28625), .A2(n273), .B1(ram[738]), .B2(n274), .ZN(
        n4979) );
  MOAI22 U13909 ( .A1(n28390), .A2(n273), .B1(ram[739]), .B2(n274), .ZN(
        n4980) );
  MOAI22 U13910 ( .A1(n28155), .A2(n273), .B1(ram[740]), .B2(n274), .ZN(
        n4981) );
  MOAI22 U13911 ( .A1(n27920), .A2(n273), .B1(ram[741]), .B2(n274), .ZN(
        n4982) );
  MOAI22 U13912 ( .A1(n27685), .A2(n273), .B1(ram[742]), .B2(n274), .ZN(
        n4983) );
  MOAI22 U13913 ( .A1(n27450), .A2(n273), .B1(ram[743]), .B2(n274), .ZN(
        n4984) );
  MOAI22 U13914 ( .A1(n29095), .A2(n275), .B1(ram[744]), .B2(n276), .ZN(
        n4985) );
  MOAI22 U13915 ( .A1(n28860), .A2(n275), .B1(ram[745]), .B2(n276), .ZN(
        n4986) );
  MOAI22 U13916 ( .A1(n28625), .A2(n275), .B1(ram[746]), .B2(n276), .ZN(
        n4987) );
  MOAI22 U13917 ( .A1(n28390), .A2(n275), .B1(ram[747]), .B2(n276), .ZN(
        n4988) );
  MOAI22 U13918 ( .A1(n28155), .A2(n275), .B1(ram[748]), .B2(n276), .ZN(
        n4989) );
  MOAI22 U13919 ( .A1(n27920), .A2(n275), .B1(ram[749]), .B2(n276), .ZN(
        n4990) );
  MOAI22 U13920 ( .A1(n27685), .A2(n275), .B1(ram[750]), .B2(n276), .ZN(
        n4991) );
  MOAI22 U13921 ( .A1(n27450), .A2(n275), .B1(ram[751]), .B2(n276), .ZN(
        n4992) );
  MOAI22 U13922 ( .A1(n29095), .A2(n277), .B1(ram[752]), .B2(n278), .ZN(
        n4993) );
  MOAI22 U13923 ( .A1(n28860), .A2(n277), .B1(ram[753]), .B2(n278), .ZN(
        n4994) );
  MOAI22 U13924 ( .A1(n28625), .A2(n277), .B1(ram[754]), .B2(n278), .ZN(
        n4995) );
  MOAI22 U13925 ( .A1(n28390), .A2(n277), .B1(ram[755]), .B2(n278), .ZN(
        n4996) );
  MOAI22 U13926 ( .A1(n28155), .A2(n277), .B1(ram[756]), .B2(n278), .ZN(
        n4997) );
  MOAI22 U13927 ( .A1(n27920), .A2(n277), .B1(ram[757]), .B2(n278), .ZN(
        n4998) );
  MOAI22 U13928 ( .A1(n27685), .A2(n277), .B1(ram[758]), .B2(n278), .ZN(
        n4999) );
  MOAI22 U13929 ( .A1(n27450), .A2(n277), .B1(ram[759]), .B2(n278), .ZN(
        n5000) );
  MOAI22 U13930 ( .A1(n29095), .A2(n279), .B1(ram[760]), .B2(n280), .ZN(
        n5001) );
  MOAI22 U13931 ( .A1(n28860), .A2(n279), .B1(ram[761]), .B2(n280), .ZN(
        n5002) );
  MOAI22 U13932 ( .A1(n28625), .A2(n279), .B1(ram[762]), .B2(n280), .ZN(
        n5003) );
  MOAI22 U13933 ( .A1(n28390), .A2(n279), .B1(ram[763]), .B2(n280), .ZN(
        n5004) );
  MOAI22 U13934 ( .A1(n28155), .A2(n279), .B1(ram[764]), .B2(n280), .ZN(
        n5005) );
  MOAI22 U13935 ( .A1(n27920), .A2(n279), .B1(ram[765]), .B2(n280), .ZN(
        n5006) );
  MOAI22 U13936 ( .A1(n27685), .A2(n279), .B1(ram[766]), .B2(n280), .ZN(
        n5007) );
  MOAI22 U13937 ( .A1(n27450), .A2(n279), .B1(ram[767]), .B2(n280), .ZN(
        n5008) );
  MOAI22 U13938 ( .A1(n29095), .A2(n281), .B1(ram[768]), .B2(n282), .ZN(
        n5009) );
  MOAI22 U13939 ( .A1(n28860), .A2(n281), .B1(ram[769]), .B2(n282), .ZN(
        n5010) );
  MOAI22 U13940 ( .A1(n28625), .A2(n281), .B1(ram[770]), .B2(n282), .ZN(
        n5011) );
  MOAI22 U13941 ( .A1(n28390), .A2(n281), .B1(ram[771]), .B2(n282), .ZN(
        n5012) );
  MOAI22 U13942 ( .A1(n28155), .A2(n281), .B1(ram[772]), .B2(n282), .ZN(
        n5013) );
  MOAI22 U13943 ( .A1(n27920), .A2(n281), .B1(ram[773]), .B2(n282), .ZN(
        n5014) );
  MOAI22 U13944 ( .A1(n27685), .A2(n281), .B1(ram[774]), .B2(n282), .ZN(
        n5015) );
  MOAI22 U13945 ( .A1(n27450), .A2(n281), .B1(ram[775]), .B2(n282), .ZN(
        n5016) );
  MOAI22 U13946 ( .A1(n29095), .A2(n283), .B1(ram[776]), .B2(n284), .ZN(
        n5017) );
  MOAI22 U13947 ( .A1(n28860), .A2(n283), .B1(ram[777]), .B2(n284), .ZN(
        n5018) );
  MOAI22 U13948 ( .A1(n28625), .A2(n283), .B1(ram[778]), .B2(n284), .ZN(
        n5019) );
  MOAI22 U13949 ( .A1(n28390), .A2(n283), .B1(ram[779]), .B2(n284), .ZN(
        n5020) );
  MOAI22 U13950 ( .A1(n28155), .A2(n283), .B1(ram[780]), .B2(n284), .ZN(
        n5021) );
  MOAI22 U13951 ( .A1(n27920), .A2(n283), .B1(ram[781]), .B2(n284), .ZN(
        n5022) );
  MOAI22 U13952 ( .A1(n27685), .A2(n283), .B1(ram[782]), .B2(n284), .ZN(
        n5023) );
  MOAI22 U13953 ( .A1(n27450), .A2(n283), .B1(ram[783]), .B2(n284), .ZN(
        n5024) );
  MOAI22 U13954 ( .A1(n29095), .A2(n285), .B1(ram[784]), .B2(n286), .ZN(
        n5025) );
  MOAI22 U13955 ( .A1(n28860), .A2(n285), .B1(ram[785]), .B2(n286), .ZN(
        n5026) );
  MOAI22 U13956 ( .A1(n28625), .A2(n285), .B1(ram[786]), .B2(n286), .ZN(
        n5027) );
  MOAI22 U13957 ( .A1(n28390), .A2(n285), .B1(ram[787]), .B2(n286), .ZN(
        n5028) );
  MOAI22 U13958 ( .A1(n28155), .A2(n285), .B1(ram[788]), .B2(n286), .ZN(
        n5029) );
  MOAI22 U13959 ( .A1(n27920), .A2(n285), .B1(ram[789]), .B2(n286), .ZN(
        n5030) );
  MOAI22 U13960 ( .A1(n27685), .A2(n285), .B1(ram[790]), .B2(n286), .ZN(
        n5031) );
  MOAI22 U13961 ( .A1(n27450), .A2(n285), .B1(ram[791]), .B2(n286), .ZN(
        n5032) );
  MOAI22 U13962 ( .A1(n29095), .A2(n287), .B1(ram[792]), .B2(n288), .ZN(
        n5033) );
  MOAI22 U13963 ( .A1(n28860), .A2(n287), .B1(ram[793]), .B2(n288), .ZN(
        n5034) );
  MOAI22 U13964 ( .A1(n28625), .A2(n287), .B1(ram[794]), .B2(n288), .ZN(
        n5035) );
  MOAI22 U13965 ( .A1(n28390), .A2(n287), .B1(ram[795]), .B2(n288), .ZN(
        n5036) );
  MOAI22 U13966 ( .A1(n28155), .A2(n287), .B1(ram[796]), .B2(n288), .ZN(
        n5037) );
  MOAI22 U13967 ( .A1(n27920), .A2(n287), .B1(ram[797]), .B2(n288), .ZN(
        n5038) );
  MOAI22 U13968 ( .A1(n27685), .A2(n287), .B1(ram[798]), .B2(n288), .ZN(
        n5039) );
  MOAI22 U13969 ( .A1(n27450), .A2(n287), .B1(ram[799]), .B2(n288), .ZN(
        n5040) );
  MOAI22 U13970 ( .A1(n29095), .A2(n289), .B1(ram[800]), .B2(n290), .ZN(
        n5041) );
  MOAI22 U13971 ( .A1(n28860), .A2(n289), .B1(ram[801]), .B2(n290), .ZN(
        n5042) );
  MOAI22 U13972 ( .A1(n28625), .A2(n289), .B1(ram[802]), .B2(n290), .ZN(
        n5043) );
  MOAI22 U13973 ( .A1(n28390), .A2(n289), .B1(ram[803]), .B2(n290), .ZN(
        n5044) );
  MOAI22 U13974 ( .A1(n28155), .A2(n289), .B1(ram[804]), .B2(n290), .ZN(
        n5045) );
  MOAI22 U13975 ( .A1(n27920), .A2(n289), .B1(ram[805]), .B2(n290), .ZN(
        n5046) );
  MOAI22 U13976 ( .A1(n27685), .A2(n289), .B1(ram[806]), .B2(n290), .ZN(
        n5047) );
  MOAI22 U13977 ( .A1(n27450), .A2(n289), .B1(ram[807]), .B2(n290), .ZN(
        n5048) );
  MOAI22 U13978 ( .A1(n29095), .A2(n291), .B1(ram[808]), .B2(n292), .ZN(
        n5049) );
  MOAI22 U13979 ( .A1(n28860), .A2(n291), .B1(ram[809]), .B2(n292), .ZN(
        n5050) );
  MOAI22 U13980 ( .A1(n28625), .A2(n291), .B1(ram[810]), .B2(n292), .ZN(
        n5051) );
  MOAI22 U13981 ( .A1(n28390), .A2(n291), .B1(ram[811]), .B2(n292), .ZN(
        n5052) );
  MOAI22 U13982 ( .A1(n28155), .A2(n291), .B1(ram[812]), .B2(n292), .ZN(
        n5053) );
  MOAI22 U13983 ( .A1(n27920), .A2(n291), .B1(ram[813]), .B2(n292), .ZN(
        n5054) );
  MOAI22 U13984 ( .A1(n27685), .A2(n291), .B1(ram[814]), .B2(n292), .ZN(
        n5055) );
  MOAI22 U13985 ( .A1(n27450), .A2(n291), .B1(ram[815]), .B2(n292), .ZN(
        n5056) );
  MOAI22 U13986 ( .A1(n29095), .A2(n293), .B1(ram[816]), .B2(n294), .ZN(
        n5057) );
  MOAI22 U13987 ( .A1(n28860), .A2(n293), .B1(ram[817]), .B2(n294), .ZN(
        n5058) );
  MOAI22 U13988 ( .A1(n28625), .A2(n293), .B1(ram[818]), .B2(n294), .ZN(
        n5059) );
  MOAI22 U13989 ( .A1(n28390), .A2(n293), .B1(ram[819]), .B2(n294), .ZN(
        n5060) );
  MOAI22 U13990 ( .A1(n28155), .A2(n293), .B1(ram[820]), .B2(n294), .ZN(
        n5061) );
  MOAI22 U13991 ( .A1(n27920), .A2(n293), .B1(ram[821]), .B2(n294), .ZN(
        n5062) );
  MOAI22 U13992 ( .A1(n27685), .A2(n293), .B1(ram[822]), .B2(n294), .ZN(
        n5063) );
  MOAI22 U13993 ( .A1(n27450), .A2(n293), .B1(ram[823]), .B2(n294), .ZN(
        n5064) );
  MOAI22 U13994 ( .A1(n29095), .A2(n295), .B1(ram[824]), .B2(n296), .ZN(
        n5065) );
  MOAI22 U13995 ( .A1(n28860), .A2(n295), .B1(ram[825]), .B2(n296), .ZN(
        n5066) );
  MOAI22 U13996 ( .A1(n28625), .A2(n295), .B1(ram[826]), .B2(n296), .ZN(
        n5067) );
  MOAI22 U13997 ( .A1(n28390), .A2(n295), .B1(ram[827]), .B2(n296), .ZN(
        n5068) );
  MOAI22 U13998 ( .A1(n28155), .A2(n295), .B1(ram[828]), .B2(n296), .ZN(
        n5069) );
  MOAI22 U13999 ( .A1(n27920), .A2(n295), .B1(ram[829]), .B2(n296), .ZN(
        n5070) );
  MOAI22 U14000 ( .A1(n27685), .A2(n295), .B1(ram[830]), .B2(n296), .ZN(
        n5071) );
  MOAI22 U14001 ( .A1(n27450), .A2(n295), .B1(ram[831]), .B2(n296), .ZN(
        n5072) );
  MOAI22 U14002 ( .A1(n29096), .A2(n297), .B1(ram[832]), .B2(n298), .ZN(
        n5073) );
  MOAI22 U14003 ( .A1(n28861), .A2(n297), .B1(ram[833]), .B2(n298), .ZN(
        n5074) );
  MOAI22 U14004 ( .A1(n28626), .A2(n297), .B1(ram[834]), .B2(n298), .ZN(
        n5075) );
  MOAI22 U14005 ( .A1(n28391), .A2(n297), .B1(ram[835]), .B2(n298), .ZN(
        n5076) );
  MOAI22 U14006 ( .A1(n28156), .A2(n297), .B1(ram[836]), .B2(n298), .ZN(
        n5077) );
  MOAI22 U14007 ( .A1(n27921), .A2(n297), .B1(ram[837]), .B2(n298), .ZN(
        n5078) );
  MOAI22 U14008 ( .A1(n27686), .A2(n297), .B1(ram[838]), .B2(n298), .ZN(
        n5079) );
  MOAI22 U14009 ( .A1(n27451), .A2(n297), .B1(ram[839]), .B2(n298), .ZN(
        n5080) );
  MOAI22 U14010 ( .A1(n29096), .A2(n299), .B1(ram[840]), .B2(n300), .ZN(
        n5081) );
  MOAI22 U14011 ( .A1(n28861), .A2(n299), .B1(ram[841]), .B2(n300), .ZN(
        n5082) );
  MOAI22 U14012 ( .A1(n28626), .A2(n299), .B1(ram[842]), .B2(n300), .ZN(
        n5083) );
  MOAI22 U14013 ( .A1(n28391), .A2(n299), .B1(ram[843]), .B2(n300), .ZN(
        n5084) );
  MOAI22 U14014 ( .A1(n28156), .A2(n299), .B1(ram[844]), .B2(n300), .ZN(
        n5085) );
  MOAI22 U14015 ( .A1(n27921), .A2(n299), .B1(ram[845]), .B2(n300), .ZN(
        n5086) );
  MOAI22 U14016 ( .A1(n27686), .A2(n299), .B1(ram[846]), .B2(n300), .ZN(
        n5087) );
  MOAI22 U14017 ( .A1(n27451), .A2(n299), .B1(ram[847]), .B2(n300), .ZN(
        n5088) );
  MOAI22 U14018 ( .A1(n29096), .A2(n301), .B1(ram[848]), .B2(n302), .ZN(
        n5089) );
  MOAI22 U14019 ( .A1(n28861), .A2(n301), .B1(ram[849]), .B2(n302), .ZN(
        n5090) );
  MOAI22 U14020 ( .A1(n28626), .A2(n301), .B1(ram[850]), .B2(n302), .ZN(
        n5091) );
  MOAI22 U14021 ( .A1(n28391), .A2(n301), .B1(ram[851]), .B2(n302), .ZN(
        n5092) );
  MOAI22 U14022 ( .A1(n28156), .A2(n301), .B1(ram[852]), .B2(n302), .ZN(
        n5093) );
  MOAI22 U14023 ( .A1(n27921), .A2(n301), .B1(ram[853]), .B2(n302), .ZN(
        n5094) );
  MOAI22 U14024 ( .A1(n27686), .A2(n301), .B1(ram[854]), .B2(n302), .ZN(
        n5095) );
  MOAI22 U14025 ( .A1(n27451), .A2(n301), .B1(ram[855]), .B2(n302), .ZN(
        n5096) );
  MOAI22 U14026 ( .A1(n29096), .A2(n303), .B1(ram[856]), .B2(n304), .ZN(
        n5097) );
  MOAI22 U14027 ( .A1(n28861), .A2(n303), .B1(ram[857]), .B2(n304), .ZN(
        n5098) );
  MOAI22 U14028 ( .A1(n28626), .A2(n303), .B1(ram[858]), .B2(n304), .ZN(
        n5099) );
  MOAI22 U14029 ( .A1(n28391), .A2(n303), .B1(ram[859]), .B2(n304), .ZN(
        n5100) );
  MOAI22 U14030 ( .A1(n28156), .A2(n303), .B1(ram[860]), .B2(n304), .ZN(
        n5101) );
  MOAI22 U14031 ( .A1(n27921), .A2(n303), .B1(ram[861]), .B2(n304), .ZN(
        n5102) );
  MOAI22 U14032 ( .A1(n27686), .A2(n303), .B1(ram[862]), .B2(n304), .ZN(
        n5103) );
  MOAI22 U14033 ( .A1(n27451), .A2(n303), .B1(ram[863]), .B2(n304), .ZN(
        n5104) );
  MOAI22 U14034 ( .A1(n29096), .A2(n305), .B1(ram[864]), .B2(n306), .ZN(
        n5105) );
  MOAI22 U14035 ( .A1(n28861), .A2(n305), .B1(ram[865]), .B2(n306), .ZN(
        n5106) );
  MOAI22 U14036 ( .A1(n28626), .A2(n305), .B1(ram[866]), .B2(n306), .ZN(
        n5107) );
  MOAI22 U14037 ( .A1(n28391), .A2(n305), .B1(ram[867]), .B2(n306), .ZN(
        n5108) );
  MOAI22 U14038 ( .A1(n28156), .A2(n305), .B1(ram[868]), .B2(n306), .ZN(
        n5109) );
  MOAI22 U14039 ( .A1(n27921), .A2(n305), .B1(ram[869]), .B2(n306), .ZN(
        n5110) );
  MOAI22 U14040 ( .A1(n27686), .A2(n305), .B1(ram[870]), .B2(n306), .ZN(
        n5111) );
  MOAI22 U14041 ( .A1(n27451), .A2(n305), .B1(ram[871]), .B2(n306), .ZN(
        n5112) );
  MOAI22 U14042 ( .A1(n29096), .A2(n307), .B1(ram[872]), .B2(n308), .ZN(
        n5113) );
  MOAI22 U14043 ( .A1(n28861), .A2(n307), .B1(ram[873]), .B2(n308), .ZN(
        n5114) );
  MOAI22 U14044 ( .A1(n28626), .A2(n307), .B1(ram[874]), .B2(n308), .ZN(
        n5115) );
  MOAI22 U14045 ( .A1(n28391), .A2(n307), .B1(ram[875]), .B2(n308), .ZN(
        n5116) );
  MOAI22 U14046 ( .A1(n28156), .A2(n307), .B1(ram[876]), .B2(n308), .ZN(
        n5117) );
  MOAI22 U14047 ( .A1(n27921), .A2(n307), .B1(ram[877]), .B2(n308), .ZN(
        n5118) );
  MOAI22 U14048 ( .A1(n27686), .A2(n307), .B1(ram[878]), .B2(n308), .ZN(
        n5119) );
  MOAI22 U14049 ( .A1(n27451), .A2(n307), .B1(ram[879]), .B2(n308), .ZN(
        n5120) );
  MOAI22 U14050 ( .A1(n29096), .A2(n309), .B1(ram[880]), .B2(n310), .ZN(
        n5121) );
  MOAI22 U14051 ( .A1(n28861), .A2(n309), .B1(ram[881]), .B2(n310), .ZN(
        n5122) );
  MOAI22 U14052 ( .A1(n28626), .A2(n309), .B1(ram[882]), .B2(n310), .ZN(
        n5123) );
  MOAI22 U14053 ( .A1(n28391), .A2(n309), .B1(ram[883]), .B2(n310), .ZN(
        n5124) );
  MOAI22 U14054 ( .A1(n28156), .A2(n309), .B1(ram[884]), .B2(n310), .ZN(
        n5125) );
  MOAI22 U14055 ( .A1(n27921), .A2(n309), .B1(ram[885]), .B2(n310), .ZN(
        n5126) );
  MOAI22 U14056 ( .A1(n27686), .A2(n309), .B1(ram[886]), .B2(n310), .ZN(
        n5127) );
  MOAI22 U14057 ( .A1(n27451), .A2(n309), .B1(ram[887]), .B2(n310), .ZN(
        n5128) );
  MOAI22 U14058 ( .A1(n29096), .A2(n311), .B1(ram[888]), .B2(n312), .ZN(
        n5129) );
  MOAI22 U14059 ( .A1(n28861), .A2(n311), .B1(ram[889]), .B2(n312), .ZN(
        n5130) );
  MOAI22 U14060 ( .A1(n28626), .A2(n311), .B1(ram[890]), .B2(n312), .ZN(
        n5131) );
  MOAI22 U14061 ( .A1(n28391), .A2(n311), .B1(ram[891]), .B2(n312), .ZN(
        n5132) );
  MOAI22 U14062 ( .A1(n28156), .A2(n311), .B1(ram[892]), .B2(n312), .ZN(
        n5133) );
  MOAI22 U14063 ( .A1(n27921), .A2(n311), .B1(ram[893]), .B2(n312), .ZN(
        n5134) );
  MOAI22 U14064 ( .A1(n27686), .A2(n311), .B1(ram[894]), .B2(n312), .ZN(
        n5135) );
  MOAI22 U14065 ( .A1(n27451), .A2(n311), .B1(ram[895]), .B2(n312), .ZN(
        n5136) );
  MOAI22 U14066 ( .A1(n29096), .A2(n313), .B1(ram[896]), .B2(n314), .ZN(
        n5137) );
  MOAI22 U14067 ( .A1(n28861), .A2(n313), .B1(ram[897]), .B2(n314), .ZN(
        n5138) );
  MOAI22 U14068 ( .A1(n28626), .A2(n313), .B1(ram[898]), .B2(n314), .ZN(
        n5139) );
  MOAI22 U14069 ( .A1(n28391), .A2(n313), .B1(ram[899]), .B2(n314), .ZN(
        n5140) );
  MOAI22 U14070 ( .A1(n28156), .A2(n313), .B1(ram[900]), .B2(n314), .ZN(
        n5141) );
  MOAI22 U14071 ( .A1(n27921), .A2(n313), .B1(ram[901]), .B2(n314), .ZN(
        n5142) );
  MOAI22 U14072 ( .A1(n27686), .A2(n313), .B1(ram[902]), .B2(n314), .ZN(
        n5143) );
  MOAI22 U14073 ( .A1(n27451), .A2(n313), .B1(ram[903]), .B2(n314), .ZN(
        n5144) );
  MOAI22 U14074 ( .A1(n29096), .A2(n315), .B1(ram[904]), .B2(n316), .ZN(
        n5145) );
  MOAI22 U14075 ( .A1(n28861), .A2(n315), .B1(ram[905]), .B2(n316), .ZN(
        n5146) );
  MOAI22 U14076 ( .A1(n28626), .A2(n315), .B1(ram[906]), .B2(n316), .ZN(
        n5147) );
  MOAI22 U14077 ( .A1(n28391), .A2(n315), .B1(ram[907]), .B2(n316), .ZN(
        n5148) );
  MOAI22 U14078 ( .A1(n28156), .A2(n315), .B1(ram[908]), .B2(n316), .ZN(
        n5149) );
  MOAI22 U14079 ( .A1(n27921), .A2(n315), .B1(ram[909]), .B2(n316), .ZN(
        n5150) );
  MOAI22 U14080 ( .A1(n27686), .A2(n315), .B1(ram[910]), .B2(n316), .ZN(
        n5151) );
  MOAI22 U14081 ( .A1(n27451), .A2(n315), .B1(ram[911]), .B2(n316), .ZN(
        n5152) );
  MOAI22 U14082 ( .A1(n29096), .A2(n317), .B1(ram[912]), .B2(n318), .ZN(
        n5153) );
  MOAI22 U14083 ( .A1(n28861), .A2(n317), .B1(ram[913]), .B2(n318), .ZN(
        n5154) );
  MOAI22 U14084 ( .A1(n28626), .A2(n317), .B1(ram[914]), .B2(n318), .ZN(
        n5155) );
  MOAI22 U14085 ( .A1(n28391), .A2(n317), .B1(ram[915]), .B2(n318), .ZN(
        n5156) );
  MOAI22 U14086 ( .A1(n28156), .A2(n317), .B1(ram[916]), .B2(n318), .ZN(
        n5157) );
  MOAI22 U14087 ( .A1(n27921), .A2(n317), .B1(ram[917]), .B2(n318), .ZN(
        n5158) );
  MOAI22 U14088 ( .A1(n27686), .A2(n317), .B1(ram[918]), .B2(n318), .ZN(
        n5159) );
  MOAI22 U14089 ( .A1(n27451), .A2(n317), .B1(ram[919]), .B2(n318), .ZN(
        n5160) );
  MOAI22 U14090 ( .A1(n29096), .A2(n319), .B1(ram[920]), .B2(n320), .ZN(
        n5161) );
  MOAI22 U14091 ( .A1(n28861), .A2(n319), .B1(ram[921]), .B2(n320), .ZN(
        n5162) );
  MOAI22 U14092 ( .A1(n28626), .A2(n319), .B1(ram[922]), .B2(n320), .ZN(
        n5163) );
  MOAI22 U14093 ( .A1(n28391), .A2(n319), .B1(ram[923]), .B2(n320), .ZN(
        n5164) );
  MOAI22 U14094 ( .A1(n28156), .A2(n319), .B1(ram[924]), .B2(n320), .ZN(
        n5165) );
  MOAI22 U14095 ( .A1(n27921), .A2(n319), .B1(ram[925]), .B2(n320), .ZN(
        n5166) );
  MOAI22 U14096 ( .A1(n27686), .A2(n319), .B1(ram[926]), .B2(n320), .ZN(
        n5167) );
  MOAI22 U14097 ( .A1(n27451), .A2(n319), .B1(ram[927]), .B2(n320), .ZN(
        n5168) );
  MOAI22 U14098 ( .A1(n29096), .A2(n321), .B1(ram[928]), .B2(n322), .ZN(
        n5169) );
  MOAI22 U14099 ( .A1(n28861), .A2(n321), .B1(ram[929]), .B2(n322), .ZN(
        n5170) );
  MOAI22 U14100 ( .A1(n28626), .A2(n321), .B1(ram[930]), .B2(n322), .ZN(
        n5171) );
  MOAI22 U14101 ( .A1(n28391), .A2(n321), .B1(ram[931]), .B2(n322), .ZN(
        n5172) );
  MOAI22 U14102 ( .A1(n28156), .A2(n321), .B1(ram[932]), .B2(n322), .ZN(
        n5173) );
  MOAI22 U14103 ( .A1(n27921), .A2(n321), .B1(ram[933]), .B2(n322), .ZN(
        n5174) );
  MOAI22 U14104 ( .A1(n27686), .A2(n321), .B1(ram[934]), .B2(n322), .ZN(
        n5175) );
  MOAI22 U14105 ( .A1(n27451), .A2(n321), .B1(ram[935]), .B2(n322), .ZN(
        n5176) );
  MOAI22 U14106 ( .A1(n29097), .A2(n323), .B1(ram[936]), .B2(n324), .ZN(
        n5177) );
  MOAI22 U14107 ( .A1(n28862), .A2(n323), .B1(ram[937]), .B2(n324), .ZN(
        n5178) );
  MOAI22 U14108 ( .A1(n28627), .A2(n323), .B1(ram[938]), .B2(n324), .ZN(
        n5179) );
  MOAI22 U14109 ( .A1(n28392), .A2(n323), .B1(ram[939]), .B2(n324), .ZN(
        n5180) );
  MOAI22 U14110 ( .A1(n28157), .A2(n323), .B1(ram[940]), .B2(n324), .ZN(
        n5181) );
  MOAI22 U14111 ( .A1(n27922), .A2(n323), .B1(ram[941]), .B2(n324), .ZN(
        n5182) );
  MOAI22 U14112 ( .A1(n27687), .A2(n323), .B1(ram[942]), .B2(n324), .ZN(
        n5183) );
  MOAI22 U14113 ( .A1(n27452), .A2(n323), .B1(ram[943]), .B2(n324), .ZN(
        n5184) );
  MOAI22 U14114 ( .A1(n29097), .A2(n325), .B1(ram[944]), .B2(n326), .ZN(
        n5185) );
  MOAI22 U14115 ( .A1(n28862), .A2(n325), .B1(ram[945]), .B2(n326), .ZN(
        n5186) );
  MOAI22 U14116 ( .A1(n28627), .A2(n325), .B1(ram[946]), .B2(n326), .ZN(
        n5187) );
  MOAI22 U14117 ( .A1(n28392), .A2(n325), .B1(ram[947]), .B2(n326), .ZN(
        n5188) );
  MOAI22 U14118 ( .A1(n28157), .A2(n325), .B1(ram[948]), .B2(n326), .ZN(
        n5189) );
  MOAI22 U14119 ( .A1(n27922), .A2(n325), .B1(ram[949]), .B2(n326), .ZN(
        n5190) );
  MOAI22 U14120 ( .A1(n27687), .A2(n325), .B1(ram[950]), .B2(n326), .ZN(
        n5191) );
  MOAI22 U14121 ( .A1(n27452), .A2(n325), .B1(ram[951]), .B2(n326), .ZN(
        n5192) );
  MOAI22 U14122 ( .A1(n29097), .A2(n327), .B1(ram[952]), .B2(n328), .ZN(
        n5193) );
  MOAI22 U14123 ( .A1(n28862), .A2(n327), .B1(ram[953]), .B2(n328), .ZN(
        n5194) );
  MOAI22 U14124 ( .A1(n28627), .A2(n327), .B1(ram[954]), .B2(n328), .ZN(
        n5195) );
  MOAI22 U14125 ( .A1(n28392), .A2(n327), .B1(ram[955]), .B2(n328), .ZN(
        n5196) );
  MOAI22 U14126 ( .A1(n28157), .A2(n327), .B1(ram[956]), .B2(n328), .ZN(
        n5197) );
  MOAI22 U14127 ( .A1(n27922), .A2(n327), .B1(ram[957]), .B2(n328), .ZN(
        n5198) );
  MOAI22 U14128 ( .A1(n27687), .A2(n327), .B1(ram[958]), .B2(n328), .ZN(
        n5199) );
  MOAI22 U14129 ( .A1(n27452), .A2(n327), .B1(ram[959]), .B2(n328), .ZN(
        n5200) );
  MOAI22 U14130 ( .A1(n29097), .A2(n329), .B1(ram[960]), .B2(n330), .ZN(
        n5201) );
  MOAI22 U14131 ( .A1(n28862), .A2(n329), .B1(ram[961]), .B2(n330), .ZN(
        n5202) );
  MOAI22 U14132 ( .A1(n28627), .A2(n329), .B1(ram[962]), .B2(n330), .ZN(
        n5203) );
  MOAI22 U14133 ( .A1(n28392), .A2(n329), .B1(ram[963]), .B2(n330), .ZN(
        n5204) );
  MOAI22 U14134 ( .A1(n28157), .A2(n329), .B1(ram[964]), .B2(n330), .ZN(
        n5205) );
  MOAI22 U14135 ( .A1(n27922), .A2(n329), .B1(ram[965]), .B2(n330), .ZN(
        n5206) );
  MOAI22 U14136 ( .A1(n27687), .A2(n329), .B1(ram[966]), .B2(n330), .ZN(
        n5207) );
  MOAI22 U14137 ( .A1(n27452), .A2(n329), .B1(ram[967]), .B2(n330), .ZN(
        n5208) );
  MOAI22 U14138 ( .A1(n29097), .A2(n331), .B1(ram[968]), .B2(n332), .ZN(
        n5209) );
  MOAI22 U14139 ( .A1(n28862), .A2(n331), .B1(ram[969]), .B2(n332), .ZN(
        n5210) );
  MOAI22 U14140 ( .A1(n28627), .A2(n331), .B1(ram[970]), .B2(n332), .ZN(
        n5211) );
  MOAI22 U14141 ( .A1(n28392), .A2(n331), .B1(ram[971]), .B2(n332), .ZN(
        n5212) );
  MOAI22 U14142 ( .A1(n28157), .A2(n331), .B1(ram[972]), .B2(n332), .ZN(
        n5213) );
  MOAI22 U14143 ( .A1(n27922), .A2(n331), .B1(ram[973]), .B2(n332), .ZN(
        n5214) );
  MOAI22 U14144 ( .A1(n27687), .A2(n331), .B1(ram[974]), .B2(n332), .ZN(
        n5215) );
  MOAI22 U14145 ( .A1(n27452), .A2(n331), .B1(ram[975]), .B2(n332), .ZN(
        n5216) );
  MOAI22 U14146 ( .A1(n29097), .A2(n333), .B1(ram[976]), .B2(n334), .ZN(
        n5217) );
  MOAI22 U14147 ( .A1(n28862), .A2(n333), .B1(ram[977]), .B2(n334), .ZN(
        n5218) );
  MOAI22 U14148 ( .A1(n28627), .A2(n333), .B1(ram[978]), .B2(n334), .ZN(
        n5219) );
  MOAI22 U14149 ( .A1(n28392), .A2(n333), .B1(ram[979]), .B2(n334), .ZN(
        n5220) );
  MOAI22 U14150 ( .A1(n28157), .A2(n333), .B1(ram[980]), .B2(n334), .ZN(
        n5221) );
  MOAI22 U14151 ( .A1(n27922), .A2(n333), .B1(ram[981]), .B2(n334), .ZN(
        n5222) );
  MOAI22 U14152 ( .A1(n27687), .A2(n333), .B1(ram[982]), .B2(n334), .ZN(
        n5223) );
  MOAI22 U14153 ( .A1(n27452), .A2(n333), .B1(ram[983]), .B2(n334), .ZN(
        n5224) );
  MOAI22 U14154 ( .A1(n29097), .A2(n335), .B1(ram[984]), .B2(n336), .ZN(
        n5225) );
  MOAI22 U14155 ( .A1(n28862), .A2(n335), .B1(ram[985]), .B2(n336), .ZN(
        n5226) );
  MOAI22 U14156 ( .A1(n28627), .A2(n335), .B1(ram[986]), .B2(n336), .ZN(
        n5227) );
  MOAI22 U14157 ( .A1(n28392), .A2(n335), .B1(ram[987]), .B2(n336), .ZN(
        n5228) );
  MOAI22 U14158 ( .A1(n28157), .A2(n335), .B1(ram[988]), .B2(n336), .ZN(
        n5229) );
  MOAI22 U14159 ( .A1(n27922), .A2(n335), .B1(ram[989]), .B2(n336), .ZN(
        n5230) );
  MOAI22 U14160 ( .A1(n27687), .A2(n335), .B1(ram[990]), .B2(n336), .ZN(
        n5231) );
  MOAI22 U14161 ( .A1(n27452), .A2(n335), .B1(ram[991]), .B2(n336), .ZN(
        n5232) );
  MOAI22 U14162 ( .A1(n29097), .A2(n337), .B1(ram[992]), .B2(n338), .ZN(
        n5233) );
  MOAI22 U14163 ( .A1(n28862), .A2(n337), .B1(ram[993]), .B2(n338), .ZN(
        n5234) );
  MOAI22 U14164 ( .A1(n28627), .A2(n337), .B1(ram[994]), .B2(n338), .ZN(
        n5235) );
  MOAI22 U14165 ( .A1(n28392), .A2(n337), .B1(ram[995]), .B2(n338), .ZN(
        n5236) );
  MOAI22 U14166 ( .A1(n28157), .A2(n337), .B1(ram[996]), .B2(n338), .ZN(
        n5237) );
  MOAI22 U14167 ( .A1(n27922), .A2(n337), .B1(ram[997]), .B2(n338), .ZN(
        n5238) );
  MOAI22 U14168 ( .A1(n27687), .A2(n337), .B1(ram[998]), .B2(n338), .ZN(
        n5239) );
  MOAI22 U14169 ( .A1(n27452), .A2(n337), .B1(ram[999]), .B2(n338), .ZN(
        n5240) );
  MOAI22 U14170 ( .A1(n29097), .A2(n339), .B1(ram[1000]), .B2(n340), .ZN(
        n5241) );
  MOAI22 U14171 ( .A1(n28862), .A2(n339), .B1(ram[1001]), .B2(n340), .ZN(
        n5242) );
  MOAI22 U14172 ( .A1(n28627), .A2(n339), .B1(ram[1002]), .B2(n340), .ZN(
        n5243) );
  MOAI22 U14173 ( .A1(n28392), .A2(n339), .B1(ram[1003]), .B2(n340), .ZN(
        n5244) );
  MOAI22 U14174 ( .A1(n28157), .A2(n339), .B1(ram[1004]), .B2(n340), .ZN(
        n5245) );
  MOAI22 U14175 ( .A1(n27922), .A2(n339), .B1(ram[1005]), .B2(n340), .ZN(
        n5246) );
  MOAI22 U14176 ( .A1(n27687), .A2(n339), .B1(ram[1006]), .B2(n340), .ZN(
        n5247) );
  MOAI22 U14177 ( .A1(n27452), .A2(n339), .B1(ram[1007]), .B2(n340), .ZN(
        n5248) );
  MOAI22 U14178 ( .A1(n29097), .A2(n341), .B1(ram[1008]), .B2(n342), .ZN(
        n5249) );
  MOAI22 U14179 ( .A1(n28862), .A2(n341), .B1(ram[1009]), .B2(n342), .ZN(
        n5250) );
  MOAI22 U14180 ( .A1(n28627), .A2(n341), .B1(ram[1010]), .B2(n342), .ZN(
        n5251) );
  MOAI22 U14181 ( .A1(n28392), .A2(n341), .B1(ram[1011]), .B2(n342), .ZN(
        n5252) );
  MOAI22 U14182 ( .A1(n28157), .A2(n341), .B1(ram[1012]), .B2(n342), .ZN(
        n5253) );
  MOAI22 U14183 ( .A1(n27922), .A2(n341), .B1(ram[1013]), .B2(n342), .ZN(
        n5254) );
  MOAI22 U14184 ( .A1(n27687), .A2(n341), .B1(ram[1014]), .B2(n342), .ZN(
        n5255) );
  MOAI22 U14185 ( .A1(n27452), .A2(n341), .B1(ram[1015]), .B2(n342), .ZN(
        n5256) );
  MOAI22 U14186 ( .A1(n29097), .A2(n343), .B1(ram[1016]), .B2(n344), .ZN(
        n5257) );
  MOAI22 U14187 ( .A1(n28862), .A2(n343), .B1(ram[1017]), .B2(n344), .ZN(
        n5258) );
  MOAI22 U14188 ( .A1(n28627), .A2(n343), .B1(ram[1018]), .B2(n344), .ZN(
        n5259) );
  MOAI22 U14189 ( .A1(n28392), .A2(n343), .B1(ram[1019]), .B2(n344), .ZN(
        n5260) );
  MOAI22 U14190 ( .A1(n28157), .A2(n343), .B1(ram[1020]), .B2(n344), .ZN(
        n5261) );
  MOAI22 U14191 ( .A1(n27922), .A2(n343), .B1(ram[1021]), .B2(n344), .ZN(
        n5262) );
  MOAI22 U14192 ( .A1(n27687), .A2(n343), .B1(ram[1022]), .B2(n344), .ZN(
        n5263) );
  MOAI22 U14193 ( .A1(n27452), .A2(n343), .B1(ram[1023]), .B2(n344), .ZN(
        n5264) );
  MOAI22 U14194 ( .A1(n29097), .A2(n346), .B1(ram[1024]), .B2(n347), .ZN(
        n5265) );
  MOAI22 U14195 ( .A1(n28862), .A2(n346), .B1(ram[1025]), .B2(n347), .ZN(
        n5266) );
  MOAI22 U14196 ( .A1(n28627), .A2(n346), .B1(ram[1026]), .B2(n347), .ZN(
        n5267) );
  MOAI22 U14197 ( .A1(n28392), .A2(n346), .B1(ram[1027]), .B2(n347), .ZN(
        n5268) );
  MOAI22 U14198 ( .A1(n28157), .A2(n346), .B1(ram[1028]), .B2(n347), .ZN(
        n5269) );
  MOAI22 U14199 ( .A1(n27922), .A2(n346), .B1(ram[1029]), .B2(n347), .ZN(
        n5270) );
  MOAI22 U14200 ( .A1(n27687), .A2(n346), .B1(ram[1030]), .B2(n347), .ZN(
        n5271) );
  MOAI22 U14201 ( .A1(n27452), .A2(n346), .B1(ram[1031]), .B2(n347), .ZN(
        n5272) );
  MOAI22 U14202 ( .A1(n29097), .A2(n349), .B1(ram[1032]), .B2(n350), .ZN(
        n5273) );
  MOAI22 U14203 ( .A1(n28862), .A2(n349), .B1(ram[1033]), .B2(n350), .ZN(
        n5274) );
  MOAI22 U14204 ( .A1(n28627), .A2(n349), .B1(ram[1034]), .B2(n350), .ZN(
        n5275) );
  MOAI22 U14205 ( .A1(n28392), .A2(n349), .B1(ram[1035]), .B2(n350), .ZN(
        n5276) );
  MOAI22 U14206 ( .A1(n28157), .A2(n349), .B1(ram[1036]), .B2(n350), .ZN(
        n5277) );
  MOAI22 U14207 ( .A1(n27922), .A2(n349), .B1(ram[1037]), .B2(n350), .ZN(
        n5278) );
  MOAI22 U14208 ( .A1(n27687), .A2(n349), .B1(ram[1038]), .B2(n350), .ZN(
        n5279) );
  MOAI22 U14209 ( .A1(n27452), .A2(n349), .B1(ram[1039]), .B2(n350), .ZN(
        n5280) );
  MOAI22 U14210 ( .A1(n29098), .A2(n351), .B1(ram[1040]), .B2(n352), .ZN(
        n5281) );
  MOAI22 U14211 ( .A1(n28863), .A2(n351), .B1(ram[1041]), .B2(n352), .ZN(
        n5282) );
  MOAI22 U14212 ( .A1(n28628), .A2(n351), .B1(ram[1042]), .B2(n352), .ZN(
        n5283) );
  MOAI22 U14213 ( .A1(n28393), .A2(n351), .B1(ram[1043]), .B2(n352), .ZN(
        n5284) );
  MOAI22 U14214 ( .A1(n28158), .A2(n351), .B1(ram[1044]), .B2(n352), .ZN(
        n5285) );
  MOAI22 U14215 ( .A1(n27923), .A2(n351), .B1(ram[1045]), .B2(n352), .ZN(
        n5286) );
  MOAI22 U14216 ( .A1(n27688), .A2(n351), .B1(ram[1046]), .B2(n352), .ZN(
        n5287) );
  MOAI22 U14217 ( .A1(n27453), .A2(n351), .B1(ram[1047]), .B2(n352), .ZN(
        n5288) );
  MOAI22 U14218 ( .A1(n29098), .A2(n353), .B1(ram[1048]), .B2(n354), .ZN(
        n5289) );
  MOAI22 U14219 ( .A1(n28863), .A2(n353), .B1(ram[1049]), .B2(n354), .ZN(
        n5290) );
  MOAI22 U14220 ( .A1(n28628), .A2(n353), .B1(ram[1050]), .B2(n354), .ZN(
        n5291) );
  MOAI22 U14221 ( .A1(n28393), .A2(n353), .B1(ram[1051]), .B2(n354), .ZN(
        n5292) );
  MOAI22 U14222 ( .A1(n28158), .A2(n353), .B1(ram[1052]), .B2(n354), .ZN(
        n5293) );
  MOAI22 U14223 ( .A1(n27923), .A2(n353), .B1(ram[1053]), .B2(n354), .ZN(
        n5294) );
  MOAI22 U14224 ( .A1(n27688), .A2(n353), .B1(ram[1054]), .B2(n354), .ZN(
        n5295) );
  MOAI22 U14225 ( .A1(n27453), .A2(n353), .B1(ram[1055]), .B2(n354), .ZN(
        n5296) );
  MOAI22 U14226 ( .A1(n29098), .A2(n355), .B1(ram[1056]), .B2(n356), .ZN(
        n5297) );
  MOAI22 U14227 ( .A1(n28863), .A2(n355), .B1(ram[1057]), .B2(n356), .ZN(
        n5298) );
  MOAI22 U14228 ( .A1(n28628), .A2(n355), .B1(ram[1058]), .B2(n356), .ZN(
        n5299) );
  MOAI22 U14229 ( .A1(n28393), .A2(n355), .B1(ram[1059]), .B2(n356), .ZN(
        n5300) );
  MOAI22 U14230 ( .A1(n28158), .A2(n355), .B1(ram[1060]), .B2(n356), .ZN(
        n5301) );
  MOAI22 U14231 ( .A1(n27923), .A2(n355), .B1(ram[1061]), .B2(n356), .ZN(
        n5302) );
  MOAI22 U14232 ( .A1(n27688), .A2(n355), .B1(ram[1062]), .B2(n356), .ZN(
        n5303) );
  MOAI22 U14233 ( .A1(n27453), .A2(n355), .B1(ram[1063]), .B2(n356), .ZN(
        n5304) );
  MOAI22 U14234 ( .A1(n29098), .A2(n357), .B1(ram[1064]), .B2(n358), .ZN(
        n5305) );
  MOAI22 U14235 ( .A1(n28863), .A2(n357), .B1(ram[1065]), .B2(n358), .ZN(
        n5306) );
  MOAI22 U14236 ( .A1(n28628), .A2(n357), .B1(ram[1066]), .B2(n358), .ZN(
        n5307) );
  MOAI22 U14237 ( .A1(n28393), .A2(n357), .B1(ram[1067]), .B2(n358), .ZN(
        n5308) );
  MOAI22 U14238 ( .A1(n28158), .A2(n357), .B1(ram[1068]), .B2(n358), .ZN(
        n5309) );
  MOAI22 U14239 ( .A1(n27923), .A2(n357), .B1(ram[1069]), .B2(n358), .ZN(
        n5310) );
  MOAI22 U14240 ( .A1(n27688), .A2(n357), .B1(ram[1070]), .B2(n358), .ZN(
        n5311) );
  MOAI22 U14241 ( .A1(n27453), .A2(n357), .B1(ram[1071]), .B2(n358), .ZN(
        n5312) );
  MOAI22 U14242 ( .A1(n29098), .A2(n359), .B1(ram[1072]), .B2(n360), .ZN(
        n5313) );
  MOAI22 U14243 ( .A1(n28863), .A2(n359), .B1(ram[1073]), .B2(n360), .ZN(
        n5314) );
  MOAI22 U14244 ( .A1(n28628), .A2(n359), .B1(ram[1074]), .B2(n360), .ZN(
        n5315) );
  MOAI22 U14245 ( .A1(n28393), .A2(n359), .B1(ram[1075]), .B2(n360), .ZN(
        n5316) );
  MOAI22 U14246 ( .A1(n28158), .A2(n359), .B1(ram[1076]), .B2(n360), .ZN(
        n5317) );
  MOAI22 U14247 ( .A1(n27923), .A2(n359), .B1(ram[1077]), .B2(n360), .ZN(
        n5318) );
  MOAI22 U14248 ( .A1(n27688), .A2(n359), .B1(ram[1078]), .B2(n360), .ZN(
        n5319) );
  MOAI22 U14249 ( .A1(n27453), .A2(n359), .B1(ram[1079]), .B2(n360), .ZN(
        n5320) );
  MOAI22 U14250 ( .A1(n29098), .A2(n361), .B1(ram[1080]), .B2(n362), .ZN(
        n5321) );
  MOAI22 U14251 ( .A1(n28863), .A2(n361), .B1(ram[1081]), .B2(n362), .ZN(
        n5322) );
  MOAI22 U14252 ( .A1(n28628), .A2(n361), .B1(ram[1082]), .B2(n362), .ZN(
        n5323) );
  MOAI22 U14253 ( .A1(n28393), .A2(n361), .B1(ram[1083]), .B2(n362), .ZN(
        n5324) );
  MOAI22 U14254 ( .A1(n28158), .A2(n361), .B1(ram[1084]), .B2(n362), .ZN(
        n5325) );
  MOAI22 U14255 ( .A1(n27923), .A2(n361), .B1(ram[1085]), .B2(n362), .ZN(
        n5326) );
  MOAI22 U14256 ( .A1(n27688), .A2(n361), .B1(ram[1086]), .B2(n362), .ZN(
        n5327) );
  MOAI22 U14257 ( .A1(n27453), .A2(n361), .B1(ram[1087]), .B2(n362), .ZN(
        n5328) );
  MOAI22 U14258 ( .A1(n29098), .A2(n363), .B1(ram[1088]), .B2(n364), .ZN(
        n5329) );
  MOAI22 U14259 ( .A1(n28863), .A2(n363), .B1(ram[1089]), .B2(n364), .ZN(
        n5330) );
  MOAI22 U14260 ( .A1(n28628), .A2(n363), .B1(ram[1090]), .B2(n364), .ZN(
        n5331) );
  MOAI22 U14261 ( .A1(n28393), .A2(n363), .B1(ram[1091]), .B2(n364), .ZN(
        n5332) );
  MOAI22 U14262 ( .A1(n28158), .A2(n363), .B1(ram[1092]), .B2(n364), .ZN(
        n5333) );
  MOAI22 U14263 ( .A1(n27923), .A2(n363), .B1(ram[1093]), .B2(n364), .ZN(
        n5334) );
  MOAI22 U14264 ( .A1(n27688), .A2(n363), .B1(ram[1094]), .B2(n364), .ZN(
        n5335) );
  MOAI22 U14265 ( .A1(n27453), .A2(n363), .B1(ram[1095]), .B2(n364), .ZN(
        n5336) );
  MOAI22 U14266 ( .A1(n29098), .A2(n365), .B1(ram[1096]), .B2(n366), .ZN(
        n5337) );
  MOAI22 U14267 ( .A1(n28863), .A2(n365), .B1(ram[1097]), .B2(n366), .ZN(
        n5338) );
  MOAI22 U14268 ( .A1(n28628), .A2(n365), .B1(ram[1098]), .B2(n366), .ZN(
        n5339) );
  MOAI22 U14269 ( .A1(n28393), .A2(n365), .B1(ram[1099]), .B2(n366), .ZN(
        n5340) );
  MOAI22 U14270 ( .A1(n28158), .A2(n365), .B1(ram[1100]), .B2(n366), .ZN(
        n5341) );
  MOAI22 U14271 ( .A1(n27923), .A2(n365), .B1(ram[1101]), .B2(n366), .ZN(
        n5342) );
  MOAI22 U14272 ( .A1(n27688), .A2(n365), .B1(ram[1102]), .B2(n366), .ZN(
        n5343) );
  MOAI22 U14273 ( .A1(n27453), .A2(n365), .B1(ram[1103]), .B2(n366), .ZN(
        n5344) );
  MOAI22 U14274 ( .A1(n29098), .A2(n367), .B1(ram[1104]), .B2(n368), .ZN(
        n5345) );
  MOAI22 U14275 ( .A1(n28863), .A2(n367), .B1(ram[1105]), .B2(n368), .ZN(
        n5346) );
  MOAI22 U14276 ( .A1(n28628), .A2(n367), .B1(ram[1106]), .B2(n368), .ZN(
        n5347) );
  MOAI22 U14277 ( .A1(n28393), .A2(n367), .B1(ram[1107]), .B2(n368), .ZN(
        n5348) );
  MOAI22 U14278 ( .A1(n28158), .A2(n367), .B1(ram[1108]), .B2(n368), .ZN(
        n5349) );
  MOAI22 U14279 ( .A1(n27923), .A2(n367), .B1(ram[1109]), .B2(n368), .ZN(
        n5350) );
  MOAI22 U14280 ( .A1(n27688), .A2(n367), .B1(ram[1110]), .B2(n368), .ZN(
        n5351) );
  MOAI22 U14281 ( .A1(n27453), .A2(n367), .B1(ram[1111]), .B2(n368), .ZN(
        n5352) );
  MOAI22 U14282 ( .A1(n29098), .A2(n369), .B1(ram[1112]), .B2(n370), .ZN(
        n5353) );
  MOAI22 U14283 ( .A1(n28863), .A2(n369), .B1(ram[1113]), .B2(n370), .ZN(
        n5354) );
  MOAI22 U14284 ( .A1(n28628), .A2(n369), .B1(ram[1114]), .B2(n370), .ZN(
        n5355) );
  MOAI22 U14285 ( .A1(n28393), .A2(n369), .B1(ram[1115]), .B2(n370), .ZN(
        n5356) );
  MOAI22 U14286 ( .A1(n28158), .A2(n369), .B1(ram[1116]), .B2(n370), .ZN(
        n5357) );
  MOAI22 U14287 ( .A1(n27923), .A2(n369), .B1(ram[1117]), .B2(n370), .ZN(
        n5358) );
  MOAI22 U14288 ( .A1(n27688), .A2(n369), .B1(ram[1118]), .B2(n370), .ZN(
        n5359) );
  MOAI22 U14289 ( .A1(n27453), .A2(n369), .B1(ram[1119]), .B2(n370), .ZN(
        n5360) );
  MOAI22 U14290 ( .A1(n29098), .A2(n371), .B1(ram[1120]), .B2(n372), .ZN(
        n5361) );
  MOAI22 U14291 ( .A1(n28863), .A2(n371), .B1(ram[1121]), .B2(n372), .ZN(
        n5362) );
  MOAI22 U14292 ( .A1(n28628), .A2(n371), .B1(ram[1122]), .B2(n372), .ZN(
        n5363) );
  MOAI22 U14293 ( .A1(n28393), .A2(n371), .B1(ram[1123]), .B2(n372), .ZN(
        n5364) );
  MOAI22 U14294 ( .A1(n28158), .A2(n371), .B1(ram[1124]), .B2(n372), .ZN(
        n5365) );
  MOAI22 U14295 ( .A1(n27923), .A2(n371), .B1(ram[1125]), .B2(n372), .ZN(
        n5366) );
  MOAI22 U14296 ( .A1(n27688), .A2(n371), .B1(ram[1126]), .B2(n372), .ZN(
        n5367) );
  MOAI22 U14297 ( .A1(n27453), .A2(n371), .B1(ram[1127]), .B2(n372), .ZN(
        n5368) );
  MOAI22 U14298 ( .A1(n29098), .A2(n373), .B1(ram[1128]), .B2(n374), .ZN(
        n5369) );
  MOAI22 U14299 ( .A1(n28863), .A2(n373), .B1(ram[1129]), .B2(n374), .ZN(
        n5370) );
  MOAI22 U14300 ( .A1(n28628), .A2(n373), .B1(ram[1130]), .B2(n374), .ZN(
        n5371) );
  MOAI22 U14301 ( .A1(n28393), .A2(n373), .B1(ram[1131]), .B2(n374), .ZN(
        n5372) );
  MOAI22 U14302 ( .A1(n28158), .A2(n373), .B1(ram[1132]), .B2(n374), .ZN(
        n5373) );
  MOAI22 U14303 ( .A1(n27923), .A2(n373), .B1(ram[1133]), .B2(n374), .ZN(
        n5374) );
  MOAI22 U14304 ( .A1(n27688), .A2(n373), .B1(ram[1134]), .B2(n374), .ZN(
        n5375) );
  MOAI22 U14305 ( .A1(n27453), .A2(n373), .B1(ram[1135]), .B2(n374), .ZN(
        n5376) );
  MOAI22 U14306 ( .A1(n29098), .A2(n375), .B1(ram[1136]), .B2(n376), .ZN(
        n5377) );
  MOAI22 U14307 ( .A1(n28863), .A2(n375), .B1(ram[1137]), .B2(n376), .ZN(
        n5378) );
  MOAI22 U14308 ( .A1(n28628), .A2(n375), .B1(ram[1138]), .B2(n376), .ZN(
        n5379) );
  MOAI22 U14309 ( .A1(n28393), .A2(n375), .B1(ram[1139]), .B2(n376), .ZN(
        n5380) );
  MOAI22 U14310 ( .A1(n28158), .A2(n375), .B1(ram[1140]), .B2(n376), .ZN(
        n5381) );
  MOAI22 U14311 ( .A1(n27923), .A2(n375), .B1(ram[1141]), .B2(n376), .ZN(
        n5382) );
  MOAI22 U14312 ( .A1(n27688), .A2(n375), .B1(ram[1142]), .B2(n376), .ZN(
        n5383) );
  MOAI22 U14313 ( .A1(n27453), .A2(n375), .B1(ram[1143]), .B2(n376), .ZN(
        n5384) );
  MOAI22 U14314 ( .A1(n29099), .A2(n377), .B1(ram[1144]), .B2(n378), .ZN(
        n5385) );
  MOAI22 U14315 ( .A1(n28864), .A2(n377), .B1(ram[1145]), .B2(n378), .ZN(
        n5386) );
  MOAI22 U14316 ( .A1(n28629), .A2(n377), .B1(ram[1146]), .B2(n378), .ZN(
        n5387) );
  MOAI22 U14317 ( .A1(n28394), .A2(n377), .B1(ram[1147]), .B2(n378), .ZN(
        n5388) );
  MOAI22 U14318 ( .A1(n28159), .A2(n377), .B1(ram[1148]), .B2(n378), .ZN(
        n5389) );
  MOAI22 U14319 ( .A1(n27924), .A2(n377), .B1(ram[1149]), .B2(n378), .ZN(
        n5390) );
  MOAI22 U14320 ( .A1(n27689), .A2(n377), .B1(ram[1150]), .B2(n378), .ZN(
        n5391) );
  MOAI22 U14321 ( .A1(n27454), .A2(n377), .B1(ram[1151]), .B2(n378), .ZN(
        n5392) );
  MOAI22 U14322 ( .A1(n29099), .A2(n379), .B1(ram[1152]), .B2(n380), .ZN(
        n5393) );
  MOAI22 U14323 ( .A1(n28864), .A2(n379), .B1(ram[1153]), .B2(n380), .ZN(
        n5394) );
  MOAI22 U14324 ( .A1(n28629), .A2(n379), .B1(ram[1154]), .B2(n380), .ZN(
        n5395) );
  MOAI22 U14325 ( .A1(n28394), .A2(n379), .B1(ram[1155]), .B2(n380), .ZN(
        n5396) );
  MOAI22 U14326 ( .A1(n28159), .A2(n379), .B1(ram[1156]), .B2(n380), .ZN(
        n5397) );
  MOAI22 U14327 ( .A1(n27924), .A2(n379), .B1(ram[1157]), .B2(n380), .ZN(
        n5398) );
  MOAI22 U14328 ( .A1(n27689), .A2(n379), .B1(ram[1158]), .B2(n380), .ZN(
        n5399) );
  MOAI22 U14329 ( .A1(n27454), .A2(n379), .B1(ram[1159]), .B2(n380), .ZN(
        n5400) );
  MOAI22 U14330 ( .A1(n29099), .A2(n381), .B1(ram[1160]), .B2(n382), .ZN(
        n5401) );
  MOAI22 U14331 ( .A1(n28864), .A2(n381), .B1(ram[1161]), .B2(n382), .ZN(
        n5402) );
  MOAI22 U14332 ( .A1(n28629), .A2(n381), .B1(ram[1162]), .B2(n382), .ZN(
        n5403) );
  MOAI22 U14333 ( .A1(n28394), .A2(n381), .B1(ram[1163]), .B2(n382), .ZN(
        n5404) );
  MOAI22 U14334 ( .A1(n28159), .A2(n381), .B1(ram[1164]), .B2(n382), .ZN(
        n5405) );
  MOAI22 U14335 ( .A1(n27924), .A2(n381), .B1(ram[1165]), .B2(n382), .ZN(
        n5406) );
  MOAI22 U14336 ( .A1(n27689), .A2(n381), .B1(ram[1166]), .B2(n382), .ZN(
        n5407) );
  MOAI22 U14337 ( .A1(n27454), .A2(n381), .B1(ram[1167]), .B2(n382), .ZN(
        n5408) );
  MOAI22 U14338 ( .A1(n29099), .A2(n383), .B1(ram[1168]), .B2(n384), .ZN(
        n5409) );
  MOAI22 U14339 ( .A1(n28864), .A2(n383), .B1(ram[1169]), .B2(n384), .ZN(
        n5410) );
  MOAI22 U14340 ( .A1(n28629), .A2(n383), .B1(ram[1170]), .B2(n384), .ZN(
        n5411) );
  MOAI22 U14341 ( .A1(n28394), .A2(n383), .B1(ram[1171]), .B2(n384), .ZN(
        n5412) );
  MOAI22 U14342 ( .A1(n28159), .A2(n383), .B1(ram[1172]), .B2(n384), .ZN(
        n5413) );
  MOAI22 U14343 ( .A1(n27924), .A2(n383), .B1(ram[1173]), .B2(n384), .ZN(
        n5414) );
  MOAI22 U14344 ( .A1(n27689), .A2(n383), .B1(ram[1174]), .B2(n384), .ZN(
        n5415) );
  MOAI22 U14345 ( .A1(n27454), .A2(n383), .B1(ram[1175]), .B2(n384), .ZN(
        n5416) );
  MOAI22 U14346 ( .A1(n29099), .A2(n385), .B1(ram[1176]), .B2(n386), .ZN(
        n5417) );
  MOAI22 U14347 ( .A1(n28864), .A2(n385), .B1(ram[1177]), .B2(n386), .ZN(
        n5418) );
  MOAI22 U14348 ( .A1(n28629), .A2(n385), .B1(ram[1178]), .B2(n386), .ZN(
        n5419) );
  MOAI22 U14349 ( .A1(n28394), .A2(n385), .B1(ram[1179]), .B2(n386), .ZN(
        n5420) );
  MOAI22 U14350 ( .A1(n28159), .A2(n385), .B1(ram[1180]), .B2(n386), .ZN(
        n5421) );
  MOAI22 U14351 ( .A1(n27924), .A2(n385), .B1(ram[1181]), .B2(n386), .ZN(
        n5422) );
  MOAI22 U14352 ( .A1(n27689), .A2(n385), .B1(ram[1182]), .B2(n386), .ZN(
        n5423) );
  MOAI22 U14353 ( .A1(n27454), .A2(n385), .B1(ram[1183]), .B2(n386), .ZN(
        n5424) );
  MOAI22 U14354 ( .A1(n29099), .A2(n387), .B1(ram[1184]), .B2(n388), .ZN(
        n5425) );
  MOAI22 U14355 ( .A1(n28864), .A2(n387), .B1(ram[1185]), .B2(n388), .ZN(
        n5426) );
  MOAI22 U14356 ( .A1(n28629), .A2(n387), .B1(ram[1186]), .B2(n388), .ZN(
        n5427) );
  MOAI22 U14357 ( .A1(n28394), .A2(n387), .B1(ram[1187]), .B2(n388), .ZN(
        n5428) );
  MOAI22 U14358 ( .A1(n28159), .A2(n387), .B1(ram[1188]), .B2(n388), .ZN(
        n5429) );
  MOAI22 U14359 ( .A1(n27924), .A2(n387), .B1(ram[1189]), .B2(n388), .ZN(
        n5430) );
  MOAI22 U14360 ( .A1(n27689), .A2(n387), .B1(ram[1190]), .B2(n388), .ZN(
        n5431) );
  MOAI22 U14361 ( .A1(n27454), .A2(n387), .B1(ram[1191]), .B2(n388), .ZN(
        n5432) );
  MOAI22 U14362 ( .A1(n29099), .A2(n389), .B1(ram[1192]), .B2(n390), .ZN(
        n5433) );
  MOAI22 U14363 ( .A1(n28864), .A2(n389), .B1(ram[1193]), .B2(n390), .ZN(
        n5434) );
  MOAI22 U14364 ( .A1(n28629), .A2(n389), .B1(ram[1194]), .B2(n390), .ZN(
        n5435) );
  MOAI22 U14365 ( .A1(n28394), .A2(n389), .B1(ram[1195]), .B2(n390), .ZN(
        n5436) );
  MOAI22 U14366 ( .A1(n28159), .A2(n389), .B1(ram[1196]), .B2(n390), .ZN(
        n5437) );
  MOAI22 U14367 ( .A1(n27924), .A2(n389), .B1(ram[1197]), .B2(n390), .ZN(
        n5438) );
  MOAI22 U14368 ( .A1(n27689), .A2(n389), .B1(ram[1198]), .B2(n390), .ZN(
        n5439) );
  MOAI22 U14369 ( .A1(n27454), .A2(n389), .B1(ram[1199]), .B2(n390), .ZN(
        n5440) );
  MOAI22 U14370 ( .A1(n29099), .A2(n391), .B1(ram[1200]), .B2(n392), .ZN(
        n5441) );
  MOAI22 U14371 ( .A1(n28864), .A2(n391), .B1(ram[1201]), .B2(n392), .ZN(
        n5442) );
  MOAI22 U14372 ( .A1(n28629), .A2(n391), .B1(ram[1202]), .B2(n392), .ZN(
        n5443) );
  MOAI22 U14373 ( .A1(n28394), .A2(n391), .B1(ram[1203]), .B2(n392), .ZN(
        n5444) );
  MOAI22 U14374 ( .A1(n28159), .A2(n391), .B1(ram[1204]), .B2(n392), .ZN(
        n5445) );
  MOAI22 U14375 ( .A1(n27924), .A2(n391), .B1(ram[1205]), .B2(n392), .ZN(
        n5446) );
  MOAI22 U14376 ( .A1(n27689), .A2(n391), .B1(ram[1206]), .B2(n392), .ZN(
        n5447) );
  MOAI22 U14377 ( .A1(n27454), .A2(n391), .B1(ram[1207]), .B2(n392), .ZN(
        n5448) );
  MOAI22 U14378 ( .A1(n29099), .A2(n393), .B1(ram[1208]), .B2(n394), .ZN(
        n5449) );
  MOAI22 U14379 ( .A1(n28864), .A2(n393), .B1(ram[1209]), .B2(n394), .ZN(
        n5450) );
  MOAI22 U14380 ( .A1(n28629), .A2(n393), .B1(ram[1210]), .B2(n394), .ZN(
        n5451) );
  MOAI22 U14381 ( .A1(n28394), .A2(n393), .B1(ram[1211]), .B2(n394), .ZN(
        n5452) );
  MOAI22 U14382 ( .A1(n28159), .A2(n393), .B1(ram[1212]), .B2(n394), .ZN(
        n5453) );
  MOAI22 U14383 ( .A1(n27924), .A2(n393), .B1(ram[1213]), .B2(n394), .ZN(
        n5454) );
  MOAI22 U14384 ( .A1(n27689), .A2(n393), .B1(ram[1214]), .B2(n394), .ZN(
        n5455) );
  MOAI22 U14385 ( .A1(n27454), .A2(n393), .B1(ram[1215]), .B2(n394), .ZN(
        n5456) );
  MOAI22 U14386 ( .A1(n29099), .A2(n395), .B1(ram[1216]), .B2(n396), .ZN(
        n5457) );
  MOAI22 U14387 ( .A1(n28864), .A2(n395), .B1(ram[1217]), .B2(n396), .ZN(
        n5458) );
  MOAI22 U14388 ( .A1(n28629), .A2(n395), .B1(ram[1218]), .B2(n396), .ZN(
        n5459) );
  MOAI22 U14389 ( .A1(n28394), .A2(n395), .B1(ram[1219]), .B2(n396), .ZN(
        n5460) );
  MOAI22 U14390 ( .A1(n28159), .A2(n395), .B1(ram[1220]), .B2(n396), .ZN(
        n5461) );
  MOAI22 U14391 ( .A1(n27924), .A2(n395), .B1(ram[1221]), .B2(n396), .ZN(
        n5462) );
  MOAI22 U14392 ( .A1(n27689), .A2(n395), .B1(ram[1222]), .B2(n396), .ZN(
        n5463) );
  MOAI22 U14393 ( .A1(n27454), .A2(n395), .B1(ram[1223]), .B2(n396), .ZN(
        n5464) );
  MOAI22 U14394 ( .A1(n29099), .A2(n397), .B1(ram[1224]), .B2(n398), .ZN(
        n5465) );
  MOAI22 U14395 ( .A1(n28864), .A2(n397), .B1(ram[1225]), .B2(n398), .ZN(
        n5466) );
  MOAI22 U14396 ( .A1(n28629), .A2(n397), .B1(ram[1226]), .B2(n398), .ZN(
        n5467) );
  MOAI22 U14397 ( .A1(n28394), .A2(n397), .B1(ram[1227]), .B2(n398), .ZN(
        n5468) );
  MOAI22 U14398 ( .A1(n28159), .A2(n397), .B1(ram[1228]), .B2(n398), .ZN(
        n5469) );
  MOAI22 U14399 ( .A1(n27924), .A2(n397), .B1(ram[1229]), .B2(n398), .ZN(
        n5470) );
  MOAI22 U14400 ( .A1(n27689), .A2(n397), .B1(ram[1230]), .B2(n398), .ZN(
        n5471) );
  MOAI22 U14401 ( .A1(n27454), .A2(n397), .B1(ram[1231]), .B2(n398), .ZN(
        n5472) );
  MOAI22 U14402 ( .A1(n29099), .A2(n399), .B1(ram[1232]), .B2(n400), .ZN(
        n5473) );
  MOAI22 U14403 ( .A1(n28864), .A2(n399), .B1(ram[1233]), .B2(n400), .ZN(
        n5474) );
  MOAI22 U14404 ( .A1(n28629), .A2(n399), .B1(ram[1234]), .B2(n400), .ZN(
        n5475) );
  MOAI22 U14405 ( .A1(n28394), .A2(n399), .B1(ram[1235]), .B2(n400), .ZN(
        n5476) );
  MOAI22 U14406 ( .A1(n28159), .A2(n399), .B1(ram[1236]), .B2(n400), .ZN(
        n5477) );
  MOAI22 U14407 ( .A1(n27924), .A2(n399), .B1(ram[1237]), .B2(n400), .ZN(
        n5478) );
  MOAI22 U14408 ( .A1(n27689), .A2(n399), .B1(ram[1238]), .B2(n400), .ZN(
        n5479) );
  MOAI22 U14409 ( .A1(n27454), .A2(n399), .B1(ram[1239]), .B2(n400), .ZN(
        n5480) );
  MOAI22 U14410 ( .A1(n29099), .A2(n401), .B1(ram[1240]), .B2(n402), .ZN(
        n5481) );
  MOAI22 U14411 ( .A1(n28864), .A2(n401), .B1(ram[1241]), .B2(n402), .ZN(
        n5482) );
  MOAI22 U14412 ( .A1(n28629), .A2(n401), .B1(ram[1242]), .B2(n402), .ZN(
        n5483) );
  MOAI22 U14413 ( .A1(n28394), .A2(n401), .B1(ram[1243]), .B2(n402), .ZN(
        n5484) );
  MOAI22 U14414 ( .A1(n28159), .A2(n401), .B1(ram[1244]), .B2(n402), .ZN(
        n5485) );
  MOAI22 U14415 ( .A1(n27924), .A2(n401), .B1(ram[1245]), .B2(n402), .ZN(
        n5486) );
  MOAI22 U14416 ( .A1(n27689), .A2(n401), .B1(ram[1246]), .B2(n402), .ZN(
        n5487) );
  MOAI22 U14417 ( .A1(n27454), .A2(n401), .B1(ram[1247]), .B2(n402), .ZN(
        n5488) );
  MOAI22 U14418 ( .A1(n29100), .A2(n403), .B1(ram[1248]), .B2(n404), .ZN(
        n5489) );
  MOAI22 U14419 ( .A1(n28865), .A2(n403), .B1(ram[1249]), .B2(n404), .ZN(
        n5490) );
  MOAI22 U14420 ( .A1(n28630), .A2(n403), .B1(ram[1250]), .B2(n404), .ZN(
        n5491) );
  MOAI22 U14421 ( .A1(n28395), .A2(n403), .B1(ram[1251]), .B2(n404), .ZN(
        n5492) );
  MOAI22 U14422 ( .A1(n28160), .A2(n403), .B1(ram[1252]), .B2(n404), .ZN(
        n5493) );
  MOAI22 U14423 ( .A1(n27925), .A2(n403), .B1(ram[1253]), .B2(n404), .ZN(
        n5494) );
  MOAI22 U14424 ( .A1(n27690), .A2(n403), .B1(ram[1254]), .B2(n404), .ZN(
        n5495) );
  MOAI22 U14425 ( .A1(n27455), .A2(n403), .B1(ram[1255]), .B2(n404), .ZN(
        n5496) );
  MOAI22 U14426 ( .A1(n29100), .A2(n405), .B1(ram[1256]), .B2(n406), .ZN(
        n5497) );
  MOAI22 U14427 ( .A1(n28865), .A2(n405), .B1(ram[1257]), .B2(n406), .ZN(
        n5498) );
  MOAI22 U14428 ( .A1(n28630), .A2(n405), .B1(ram[1258]), .B2(n406), .ZN(
        n5499) );
  MOAI22 U14429 ( .A1(n28395), .A2(n405), .B1(ram[1259]), .B2(n406), .ZN(
        n5500) );
  MOAI22 U14430 ( .A1(n28160), .A2(n405), .B1(ram[1260]), .B2(n406), .ZN(
        n5501) );
  MOAI22 U14431 ( .A1(n27925), .A2(n405), .B1(ram[1261]), .B2(n406), .ZN(
        n5502) );
  MOAI22 U14432 ( .A1(n27690), .A2(n405), .B1(ram[1262]), .B2(n406), .ZN(
        n5503) );
  MOAI22 U14433 ( .A1(n27455), .A2(n405), .B1(ram[1263]), .B2(n406), .ZN(
        n5504) );
  MOAI22 U14434 ( .A1(n29100), .A2(n407), .B1(ram[1264]), .B2(n408), .ZN(
        n5505) );
  MOAI22 U14435 ( .A1(n28865), .A2(n407), .B1(ram[1265]), .B2(n408), .ZN(
        n5506) );
  MOAI22 U14436 ( .A1(n28630), .A2(n407), .B1(ram[1266]), .B2(n408), .ZN(
        n5507) );
  MOAI22 U14437 ( .A1(n28395), .A2(n407), .B1(ram[1267]), .B2(n408), .ZN(
        n5508) );
  MOAI22 U14438 ( .A1(n28160), .A2(n407), .B1(ram[1268]), .B2(n408), .ZN(
        n5509) );
  MOAI22 U14439 ( .A1(n27925), .A2(n407), .B1(ram[1269]), .B2(n408), .ZN(
        n5510) );
  MOAI22 U14440 ( .A1(n27690), .A2(n407), .B1(ram[1270]), .B2(n408), .ZN(
        n5511) );
  MOAI22 U14441 ( .A1(n27455), .A2(n407), .B1(ram[1271]), .B2(n408), .ZN(
        n5512) );
  MOAI22 U14442 ( .A1(n29100), .A2(n409), .B1(ram[1272]), .B2(n410), .ZN(
        n5513) );
  MOAI22 U14443 ( .A1(n28865), .A2(n409), .B1(ram[1273]), .B2(n410), .ZN(
        n5514) );
  MOAI22 U14444 ( .A1(n28630), .A2(n409), .B1(ram[1274]), .B2(n410), .ZN(
        n5515) );
  MOAI22 U14445 ( .A1(n28395), .A2(n409), .B1(ram[1275]), .B2(n410), .ZN(
        n5516) );
  MOAI22 U14446 ( .A1(n28160), .A2(n409), .B1(ram[1276]), .B2(n410), .ZN(
        n5517) );
  MOAI22 U14447 ( .A1(n27925), .A2(n409), .B1(ram[1277]), .B2(n410), .ZN(
        n5518) );
  MOAI22 U14448 ( .A1(n27690), .A2(n409), .B1(ram[1278]), .B2(n410), .ZN(
        n5519) );
  MOAI22 U14449 ( .A1(n27455), .A2(n409), .B1(ram[1279]), .B2(n410), .ZN(
        n5520) );
  MOAI22 U14450 ( .A1(n29100), .A2(n411), .B1(ram[1280]), .B2(n412), .ZN(
        n5521) );
  MOAI22 U14451 ( .A1(n28865), .A2(n411), .B1(ram[1281]), .B2(n412), .ZN(
        n5522) );
  MOAI22 U14452 ( .A1(n28630), .A2(n411), .B1(ram[1282]), .B2(n412), .ZN(
        n5523) );
  MOAI22 U14453 ( .A1(n28395), .A2(n411), .B1(ram[1283]), .B2(n412), .ZN(
        n5524) );
  MOAI22 U14454 ( .A1(n28160), .A2(n411), .B1(ram[1284]), .B2(n412), .ZN(
        n5525) );
  MOAI22 U14455 ( .A1(n27925), .A2(n411), .B1(ram[1285]), .B2(n412), .ZN(
        n5526) );
  MOAI22 U14456 ( .A1(n27690), .A2(n411), .B1(ram[1286]), .B2(n412), .ZN(
        n5527) );
  MOAI22 U14457 ( .A1(n27455), .A2(n411), .B1(ram[1287]), .B2(n412), .ZN(
        n5528) );
  MOAI22 U14458 ( .A1(n29100), .A2(n413), .B1(ram[1288]), .B2(n414), .ZN(
        n5529) );
  MOAI22 U14459 ( .A1(n28865), .A2(n413), .B1(ram[1289]), .B2(n414), .ZN(
        n5530) );
  MOAI22 U14460 ( .A1(n28630), .A2(n413), .B1(ram[1290]), .B2(n414), .ZN(
        n5531) );
  MOAI22 U14461 ( .A1(n28395), .A2(n413), .B1(ram[1291]), .B2(n414), .ZN(
        n5532) );
  MOAI22 U14462 ( .A1(n28160), .A2(n413), .B1(ram[1292]), .B2(n414), .ZN(
        n5533) );
  MOAI22 U14463 ( .A1(n27925), .A2(n413), .B1(ram[1293]), .B2(n414), .ZN(
        n5534) );
  MOAI22 U14464 ( .A1(n27690), .A2(n413), .B1(ram[1294]), .B2(n414), .ZN(
        n5535) );
  MOAI22 U14465 ( .A1(n27455), .A2(n413), .B1(ram[1295]), .B2(n414), .ZN(
        n5536) );
  MOAI22 U14466 ( .A1(n29100), .A2(n415), .B1(ram[1296]), .B2(n416), .ZN(
        n5537) );
  MOAI22 U14467 ( .A1(n28865), .A2(n415), .B1(ram[1297]), .B2(n416), .ZN(
        n5538) );
  MOAI22 U14468 ( .A1(n28630), .A2(n415), .B1(ram[1298]), .B2(n416), .ZN(
        n5539) );
  MOAI22 U14469 ( .A1(n28395), .A2(n415), .B1(ram[1299]), .B2(n416), .ZN(
        n5540) );
  MOAI22 U14470 ( .A1(n28160), .A2(n415), .B1(ram[1300]), .B2(n416), .ZN(
        n5541) );
  MOAI22 U14471 ( .A1(n27925), .A2(n415), .B1(ram[1301]), .B2(n416), .ZN(
        n5542) );
  MOAI22 U14472 ( .A1(n27690), .A2(n415), .B1(ram[1302]), .B2(n416), .ZN(
        n5543) );
  MOAI22 U14473 ( .A1(n27455), .A2(n415), .B1(ram[1303]), .B2(n416), .ZN(
        n5544) );
  MOAI22 U14474 ( .A1(n29100), .A2(n417), .B1(ram[1304]), .B2(n418), .ZN(
        n5545) );
  MOAI22 U14475 ( .A1(n28865), .A2(n417), .B1(ram[1305]), .B2(n418), .ZN(
        n5546) );
  MOAI22 U14476 ( .A1(n28630), .A2(n417), .B1(ram[1306]), .B2(n418), .ZN(
        n5547) );
  MOAI22 U14477 ( .A1(n28395), .A2(n417), .B1(ram[1307]), .B2(n418), .ZN(
        n5548) );
  MOAI22 U14478 ( .A1(n28160), .A2(n417), .B1(ram[1308]), .B2(n418), .ZN(
        n5549) );
  MOAI22 U14479 ( .A1(n27925), .A2(n417), .B1(ram[1309]), .B2(n418), .ZN(
        n5550) );
  MOAI22 U14480 ( .A1(n27690), .A2(n417), .B1(ram[1310]), .B2(n418), .ZN(
        n5551) );
  MOAI22 U14481 ( .A1(n27455), .A2(n417), .B1(ram[1311]), .B2(n418), .ZN(
        n5552) );
  MOAI22 U14482 ( .A1(n29100), .A2(n419), .B1(ram[1312]), .B2(n420), .ZN(
        n5553) );
  MOAI22 U14483 ( .A1(n28865), .A2(n419), .B1(ram[1313]), .B2(n420), .ZN(
        n5554) );
  MOAI22 U14484 ( .A1(n28630), .A2(n419), .B1(ram[1314]), .B2(n420), .ZN(
        n5555) );
  MOAI22 U14485 ( .A1(n28395), .A2(n419), .B1(ram[1315]), .B2(n420), .ZN(
        n5556) );
  MOAI22 U14486 ( .A1(n28160), .A2(n419), .B1(ram[1316]), .B2(n420), .ZN(
        n5557) );
  MOAI22 U14487 ( .A1(n27925), .A2(n419), .B1(ram[1317]), .B2(n420), .ZN(
        n5558) );
  MOAI22 U14488 ( .A1(n27690), .A2(n419), .B1(ram[1318]), .B2(n420), .ZN(
        n5559) );
  MOAI22 U14489 ( .A1(n27455), .A2(n419), .B1(ram[1319]), .B2(n420), .ZN(
        n5560) );
  MOAI22 U14490 ( .A1(n29100), .A2(n421), .B1(ram[1320]), .B2(n422), .ZN(
        n5561) );
  MOAI22 U14491 ( .A1(n28865), .A2(n421), .B1(ram[1321]), .B2(n422), .ZN(
        n5562) );
  MOAI22 U14492 ( .A1(n28630), .A2(n421), .B1(ram[1322]), .B2(n422), .ZN(
        n5563) );
  MOAI22 U14493 ( .A1(n28395), .A2(n421), .B1(ram[1323]), .B2(n422), .ZN(
        n5564) );
  MOAI22 U14494 ( .A1(n28160), .A2(n421), .B1(ram[1324]), .B2(n422), .ZN(
        n5565) );
  MOAI22 U14495 ( .A1(n27925), .A2(n421), .B1(ram[1325]), .B2(n422), .ZN(
        n5566) );
  MOAI22 U14496 ( .A1(n27690), .A2(n421), .B1(ram[1326]), .B2(n422), .ZN(
        n5567) );
  MOAI22 U14497 ( .A1(n27455), .A2(n421), .B1(ram[1327]), .B2(n422), .ZN(
        n5568) );
  MOAI22 U14498 ( .A1(n29100), .A2(n423), .B1(ram[1328]), .B2(n424), .ZN(
        n5569) );
  MOAI22 U14499 ( .A1(n28865), .A2(n423), .B1(ram[1329]), .B2(n424), .ZN(
        n5570) );
  MOAI22 U14500 ( .A1(n28630), .A2(n423), .B1(ram[1330]), .B2(n424), .ZN(
        n5571) );
  MOAI22 U14501 ( .A1(n28395), .A2(n423), .B1(ram[1331]), .B2(n424), .ZN(
        n5572) );
  MOAI22 U14502 ( .A1(n28160), .A2(n423), .B1(ram[1332]), .B2(n424), .ZN(
        n5573) );
  MOAI22 U14503 ( .A1(n27925), .A2(n423), .B1(ram[1333]), .B2(n424), .ZN(
        n5574) );
  MOAI22 U14504 ( .A1(n27690), .A2(n423), .B1(ram[1334]), .B2(n424), .ZN(
        n5575) );
  MOAI22 U14505 ( .A1(n27455), .A2(n423), .B1(ram[1335]), .B2(n424), .ZN(
        n5576) );
  MOAI22 U14506 ( .A1(n29100), .A2(n425), .B1(ram[1336]), .B2(n426), .ZN(
        n5577) );
  MOAI22 U14507 ( .A1(n28865), .A2(n425), .B1(ram[1337]), .B2(n426), .ZN(
        n5578) );
  MOAI22 U14508 ( .A1(n28630), .A2(n425), .B1(ram[1338]), .B2(n426), .ZN(
        n5579) );
  MOAI22 U14509 ( .A1(n28395), .A2(n425), .B1(ram[1339]), .B2(n426), .ZN(
        n5580) );
  MOAI22 U14510 ( .A1(n28160), .A2(n425), .B1(ram[1340]), .B2(n426), .ZN(
        n5581) );
  MOAI22 U14511 ( .A1(n27925), .A2(n425), .B1(ram[1341]), .B2(n426), .ZN(
        n5582) );
  MOAI22 U14512 ( .A1(n27690), .A2(n425), .B1(ram[1342]), .B2(n426), .ZN(
        n5583) );
  MOAI22 U14513 ( .A1(n27455), .A2(n425), .B1(ram[1343]), .B2(n426), .ZN(
        n5584) );
  MOAI22 U14514 ( .A1(n29100), .A2(n427), .B1(ram[1344]), .B2(n428), .ZN(
        n5585) );
  MOAI22 U14515 ( .A1(n28865), .A2(n427), .B1(ram[1345]), .B2(n428), .ZN(
        n5586) );
  MOAI22 U14516 ( .A1(n28630), .A2(n427), .B1(ram[1346]), .B2(n428), .ZN(
        n5587) );
  MOAI22 U14517 ( .A1(n28395), .A2(n427), .B1(ram[1347]), .B2(n428), .ZN(
        n5588) );
  MOAI22 U14518 ( .A1(n28160), .A2(n427), .B1(ram[1348]), .B2(n428), .ZN(
        n5589) );
  MOAI22 U14519 ( .A1(n27925), .A2(n427), .B1(ram[1349]), .B2(n428), .ZN(
        n5590) );
  MOAI22 U14520 ( .A1(n27690), .A2(n427), .B1(ram[1350]), .B2(n428), .ZN(
        n5591) );
  MOAI22 U14521 ( .A1(n27455), .A2(n427), .B1(ram[1351]), .B2(n428), .ZN(
        n5592) );
  MOAI22 U14522 ( .A1(n29101), .A2(n429), .B1(ram[1352]), .B2(n430), .ZN(
        n5593) );
  MOAI22 U14523 ( .A1(n28866), .A2(n429), .B1(ram[1353]), .B2(n430), .ZN(
        n5594) );
  MOAI22 U14524 ( .A1(n28631), .A2(n429), .B1(ram[1354]), .B2(n430), .ZN(
        n5595) );
  MOAI22 U14525 ( .A1(n28396), .A2(n429), .B1(ram[1355]), .B2(n430), .ZN(
        n5596) );
  MOAI22 U14526 ( .A1(n28161), .A2(n429), .B1(ram[1356]), .B2(n430), .ZN(
        n5597) );
  MOAI22 U14527 ( .A1(n27926), .A2(n429), .B1(ram[1357]), .B2(n430), .ZN(
        n5598) );
  MOAI22 U14528 ( .A1(n27691), .A2(n429), .B1(ram[1358]), .B2(n430), .ZN(
        n5599) );
  MOAI22 U14529 ( .A1(n27456), .A2(n429), .B1(ram[1359]), .B2(n430), .ZN(
        n5600) );
  MOAI22 U14530 ( .A1(n29101), .A2(n431), .B1(ram[1360]), .B2(n432), .ZN(
        n5601) );
  MOAI22 U14531 ( .A1(n28866), .A2(n431), .B1(ram[1361]), .B2(n432), .ZN(
        n5602) );
  MOAI22 U14532 ( .A1(n28631), .A2(n431), .B1(ram[1362]), .B2(n432), .ZN(
        n5603) );
  MOAI22 U14533 ( .A1(n28396), .A2(n431), .B1(ram[1363]), .B2(n432), .ZN(
        n5604) );
  MOAI22 U14534 ( .A1(n28161), .A2(n431), .B1(ram[1364]), .B2(n432), .ZN(
        n5605) );
  MOAI22 U14535 ( .A1(n27926), .A2(n431), .B1(ram[1365]), .B2(n432), .ZN(
        n5606) );
  MOAI22 U14536 ( .A1(n27691), .A2(n431), .B1(ram[1366]), .B2(n432), .ZN(
        n5607) );
  MOAI22 U14537 ( .A1(n27456), .A2(n431), .B1(ram[1367]), .B2(n432), .ZN(
        n5608) );
  MOAI22 U14538 ( .A1(n29101), .A2(n433), .B1(ram[1368]), .B2(n434), .ZN(
        n5609) );
  MOAI22 U14539 ( .A1(n28866), .A2(n433), .B1(ram[1369]), .B2(n434), .ZN(
        n5610) );
  MOAI22 U14540 ( .A1(n28631), .A2(n433), .B1(ram[1370]), .B2(n434), .ZN(
        n5611) );
  MOAI22 U14541 ( .A1(n28396), .A2(n433), .B1(ram[1371]), .B2(n434), .ZN(
        n5612) );
  MOAI22 U14542 ( .A1(n28161), .A2(n433), .B1(ram[1372]), .B2(n434), .ZN(
        n5613) );
  MOAI22 U14543 ( .A1(n27926), .A2(n433), .B1(ram[1373]), .B2(n434), .ZN(
        n5614) );
  MOAI22 U14544 ( .A1(n27691), .A2(n433), .B1(ram[1374]), .B2(n434), .ZN(
        n5615) );
  MOAI22 U14545 ( .A1(n27456), .A2(n433), .B1(ram[1375]), .B2(n434), .ZN(
        n5616) );
  MOAI22 U14546 ( .A1(n29101), .A2(n435), .B1(ram[1376]), .B2(n436), .ZN(
        n5617) );
  MOAI22 U14547 ( .A1(n28866), .A2(n435), .B1(ram[1377]), .B2(n436), .ZN(
        n5618) );
  MOAI22 U14548 ( .A1(n28631), .A2(n435), .B1(ram[1378]), .B2(n436), .ZN(
        n5619) );
  MOAI22 U14549 ( .A1(n28396), .A2(n435), .B1(ram[1379]), .B2(n436), .ZN(
        n5620) );
  MOAI22 U14550 ( .A1(n28161), .A2(n435), .B1(ram[1380]), .B2(n436), .ZN(
        n5621) );
  MOAI22 U14551 ( .A1(n27926), .A2(n435), .B1(ram[1381]), .B2(n436), .ZN(
        n5622) );
  MOAI22 U14552 ( .A1(n27691), .A2(n435), .B1(ram[1382]), .B2(n436), .ZN(
        n5623) );
  MOAI22 U14553 ( .A1(n27456), .A2(n435), .B1(ram[1383]), .B2(n436), .ZN(
        n5624) );
  MOAI22 U14554 ( .A1(n29101), .A2(n437), .B1(ram[1384]), .B2(n438), .ZN(
        n5625) );
  MOAI22 U14555 ( .A1(n28866), .A2(n437), .B1(ram[1385]), .B2(n438), .ZN(
        n5626) );
  MOAI22 U14556 ( .A1(n28631), .A2(n437), .B1(ram[1386]), .B2(n438), .ZN(
        n5627) );
  MOAI22 U14557 ( .A1(n28396), .A2(n437), .B1(ram[1387]), .B2(n438), .ZN(
        n5628) );
  MOAI22 U14558 ( .A1(n28161), .A2(n437), .B1(ram[1388]), .B2(n438), .ZN(
        n5629) );
  MOAI22 U14559 ( .A1(n27926), .A2(n437), .B1(ram[1389]), .B2(n438), .ZN(
        n5630) );
  MOAI22 U14560 ( .A1(n27691), .A2(n437), .B1(ram[1390]), .B2(n438), .ZN(
        n5631) );
  MOAI22 U14561 ( .A1(n27456), .A2(n437), .B1(ram[1391]), .B2(n438), .ZN(
        n5632) );
  MOAI22 U14562 ( .A1(n29101), .A2(n439), .B1(ram[1392]), .B2(n440), .ZN(
        n5633) );
  MOAI22 U14563 ( .A1(n28866), .A2(n439), .B1(ram[1393]), .B2(n440), .ZN(
        n5634) );
  MOAI22 U14564 ( .A1(n28631), .A2(n439), .B1(ram[1394]), .B2(n440), .ZN(
        n5635) );
  MOAI22 U14565 ( .A1(n28396), .A2(n439), .B1(ram[1395]), .B2(n440), .ZN(
        n5636) );
  MOAI22 U14566 ( .A1(n28161), .A2(n439), .B1(ram[1396]), .B2(n440), .ZN(
        n5637) );
  MOAI22 U14567 ( .A1(n27926), .A2(n439), .B1(ram[1397]), .B2(n440), .ZN(
        n5638) );
  MOAI22 U14568 ( .A1(n27691), .A2(n439), .B1(ram[1398]), .B2(n440), .ZN(
        n5639) );
  MOAI22 U14569 ( .A1(n27456), .A2(n439), .B1(ram[1399]), .B2(n440), .ZN(
        n5640) );
  MOAI22 U14570 ( .A1(n29101), .A2(n441), .B1(ram[1400]), .B2(n442), .ZN(
        n5641) );
  MOAI22 U14571 ( .A1(n28866), .A2(n441), .B1(ram[1401]), .B2(n442), .ZN(
        n5642) );
  MOAI22 U14572 ( .A1(n28631), .A2(n441), .B1(ram[1402]), .B2(n442), .ZN(
        n5643) );
  MOAI22 U14573 ( .A1(n28396), .A2(n441), .B1(ram[1403]), .B2(n442), .ZN(
        n5644) );
  MOAI22 U14574 ( .A1(n28161), .A2(n441), .B1(ram[1404]), .B2(n442), .ZN(
        n5645) );
  MOAI22 U14575 ( .A1(n27926), .A2(n441), .B1(ram[1405]), .B2(n442), .ZN(
        n5646) );
  MOAI22 U14576 ( .A1(n27691), .A2(n441), .B1(ram[1406]), .B2(n442), .ZN(
        n5647) );
  MOAI22 U14577 ( .A1(n27456), .A2(n441), .B1(ram[1407]), .B2(n442), .ZN(
        n5648) );
  MOAI22 U14578 ( .A1(n29101), .A2(n443), .B1(ram[1408]), .B2(n444), .ZN(
        n5649) );
  MOAI22 U14579 ( .A1(n28866), .A2(n443), .B1(ram[1409]), .B2(n444), .ZN(
        n5650) );
  MOAI22 U14580 ( .A1(n28631), .A2(n443), .B1(ram[1410]), .B2(n444), .ZN(
        n5651) );
  MOAI22 U14581 ( .A1(n28396), .A2(n443), .B1(ram[1411]), .B2(n444), .ZN(
        n5652) );
  MOAI22 U14582 ( .A1(n28161), .A2(n443), .B1(ram[1412]), .B2(n444), .ZN(
        n5653) );
  MOAI22 U14583 ( .A1(n27926), .A2(n443), .B1(ram[1413]), .B2(n444), .ZN(
        n5654) );
  MOAI22 U14584 ( .A1(n27691), .A2(n443), .B1(ram[1414]), .B2(n444), .ZN(
        n5655) );
  MOAI22 U14585 ( .A1(n27456), .A2(n443), .B1(ram[1415]), .B2(n444), .ZN(
        n5656) );
  MOAI22 U14586 ( .A1(n29101), .A2(n445), .B1(ram[1416]), .B2(n446), .ZN(
        n5657) );
  MOAI22 U14587 ( .A1(n28866), .A2(n445), .B1(ram[1417]), .B2(n446), .ZN(
        n5658) );
  MOAI22 U14588 ( .A1(n28631), .A2(n445), .B1(ram[1418]), .B2(n446), .ZN(
        n5659) );
  MOAI22 U14589 ( .A1(n28396), .A2(n445), .B1(ram[1419]), .B2(n446), .ZN(
        n5660) );
  MOAI22 U14590 ( .A1(n28161), .A2(n445), .B1(ram[1420]), .B2(n446), .ZN(
        n5661) );
  MOAI22 U14591 ( .A1(n27926), .A2(n445), .B1(ram[1421]), .B2(n446), .ZN(
        n5662) );
  MOAI22 U14592 ( .A1(n27691), .A2(n445), .B1(ram[1422]), .B2(n446), .ZN(
        n5663) );
  MOAI22 U14593 ( .A1(n27456), .A2(n445), .B1(ram[1423]), .B2(n446), .ZN(
        n5664) );
  MOAI22 U14594 ( .A1(n29101), .A2(n447), .B1(ram[1424]), .B2(n448), .ZN(
        n5665) );
  MOAI22 U14595 ( .A1(n28866), .A2(n447), .B1(ram[1425]), .B2(n448), .ZN(
        n5666) );
  MOAI22 U14596 ( .A1(n28631), .A2(n447), .B1(ram[1426]), .B2(n448), .ZN(
        n5667) );
  MOAI22 U14597 ( .A1(n28396), .A2(n447), .B1(ram[1427]), .B2(n448), .ZN(
        n5668) );
  MOAI22 U14598 ( .A1(n28161), .A2(n447), .B1(ram[1428]), .B2(n448), .ZN(
        n5669) );
  MOAI22 U14599 ( .A1(n27926), .A2(n447), .B1(ram[1429]), .B2(n448), .ZN(
        n5670) );
  MOAI22 U14600 ( .A1(n27691), .A2(n447), .B1(ram[1430]), .B2(n448), .ZN(
        n5671) );
  MOAI22 U14601 ( .A1(n27456), .A2(n447), .B1(ram[1431]), .B2(n448), .ZN(
        n5672) );
  MOAI22 U14602 ( .A1(n29101), .A2(n449), .B1(ram[1432]), .B2(n450), .ZN(
        n5673) );
  MOAI22 U14603 ( .A1(n28866), .A2(n449), .B1(ram[1433]), .B2(n450), .ZN(
        n5674) );
  MOAI22 U14604 ( .A1(n28631), .A2(n449), .B1(ram[1434]), .B2(n450), .ZN(
        n5675) );
  MOAI22 U14605 ( .A1(n28396), .A2(n449), .B1(ram[1435]), .B2(n450), .ZN(
        n5676) );
  MOAI22 U14606 ( .A1(n28161), .A2(n449), .B1(ram[1436]), .B2(n450), .ZN(
        n5677) );
  MOAI22 U14607 ( .A1(n27926), .A2(n449), .B1(ram[1437]), .B2(n450), .ZN(
        n5678) );
  MOAI22 U14608 ( .A1(n27691), .A2(n449), .B1(ram[1438]), .B2(n450), .ZN(
        n5679) );
  MOAI22 U14609 ( .A1(n27456), .A2(n449), .B1(ram[1439]), .B2(n450), .ZN(
        n5680) );
  MOAI22 U14610 ( .A1(n29101), .A2(n451), .B1(ram[1440]), .B2(n452), .ZN(
        n5681) );
  MOAI22 U14611 ( .A1(n28866), .A2(n451), .B1(ram[1441]), .B2(n452), .ZN(
        n5682) );
  MOAI22 U14612 ( .A1(n28631), .A2(n451), .B1(ram[1442]), .B2(n452), .ZN(
        n5683) );
  MOAI22 U14613 ( .A1(n28396), .A2(n451), .B1(ram[1443]), .B2(n452), .ZN(
        n5684) );
  MOAI22 U14614 ( .A1(n28161), .A2(n451), .B1(ram[1444]), .B2(n452), .ZN(
        n5685) );
  MOAI22 U14615 ( .A1(n27926), .A2(n451), .B1(ram[1445]), .B2(n452), .ZN(
        n5686) );
  MOAI22 U14616 ( .A1(n27691), .A2(n451), .B1(ram[1446]), .B2(n452), .ZN(
        n5687) );
  MOAI22 U14617 ( .A1(n27456), .A2(n451), .B1(ram[1447]), .B2(n452), .ZN(
        n5688) );
  MOAI22 U14618 ( .A1(n29101), .A2(n453), .B1(ram[1448]), .B2(n454), .ZN(
        n5689) );
  MOAI22 U14619 ( .A1(n28866), .A2(n453), .B1(ram[1449]), .B2(n454), .ZN(
        n5690) );
  MOAI22 U14620 ( .A1(n28631), .A2(n453), .B1(ram[1450]), .B2(n454), .ZN(
        n5691) );
  MOAI22 U14621 ( .A1(n28396), .A2(n453), .B1(ram[1451]), .B2(n454), .ZN(
        n5692) );
  MOAI22 U14622 ( .A1(n28161), .A2(n453), .B1(ram[1452]), .B2(n454), .ZN(
        n5693) );
  MOAI22 U14623 ( .A1(n27926), .A2(n453), .B1(ram[1453]), .B2(n454), .ZN(
        n5694) );
  MOAI22 U14624 ( .A1(n27691), .A2(n453), .B1(ram[1454]), .B2(n454), .ZN(
        n5695) );
  MOAI22 U14625 ( .A1(n27456), .A2(n453), .B1(ram[1455]), .B2(n454), .ZN(
        n5696) );
  MOAI22 U14626 ( .A1(n29102), .A2(n455), .B1(ram[1456]), .B2(n456), .ZN(
        n5697) );
  MOAI22 U14627 ( .A1(n28867), .A2(n455), .B1(ram[1457]), .B2(n456), .ZN(
        n5698) );
  MOAI22 U14628 ( .A1(n28632), .A2(n455), .B1(ram[1458]), .B2(n456), .ZN(
        n5699) );
  MOAI22 U14629 ( .A1(n28397), .A2(n455), .B1(ram[1459]), .B2(n456), .ZN(
        n5700) );
  MOAI22 U14630 ( .A1(n28162), .A2(n455), .B1(ram[1460]), .B2(n456), .ZN(
        n5701) );
  MOAI22 U14631 ( .A1(n27927), .A2(n455), .B1(ram[1461]), .B2(n456), .ZN(
        n5702) );
  MOAI22 U14632 ( .A1(n27692), .A2(n455), .B1(ram[1462]), .B2(n456), .ZN(
        n5703) );
  MOAI22 U14633 ( .A1(n27457), .A2(n455), .B1(ram[1463]), .B2(n456), .ZN(
        n5704) );
  MOAI22 U14634 ( .A1(n29102), .A2(n457), .B1(ram[1464]), .B2(n458), .ZN(
        n5705) );
  MOAI22 U14635 ( .A1(n28867), .A2(n457), .B1(ram[1465]), .B2(n458), .ZN(
        n5706) );
  MOAI22 U14636 ( .A1(n28632), .A2(n457), .B1(ram[1466]), .B2(n458), .ZN(
        n5707) );
  MOAI22 U14637 ( .A1(n28397), .A2(n457), .B1(ram[1467]), .B2(n458), .ZN(
        n5708) );
  MOAI22 U14638 ( .A1(n28162), .A2(n457), .B1(ram[1468]), .B2(n458), .ZN(
        n5709) );
  MOAI22 U14639 ( .A1(n27927), .A2(n457), .B1(ram[1469]), .B2(n458), .ZN(
        n5710) );
  MOAI22 U14640 ( .A1(n27692), .A2(n457), .B1(ram[1470]), .B2(n458), .ZN(
        n5711) );
  MOAI22 U14641 ( .A1(n27457), .A2(n457), .B1(ram[1471]), .B2(n458), .ZN(
        n5712) );
  MOAI22 U14642 ( .A1(n29102), .A2(n459), .B1(ram[1472]), .B2(n460), .ZN(
        n5713) );
  MOAI22 U14643 ( .A1(n28867), .A2(n459), .B1(ram[1473]), .B2(n460), .ZN(
        n5714) );
  MOAI22 U14644 ( .A1(n28632), .A2(n459), .B1(ram[1474]), .B2(n460), .ZN(
        n5715) );
  MOAI22 U14645 ( .A1(n28397), .A2(n459), .B1(ram[1475]), .B2(n460), .ZN(
        n5716) );
  MOAI22 U14646 ( .A1(n28162), .A2(n459), .B1(ram[1476]), .B2(n460), .ZN(
        n5717) );
  MOAI22 U14647 ( .A1(n27927), .A2(n459), .B1(ram[1477]), .B2(n460), .ZN(
        n5718) );
  MOAI22 U14648 ( .A1(n27692), .A2(n459), .B1(ram[1478]), .B2(n460), .ZN(
        n5719) );
  MOAI22 U14649 ( .A1(n27457), .A2(n459), .B1(ram[1479]), .B2(n460), .ZN(
        n5720) );
  MOAI22 U14650 ( .A1(n29102), .A2(n461), .B1(ram[1480]), .B2(n462), .ZN(
        n5721) );
  MOAI22 U14651 ( .A1(n28867), .A2(n461), .B1(ram[1481]), .B2(n462), .ZN(
        n5722) );
  MOAI22 U14652 ( .A1(n28632), .A2(n461), .B1(ram[1482]), .B2(n462), .ZN(
        n5723) );
  MOAI22 U14653 ( .A1(n28397), .A2(n461), .B1(ram[1483]), .B2(n462), .ZN(
        n5724) );
  MOAI22 U14654 ( .A1(n28162), .A2(n461), .B1(ram[1484]), .B2(n462), .ZN(
        n5725) );
  MOAI22 U14655 ( .A1(n27927), .A2(n461), .B1(ram[1485]), .B2(n462), .ZN(
        n5726) );
  MOAI22 U14656 ( .A1(n27692), .A2(n461), .B1(ram[1486]), .B2(n462), .ZN(
        n5727) );
  MOAI22 U14657 ( .A1(n27457), .A2(n461), .B1(ram[1487]), .B2(n462), .ZN(
        n5728) );
  MOAI22 U14658 ( .A1(n29102), .A2(n463), .B1(ram[1488]), .B2(n464), .ZN(
        n5729) );
  MOAI22 U14659 ( .A1(n28867), .A2(n463), .B1(ram[1489]), .B2(n464), .ZN(
        n5730) );
  MOAI22 U14660 ( .A1(n28632), .A2(n463), .B1(ram[1490]), .B2(n464), .ZN(
        n5731) );
  MOAI22 U14661 ( .A1(n28397), .A2(n463), .B1(ram[1491]), .B2(n464), .ZN(
        n5732) );
  MOAI22 U14662 ( .A1(n28162), .A2(n463), .B1(ram[1492]), .B2(n464), .ZN(
        n5733) );
  MOAI22 U14663 ( .A1(n27927), .A2(n463), .B1(ram[1493]), .B2(n464), .ZN(
        n5734) );
  MOAI22 U14664 ( .A1(n27692), .A2(n463), .B1(ram[1494]), .B2(n464), .ZN(
        n5735) );
  MOAI22 U14665 ( .A1(n27457), .A2(n463), .B1(ram[1495]), .B2(n464), .ZN(
        n5736) );
  MOAI22 U14666 ( .A1(n29102), .A2(n465), .B1(ram[1496]), .B2(n466), .ZN(
        n5737) );
  MOAI22 U14667 ( .A1(n28867), .A2(n465), .B1(ram[1497]), .B2(n466), .ZN(
        n5738) );
  MOAI22 U14668 ( .A1(n28632), .A2(n465), .B1(ram[1498]), .B2(n466), .ZN(
        n5739) );
  MOAI22 U14669 ( .A1(n28397), .A2(n465), .B1(ram[1499]), .B2(n466), .ZN(
        n5740) );
  MOAI22 U14670 ( .A1(n28162), .A2(n465), .B1(ram[1500]), .B2(n466), .ZN(
        n5741) );
  MOAI22 U14671 ( .A1(n27927), .A2(n465), .B1(ram[1501]), .B2(n466), .ZN(
        n5742) );
  MOAI22 U14672 ( .A1(n27692), .A2(n465), .B1(ram[1502]), .B2(n466), .ZN(
        n5743) );
  MOAI22 U14673 ( .A1(n27457), .A2(n465), .B1(ram[1503]), .B2(n466), .ZN(
        n5744) );
  MOAI22 U14674 ( .A1(n29102), .A2(n467), .B1(ram[1504]), .B2(n468), .ZN(
        n5745) );
  MOAI22 U14675 ( .A1(n28867), .A2(n467), .B1(ram[1505]), .B2(n468), .ZN(
        n5746) );
  MOAI22 U14676 ( .A1(n28632), .A2(n467), .B1(ram[1506]), .B2(n468), .ZN(
        n5747) );
  MOAI22 U14677 ( .A1(n28397), .A2(n467), .B1(ram[1507]), .B2(n468), .ZN(
        n5748) );
  MOAI22 U14678 ( .A1(n28162), .A2(n467), .B1(ram[1508]), .B2(n468), .ZN(
        n5749) );
  MOAI22 U14679 ( .A1(n27927), .A2(n467), .B1(ram[1509]), .B2(n468), .ZN(
        n5750) );
  MOAI22 U14680 ( .A1(n27692), .A2(n467), .B1(ram[1510]), .B2(n468), .ZN(
        n5751) );
  MOAI22 U14681 ( .A1(n27457), .A2(n467), .B1(ram[1511]), .B2(n468), .ZN(
        n5752) );
  MOAI22 U14682 ( .A1(n29102), .A2(n469), .B1(ram[1512]), .B2(n470), .ZN(
        n5753) );
  MOAI22 U14683 ( .A1(n28867), .A2(n469), .B1(ram[1513]), .B2(n470), .ZN(
        n5754) );
  MOAI22 U14684 ( .A1(n28632), .A2(n469), .B1(ram[1514]), .B2(n470), .ZN(
        n5755) );
  MOAI22 U14685 ( .A1(n28397), .A2(n469), .B1(ram[1515]), .B2(n470), .ZN(
        n5756) );
  MOAI22 U14686 ( .A1(n28162), .A2(n469), .B1(ram[1516]), .B2(n470), .ZN(
        n5757) );
  MOAI22 U14687 ( .A1(n27927), .A2(n469), .B1(ram[1517]), .B2(n470), .ZN(
        n5758) );
  MOAI22 U14688 ( .A1(n27692), .A2(n469), .B1(ram[1518]), .B2(n470), .ZN(
        n5759) );
  MOAI22 U14689 ( .A1(n27457), .A2(n469), .B1(ram[1519]), .B2(n470), .ZN(
        n5760) );
  MOAI22 U14690 ( .A1(n29102), .A2(n471), .B1(ram[1520]), .B2(n472), .ZN(
        n5761) );
  MOAI22 U14691 ( .A1(n28867), .A2(n471), .B1(ram[1521]), .B2(n472), .ZN(
        n5762) );
  MOAI22 U14692 ( .A1(n28632), .A2(n471), .B1(ram[1522]), .B2(n472), .ZN(
        n5763) );
  MOAI22 U14693 ( .A1(n28397), .A2(n471), .B1(ram[1523]), .B2(n472), .ZN(
        n5764) );
  MOAI22 U14694 ( .A1(n28162), .A2(n471), .B1(ram[1524]), .B2(n472), .ZN(
        n5765) );
  MOAI22 U14695 ( .A1(n27927), .A2(n471), .B1(ram[1525]), .B2(n472), .ZN(
        n5766) );
  MOAI22 U14696 ( .A1(n27692), .A2(n471), .B1(ram[1526]), .B2(n472), .ZN(
        n5767) );
  MOAI22 U14697 ( .A1(n27457), .A2(n471), .B1(ram[1527]), .B2(n472), .ZN(
        n5768) );
  MOAI22 U14698 ( .A1(n29102), .A2(n473), .B1(ram[1528]), .B2(n474), .ZN(
        n5769) );
  MOAI22 U14699 ( .A1(n28867), .A2(n473), .B1(ram[1529]), .B2(n474), .ZN(
        n5770) );
  MOAI22 U14700 ( .A1(n28632), .A2(n473), .B1(ram[1530]), .B2(n474), .ZN(
        n5771) );
  MOAI22 U14701 ( .A1(n28397), .A2(n473), .B1(ram[1531]), .B2(n474), .ZN(
        n5772) );
  MOAI22 U14702 ( .A1(n28162), .A2(n473), .B1(ram[1532]), .B2(n474), .ZN(
        n5773) );
  MOAI22 U14703 ( .A1(n27927), .A2(n473), .B1(ram[1533]), .B2(n474), .ZN(
        n5774) );
  MOAI22 U14704 ( .A1(n27692), .A2(n473), .B1(ram[1534]), .B2(n474), .ZN(
        n5775) );
  MOAI22 U14705 ( .A1(n27457), .A2(n473), .B1(ram[1535]), .B2(n474), .ZN(
        n5776) );
  MOAI22 U14706 ( .A1(n29102), .A2(n476), .B1(ram[1536]), .B2(n477), .ZN(
        n5777) );
  MOAI22 U14707 ( .A1(n28867), .A2(n476), .B1(ram[1537]), .B2(n477), .ZN(
        n5778) );
  MOAI22 U14708 ( .A1(n28632), .A2(n476), .B1(ram[1538]), .B2(n477), .ZN(
        n5779) );
  MOAI22 U14709 ( .A1(n28397), .A2(n476), .B1(ram[1539]), .B2(n477), .ZN(
        n5780) );
  MOAI22 U14710 ( .A1(n28162), .A2(n476), .B1(ram[1540]), .B2(n477), .ZN(
        n5781) );
  MOAI22 U14711 ( .A1(n27927), .A2(n476), .B1(ram[1541]), .B2(n477), .ZN(
        n5782) );
  MOAI22 U14712 ( .A1(n27692), .A2(n476), .B1(ram[1542]), .B2(n477), .ZN(
        n5783) );
  MOAI22 U14713 ( .A1(n27457), .A2(n476), .B1(ram[1543]), .B2(n477), .ZN(
        n5784) );
  MOAI22 U14714 ( .A1(n29102), .A2(n479), .B1(ram[1544]), .B2(n480), .ZN(
        n5785) );
  MOAI22 U14715 ( .A1(n28867), .A2(n479), .B1(ram[1545]), .B2(n480), .ZN(
        n5786) );
  MOAI22 U14716 ( .A1(n28632), .A2(n479), .B1(ram[1546]), .B2(n480), .ZN(
        n5787) );
  MOAI22 U14717 ( .A1(n28397), .A2(n479), .B1(ram[1547]), .B2(n480), .ZN(
        n5788) );
  MOAI22 U14718 ( .A1(n28162), .A2(n479), .B1(ram[1548]), .B2(n480), .ZN(
        n5789) );
  MOAI22 U14719 ( .A1(n27927), .A2(n479), .B1(ram[1549]), .B2(n480), .ZN(
        n5790) );
  MOAI22 U14720 ( .A1(n27692), .A2(n479), .B1(ram[1550]), .B2(n480), .ZN(
        n5791) );
  MOAI22 U14721 ( .A1(n27457), .A2(n479), .B1(ram[1551]), .B2(n480), .ZN(
        n5792) );
  MOAI22 U14722 ( .A1(n29102), .A2(n481), .B1(ram[1552]), .B2(n482), .ZN(
        n5793) );
  MOAI22 U14723 ( .A1(n28867), .A2(n481), .B1(ram[1553]), .B2(n482), .ZN(
        n5794) );
  MOAI22 U14724 ( .A1(n28632), .A2(n481), .B1(ram[1554]), .B2(n482), .ZN(
        n5795) );
  MOAI22 U14725 ( .A1(n28397), .A2(n481), .B1(ram[1555]), .B2(n482), .ZN(
        n5796) );
  MOAI22 U14726 ( .A1(n28162), .A2(n481), .B1(ram[1556]), .B2(n482), .ZN(
        n5797) );
  MOAI22 U14727 ( .A1(n27927), .A2(n481), .B1(ram[1557]), .B2(n482), .ZN(
        n5798) );
  MOAI22 U14728 ( .A1(n27692), .A2(n481), .B1(ram[1558]), .B2(n482), .ZN(
        n5799) );
  MOAI22 U14729 ( .A1(n27457), .A2(n481), .B1(ram[1559]), .B2(n482), .ZN(
        n5800) );
  MOAI22 U14730 ( .A1(n29103), .A2(n483), .B1(ram[1560]), .B2(n484), .ZN(
        n5801) );
  MOAI22 U14731 ( .A1(n28868), .A2(n483), .B1(ram[1561]), .B2(n484), .ZN(
        n5802) );
  MOAI22 U14732 ( .A1(n28633), .A2(n483), .B1(ram[1562]), .B2(n484), .ZN(
        n5803) );
  MOAI22 U14733 ( .A1(n28398), .A2(n483), .B1(ram[1563]), .B2(n484), .ZN(
        n5804) );
  MOAI22 U14734 ( .A1(n28163), .A2(n483), .B1(ram[1564]), .B2(n484), .ZN(
        n5805) );
  MOAI22 U14735 ( .A1(n27928), .A2(n483), .B1(ram[1565]), .B2(n484), .ZN(
        n5806) );
  MOAI22 U14736 ( .A1(n27693), .A2(n483), .B1(ram[1566]), .B2(n484), .ZN(
        n5807) );
  MOAI22 U14737 ( .A1(n27458), .A2(n483), .B1(ram[1567]), .B2(n484), .ZN(
        n5808) );
  MOAI22 U14738 ( .A1(n29103), .A2(n485), .B1(ram[1568]), .B2(n486), .ZN(
        n5809) );
  MOAI22 U14739 ( .A1(n28868), .A2(n485), .B1(ram[1569]), .B2(n486), .ZN(
        n5810) );
  MOAI22 U14740 ( .A1(n28633), .A2(n485), .B1(ram[1570]), .B2(n486), .ZN(
        n5811) );
  MOAI22 U14741 ( .A1(n28398), .A2(n485), .B1(ram[1571]), .B2(n486), .ZN(
        n5812) );
  MOAI22 U14742 ( .A1(n28163), .A2(n485), .B1(ram[1572]), .B2(n486), .ZN(
        n5813) );
  MOAI22 U14743 ( .A1(n27928), .A2(n485), .B1(ram[1573]), .B2(n486), .ZN(
        n5814) );
  MOAI22 U14744 ( .A1(n27693), .A2(n485), .B1(ram[1574]), .B2(n486), .ZN(
        n5815) );
  MOAI22 U14745 ( .A1(n27458), .A2(n485), .B1(ram[1575]), .B2(n486), .ZN(
        n5816) );
  MOAI22 U14746 ( .A1(n29103), .A2(n487), .B1(ram[1576]), .B2(n488), .ZN(
        n5817) );
  MOAI22 U14747 ( .A1(n28868), .A2(n487), .B1(ram[1577]), .B2(n488), .ZN(
        n5818) );
  MOAI22 U14748 ( .A1(n28633), .A2(n487), .B1(ram[1578]), .B2(n488), .ZN(
        n5819) );
  MOAI22 U14749 ( .A1(n28398), .A2(n487), .B1(ram[1579]), .B2(n488), .ZN(
        n5820) );
  MOAI22 U14750 ( .A1(n28163), .A2(n487), .B1(ram[1580]), .B2(n488), .ZN(
        n5821) );
  MOAI22 U14751 ( .A1(n27928), .A2(n487), .B1(ram[1581]), .B2(n488), .ZN(
        n5822) );
  MOAI22 U14752 ( .A1(n27693), .A2(n487), .B1(ram[1582]), .B2(n488), .ZN(
        n5823) );
  MOAI22 U14753 ( .A1(n27458), .A2(n487), .B1(ram[1583]), .B2(n488), .ZN(
        n5824) );
  MOAI22 U14754 ( .A1(n29103), .A2(n489), .B1(ram[1584]), .B2(n490), .ZN(
        n5825) );
  MOAI22 U14755 ( .A1(n28868), .A2(n489), .B1(ram[1585]), .B2(n490), .ZN(
        n5826) );
  MOAI22 U14756 ( .A1(n28633), .A2(n489), .B1(ram[1586]), .B2(n490), .ZN(
        n5827) );
  MOAI22 U14757 ( .A1(n28398), .A2(n489), .B1(ram[1587]), .B2(n490), .ZN(
        n5828) );
  MOAI22 U14758 ( .A1(n28163), .A2(n489), .B1(ram[1588]), .B2(n490), .ZN(
        n5829) );
  MOAI22 U14759 ( .A1(n27928), .A2(n489), .B1(ram[1589]), .B2(n490), .ZN(
        n5830) );
  MOAI22 U14760 ( .A1(n27693), .A2(n489), .B1(ram[1590]), .B2(n490), .ZN(
        n5831) );
  MOAI22 U14761 ( .A1(n27458), .A2(n489), .B1(ram[1591]), .B2(n490), .ZN(
        n5832) );
  MOAI22 U14762 ( .A1(n29103), .A2(n491), .B1(ram[1592]), .B2(n492), .ZN(
        n5833) );
  MOAI22 U14763 ( .A1(n28868), .A2(n491), .B1(ram[1593]), .B2(n492), .ZN(
        n5834) );
  MOAI22 U14764 ( .A1(n28633), .A2(n491), .B1(ram[1594]), .B2(n492), .ZN(
        n5835) );
  MOAI22 U14765 ( .A1(n28398), .A2(n491), .B1(ram[1595]), .B2(n492), .ZN(
        n5836) );
  MOAI22 U14766 ( .A1(n28163), .A2(n491), .B1(ram[1596]), .B2(n492), .ZN(
        n5837) );
  MOAI22 U14767 ( .A1(n27928), .A2(n491), .B1(ram[1597]), .B2(n492), .ZN(
        n5838) );
  MOAI22 U14768 ( .A1(n27693), .A2(n491), .B1(ram[1598]), .B2(n492), .ZN(
        n5839) );
  MOAI22 U14769 ( .A1(n27458), .A2(n491), .B1(ram[1599]), .B2(n492), .ZN(
        n5840) );
  MOAI22 U14770 ( .A1(n29103), .A2(n493), .B1(ram[1600]), .B2(n494), .ZN(
        n5841) );
  MOAI22 U14771 ( .A1(n28868), .A2(n493), .B1(ram[1601]), .B2(n494), .ZN(
        n5842) );
  MOAI22 U14772 ( .A1(n28633), .A2(n493), .B1(ram[1602]), .B2(n494), .ZN(
        n5843) );
  MOAI22 U14773 ( .A1(n28398), .A2(n493), .B1(ram[1603]), .B2(n494), .ZN(
        n5844) );
  MOAI22 U14774 ( .A1(n28163), .A2(n493), .B1(ram[1604]), .B2(n494), .ZN(
        n5845) );
  MOAI22 U14775 ( .A1(n27928), .A2(n493), .B1(ram[1605]), .B2(n494), .ZN(
        n5846) );
  MOAI22 U14776 ( .A1(n27693), .A2(n493), .B1(ram[1606]), .B2(n494), .ZN(
        n5847) );
  MOAI22 U14777 ( .A1(n27458), .A2(n493), .B1(ram[1607]), .B2(n494), .ZN(
        n5848) );
  MOAI22 U14778 ( .A1(n29103), .A2(n495), .B1(ram[1608]), .B2(n496), .ZN(
        n5849) );
  MOAI22 U14779 ( .A1(n28868), .A2(n495), .B1(ram[1609]), .B2(n496), .ZN(
        n5850) );
  MOAI22 U14780 ( .A1(n28633), .A2(n495), .B1(ram[1610]), .B2(n496), .ZN(
        n5851) );
  MOAI22 U14781 ( .A1(n28398), .A2(n495), .B1(ram[1611]), .B2(n496), .ZN(
        n5852) );
  MOAI22 U14782 ( .A1(n28163), .A2(n495), .B1(ram[1612]), .B2(n496), .ZN(
        n5853) );
  MOAI22 U14783 ( .A1(n27928), .A2(n495), .B1(ram[1613]), .B2(n496), .ZN(
        n5854) );
  MOAI22 U14784 ( .A1(n27693), .A2(n495), .B1(ram[1614]), .B2(n496), .ZN(
        n5855) );
  MOAI22 U14785 ( .A1(n27458), .A2(n495), .B1(ram[1615]), .B2(n496), .ZN(
        n5856) );
  MOAI22 U14786 ( .A1(n29103), .A2(n497), .B1(ram[1616]), .B2(n498), .ZN(
        n5857) );
  MOAI22 U14787 ( .A1(n28868), .A2(n497), .B1(ram[1617]), .B2(n498), .ZN(
        n5858) );
  MOAI22 U14788 ( .A1(n28633), .A2(n497), .B1(ram[1618]), .B2(n498), .ZN(
        n5859) );
  MOAI22 U14789 ( .A1(n28398), .A2(n497), .B1(ram[1619]), .B2(n498), .ZN(
        n5860) );
  MOAI22 U14790 ( .A1(n28163), .A2(n497), .B1(ram[1620]), .B2(n498), .ZN(
        n5861) );
  MOAI22 U14791 ( .A1(n27928), .A2(n497), .B1(ram[1621]), .B2(n498), .ZN(
        n5862) );
  MOAI22 U14792 ( .A1(n27693), .A2(n497), .B1(ram[1622]), .B2(n498), .ZN(
        n5863) );
  MOAI22 U14793 ( .A1(n27458), .A2(n497), .B1(ram[1623]), .B2(n498), .ZN(
        n5864) );
  MOAI22 U14794 ( .A1(n29103), .A2(n499), .B1(ram[1624]), .B2(n500), .ZN(
        n5865) );
  MOAI22 U14795 ( .A1(n28868), .A2(n499), .B1(ram[1625]), .B2(n500), .ZN(
        n5866) );
  MOAI22 U14796 ( .A1(n28633), .A2(n499), .B1(ram[1626]), .B2(n500), .ZN(
        n5867) );
  MOAI22 U14797 ( .A1(n28398), .A2(n499), .B1(ram[1627]), .B2(n500), .ZN(
        n5868) );
  MOAI22 U14798 ( .A1(n28163), .A2(n499), .B1(ram[1628]), .B2(n500), .ZN(
        n5869) );
  MOAI22 U14799 ( .A1(n27928), .A2(n499), .B1(ram[1629]), .B2(n500), .ZN(
        n5870) );
  MOAI22 U14800 ( .A1(n27693), .A2(n499), .B1(ram[1630]), .B2(n500), .ZN(
        n5871) );
  MOAI22 U14801 ( .A1(n27458), .A2(n499), .B1(ram[1631]), .B2(n500), .ZN(
        n5872) );
  MOAI22 U14802 ( .A1(n29103), .A2(n501), .B1(ram[1632]), .B2(n502), .ZN(
        n5873) );
  MOAI22 U14803 ( .A1(n28868), .A2(n501), .B1(ram[1633]), .B2(n502), .ZN(
        n5874) );
  MOAI22 U14804 ( .A1(n28633), .A2(n501), .B1(ram[1634]), .B2(n502), .ZN(
        n5875) );
  MOAI22 U14805 ( .A1(n28398), .A2(n501), .B1(ram[1635]), .B2(n502), .ZN(
        n5876) );
  MOAI22 U14806 ( .A1(n28163), .A2(n501), .B1(ram[1636]), .B2(n502), .ZN(
        n5877) );
  MOAI22 U14807 ( .A1(n27928), .A2(n501), .B1(ram[1637]), .B2(n502), .ZN(
        n5878) );
  MOAI22 U14808 ( .A1(n27693), .A2(n501), .B1(ram[1638]), .B2(n502), .ZN(
        n5879) );
  MOAI22 U14809 ( .A1(n27458), .A2(n501), .B1(ram[1639]), .B2(n502), .ZN(
        n5880) );
  MOAI22 U14810 ( .A1(n29103), .A2(n503), .B1(ram[1640]), .B2(n504), .ZN(
        n5881) );
  MOAI22 U14811 ( .A1(n28868), .A2(n503), .B1(ram[1641]), .B2(n504), .ZN(
        n5882) );
  MOAI22 U14812 ( .A1(n28633), .A2(n503), .B1(ram[1642]), .B2(n504), .ZN(
        n5883) );
  MOAI22 U14813 ( .A1(n28398), .A2(n503), .B1(ram[1643]), .B2(n504), .ZN(
        n5884) );
  MOAI22 U14814 ( .A1(n28163), .A2(n503), .B1(ram[1644]), .B2(n504), .ZN(
        n5885) );
  MOAI22 U14815 ( .A1(n27928), .A2(n503), .B1(ram[1645]), .B2(n504), .ZN(
        n5886) );
  MOAI22 U14816 ( .A1(n27693), .A2(n503), .B1(ram[1646]), .B2(n504), .ZN(
        n5887) );
  MOAI22 U14817 ( .A1(n27458), .A2(n503), .B1(ram[1647]), .B2(n504), .ZN(
        n5888) );
  MOAI22 U14818 ( .A1(n29103), .A2(n505), .B1(ram[1648]), .B2(n506), .ZN(
        n5889) );
  MOAI22 U14819 ( .A1(n28868), .A2(n505), .B1(ram[1649]), .B2(n506), .ZN(
        n5890) );
  MOAI22 U14820 ( .A1(n28633), .A2(n505), .B1(ram[1650]), .B2(n506), .ZN(
        n5891) );
  MOAI22 U14821 ( .A1(n28398), .A2(n505), .B1(ram[1651]), .B2(n506), .ZN(
        n5892) );
  MOAI22 U14822 ( .A1(n28163), .A2(n505), .B1(ram[1652]), .B2(n506), .ZN(
        n5893) );
  MOAI22 U14823 ( .A1(n27928), .A2(n505), .B1(ram[1653]), .B2(n506), .ZN(
        n5894) );
  MOAI22 U14824 ( .A1(n27693), .A2(n505), .B1(ram[1654]), .B2(n506), .ZN(
        n5895) );
  MOAI22 U14825 ( .A1(n27458), .A2(n505), .B1(ram[1655]), .B2(n506), .ZN(
        n5896) );
  MOAI22 U14826 ( .A1(n29103), .A2(n507), .B1(ram[1656]), .B2(n508), .ZN(
        n5897) );
  MOAI22 U14827 ( .A1(n28868), .A2(n507), .B1(ram[1657]), .B2(n508), .ZN(
        n5898) );
  MOAI22 U14828 ( .A1(n28633), .A2(n507), .B1(ram[1658]), .B2(n508), .ZN(
        n5899) );
  MOAI22 U14829 ( .A1(n28398), .A2(n507), .B1(ram[1659]), .B2(n508), .ZN(
        n5900) );
  MOAI22 U14830 ( .A1(n28163), .A2(n507), .B1(ram[1660]), .B2(n508), .ZN(
        n5901) );
  MOAI22 U14831 ( .A1(n27928), .A2(n507), .B1(ram[1661]), .B2(n508), .ZN(
        n5902) );
  MOAI22 U14832 ( .A1(n27693), .A2(n507), .B1(ram[1662]), .B2(n508), .ZN(
        n5903) );
  MOAI22 U14833 ( .A1(n27458), .A2(n507), .B1(ram[1663]), .B2(n508), .ZN(
        n5904) );
  MOAI22 U14834 ( .A1(n29104), .A2(n509), .B1(ram[1664]), .B2(n510), .ZN(
        n5905) );
  MOAI22 U14835 ( .A1(n28869), .A2(n509), .B1(ram[1665]), .B2(n510), .ZN(
        n5906) );
  MOAI22 U14836 ( .A1(n28634), .A2(n509), .B1(ram[1666]), .B2(n510), .ZN(
        n5907) );
  MOAI22 U14837 ( .A1(n28399), .A2(n509), .B1(ram[1667]), .B2(n510), .ZN(
        n5908) );
  MOAI22 U14838 ( .A1(n28164), .A2(n509), .B1(ram[1668]), .B2(n510), .ZN(
        n5909) );
  MOAI22 U14839 ( .A1(n27929), .A2(n509), .B1(ram[1669]), .B2(n510), .ZN(
        n5910) );
  MOAI22 U14840 ( .A1(n27694), .A2(n509), .B1(ram[1670]), .B2(n510), .ZN(
        n5911) );
  MOAI22 U14841 ( .A1(n27459), .A2(n509), .B1(ram[1671]), .B2(n510), .ZN(
        n5912) );
  MOAI22 U14842 ( .A1(n29104), .A2(n511), .B1(ram[1672]), .B2(n512), .ZN(
        n5913) );
  MOAI22 U14843 ( .A1(n28869), .A2(n511), .B1(ram[1673]), .B2(n512), .ZN(
        n5914) );
  MOAI22 U14844 ( .A1(n28634), .A2(n511), .B1(ram[1674]), .B2(n512), .ZN(
        n5915) );
  MOAI22 U14845 ( .A1(n28399), .A2(n511), .B1(ram[1675]), .B2(n512), .ZN(
        n5916) );
  MOAI22 U14846 ( .A1(n28164), .A2(n511), .B1(ram[1676]), .B2(n512), .ZN(
        n5917) );
  MOAI22 U14847 ( .A1(n27929), .A2(n511), .B1(ram[1677]), .B2(n512), .ZN(
        n5918) );
  MOAI22 U14848 ( .A1(n27694), .A2(n511), .B1(ram[1678]), .B2(n512), .ZN(
        n5919) );
  MOAI22 U14849 ( .A1(n27459), .A2(n511), .B1(ram[1679]), .B2(n512), .ZN(
        n5920) );
  MOAI22 U14850 ( .A1(n29104), .A2(n513), .B1(ram[1680]), .B2(n514), .ZN(
        n5921) );
  MOAI22 U14851 ( .A1(n28869), .A2(n513), .B1(ram[1681]), .B2(n514), .ZN(
        n5922) );
  MOAI22 U14852 ( .A1(n28634), .A2(n513), .B1(ram[1682]), .B2(n514), .ZN(
        n5923) );
  MOAI22 U14853 ( .A1(n28399), .A2(n513), .B1(ram[1683]), .B2(n514), .ZN(
        n5924) );
  MOAI22 U14854 ( .A1(n28164), .A2(n513), .B1(ram[1684]), .B2(n514), .ZN(
        n5925) );
  MOAI22 U14855 ( .A1(n27929), .A2(n513), .B1(ram[1685]), .B2(n514), .ZN(
        n5926) );
  MOAI22 U14856 ( .A1(n27694), .A2(n513), .B1(ram[1686]), .B2(n514), .ZN(
        n5927) );
  MOAI22 U14857 ( .A1(n27459), .A2(n513), .B1(ram[1687]), .B2(n514), .ZN(
        n5928) );
  MOAI22 U14858 ( .A1(n29104), .A2(n515), .B1(ram[1688]), .B2(n516), .ZN(
        n5929) );
  MOAI22 U14859 ( .A1(n28869), .A2(n515), .B1(ram[1689]), .B2(n516), .ZN(
        n5930) );
  MOAI22 U14860 ( .A1(n28634), .A2(n515), .B1(ram[1690]), .B2(n516), .ZN(
        n5931) );
  MOAI22 U14861 ( .A1(n28399), .A2(n515), .B1(ram[1691]), .B2(n516), .ZN(
        n5932) );
  MOAI22 U14862 ( .A1(n28164), .A2(n515), .B1(ram[1692]), .B2(n516), .ZN(
        n5933) );
  MOAI22 U14863 ( .A1(n27929), .A2(n515), .B1(ram[1693]), .B2(n516), .ZN(
        n5934) );
  MOAI22 U14864 ( .A1(n27694), .A2(n515), .B1(ram[1694]), .B2(n516), .ZN(
        n5935) );
  MOAI22 U14865 ( .A1(n27459), .A2(n515), .B1(ram[1695]), .B2(n516), .ZN(
        n5936) );
  MOAI22 U14866 ( .A1(n29104), .A2(n517), .B1(ram[1696]), .B2(n518), .ZN(
        n5937) );
  MOAI22 U14867 ( .A1(n28869), .A2(n517), .B1(ram[1697]), .B2(n518), .ZN(
        n5938) );
  MOAI22 U14868 ( .A1(n28634), .A2(n517), .B1(ram[1698]), .B2(n518), .ZN(
        n5939) );
  MOAI22 U14869 ( .A1(n28399), .A2(n517), .B1(ram[1699]), .B2(n518), .ZN(
        n5940) );
  MOAI22 U14870 ( .A1(n28164), .A2(n517), .B1(ram[1700]), .B2(n518), .ZN(
        n5941) );
  MOAI22 U14871 ( .A1(n27929), .A2(n517), .B1(ram[1701]), .B2(n518), .ZN(
        n5942) );
  MOAI22 U14872 ( .A1(n27694), .A2(n517), .B1(ram[1702]), .B2(n518), .ZN(
        n5943) );
  MOAI22 U14873 ( .A1(n27459), .A2(n517), .B1(ram[1703]), .B2(n518), .ZN(
        n5944) );
  MOAI22 U14874 ( .A1(n29104), .A2(n519), .B1(ram[1704]), .B2(n520), .ZN(
        n5945) );
  MOAI22 U14875 ( .A1(n28869), .A2(n519), .B1(ram[1705]), .B2(n520), .ZN(
        n5946) );
  MOAI22 U14876 ( .A1(n28634), .A2(n519), .B1(ram[1706]), .B2(n520), .ZN(
        n5947) );
  MOAI22 U14877 ( .A1(n28399), .A2(n519), .B1(ram[1707]), .B2(n520), .ZN(
        n5948) );
  MOAI22 U14878 ( .A1(n28164), .A2(n519), .B1(ram[1708]), .B2(n520), .ZN(
        n5949) );
  MOAI22 U14879 ( .A1(n27929), .A2(n519), .B1(ram[1709]), .B2(n520), .ZN(
        n5950) );
  MOAI22 U14880 ( .A1(n27694), .A2(n519), .B1(ram[1710]), .B2(n520), .ZN(
        n5951) );
  MOAI22 U14881 ( .A1(n27459), .A2(n519), .B1(ram[1711]), .B2(n520), .ZN(
        n5952) );
  MOAI22 U14882 ( .A1(n29104), .A2(n521), .B1(ram[1712]), .B2(n522), .ZN(
        n5953) );
  MOAI22 U14883 ( .A1(n28869), .A2(n521), .B1(ram[1713]), .B2(n522), .ZN(
        n5954) );
  MOAI22 U14884 ( .A1(n28634), .A2(n521), .B1(ram[1714]), .B2(n522), .ZN(
        n5955) );
  MOAI22 U14885 ( .A1(n28399), .A2(n521), .B1(ram[1715]), .B2(n522), .ZN(
        n5956) );
  MOAI22 U14886 ( .A1(n28164), .A2(n521), .B1(ram[1716]), .B2(n522), .ZN(
        n5957) );
  MOAI22 U14887 ( .A1(n27929), .A2(n521), .B1(ram[1717]), .B2(n522), .ZN(
        n5958) );
  MOAI22 U14888 ( .A1(n27694), .A2(n521), .B1(ram[1718]), .B2(n522), .ZN(
        n5959) );
  MOAI22 U14889 ( .A1(n27459), .A2(n521), .B1(ram[1719]), .B2(n522), .ZN(
        n5960) );
  MOAI22 U14890 ( .A1(n29104), .A2(n523), .B1(ram[1720]), .B2(n524), .ZN(
        n5961) );
  MOAI22 U14891 ( .A1(n28869), .A2(n523), .B1(ram[1721]), .B2(n524), .ZN(
        n5962) );
  MOAI22 U14892 ( .A1(n28634), .A2(n523), .B1(ram[1722]), .B2(n524), .ZN(
        n5963) );
  MOAI22 U14893 ( .A1(n28399), .A2(n523), .B1(ram[1723]), .B2(n524), .ZN(
        n5964) );
  MOAI22 U14894 ( .A1(n28164), .A2(n523), .B1(ram[1724]), .B2(n524), .ZN(
        n5965) );
  MOAI22 U14895 ( .A1(n27929), .A2(n523), .B1(ram[1725]), .B2(n524), .ZN(
        n5966) );
  MOAI22 U14896 ( .A1(n27694), .A2(n523), .B1(ram[1726]), .B2(n524), .ZN(
        n5967) );
  MOAI22 U14897 ( .A1(n27459), .A2(n523), .B1(ram[1727]), .B2(n524), .ZN(
        n5968) );
  MOAI22 U14898 ( .A1(n29104), .A2(n525), .B1(ram[1728]), .B2(n526), .ZN(
        n5969) );
  MOAI22 U14899 ( .A1(n28869), .A2(n525), .B1(ram[1729]), .B2(n526), .ZN(
        n5970) );
  MOAI22 U14900 ( .A1(n28634), .A2(n525), .B1(ram[1730]), .B2(n526), .ZN(
        n5971) );
  MOAI22 U14901 ( .A1(n28399), .A2(n525), .B1(ram[1731]), .B2(n526), .ZN(
        n5972) );
  MOAI22 U14902 ( .A1(n28164), .A2(n525), .B1(ram[1732]), .B2(n526), .ZN(
        n5973) );
  MOAI22 U14903 ( .A1(n27929), .A2(n525), .B1(ram[1733]), .B2(n526), .ZN(
        n5974) );
  MOAI22 U14904 ( .A1(n27694), .A2(n525), .B1(ram[1734]), .B2(n526), .ZN(
        n5975) );
  MOAI22 U14905 ( .A1(n27459), .A2(n525), .B1(ram[1735]), .B2(n526), .ZN(
        n5976) );
  MOAI22 U14906 ( .A1(n29104), .A2(n527), .B1(ram[1736]), .B2(n528), .ZN(
        n5977) );
  MOAI22 U14907 ( .A1(n28869), .A2(n527), .B1(ram[1737]), .B2(n528), .ZN(
        n5978) );
  MOAI22 U14908 ( .A1(n28634), .A2(n527), .B1(ram[1738]), .B2(n528), .ZN(
        n5979) );
  MOAI22 U14909 ( .A1(n28399), .A2(n527), .B1(ram[1739]), .B2(n528), .ZN(
        n5980) );
  MOAI22 U14910 ( .A1(n28164), .A2(n527), .B1(ram[1740]), .B2(n528), .ZN(
        n5981) );
  MOAI22 U14911 ( .A1(n27929), .A2(n527), .B1(ram[1741]), .B2(n528), .ZN(
        n5982) );
  MOAI22 U14912 ( .A1(n27694), .A2(n527), .B1(ram[1742]), .B2(n528), .ZN(
        n5983) );
  MOAI22 U14913 ( .A1(n27459), .A2(n527), .B1(ram[1743]), .B2(n528), .ZN(
        n5984) );
  MOAI22 U14914 ( .A1(n29104), .A2(n529), .B1(ram[1744]), .B2(n530), .ZN(
        n5985) );
  MOAI22 U14915 ( .A1(n28869), .A2(n529), .B1(ram[1745]), .B2(n530), .ZN(
        n5986) );
  MOAI22 U14916 ( .A1(n28634), .A2(n529), .B1(ram[1746]), .B2(n530), .ZN(
        n5987) );
  MOAI22 U14917 ( .A1(n28399), .A2(n529), .B1(ram[1747]), .B2(n530), .ZN(
        n5988) );
  MOAI22 U14918 ( .A1(n28164), .A2(n529), .B1(ram[1748]), .B2(n530), .ZN(
        n5989) );
  MOAI22 U14919 ( .A1(n27929), .A2(n529), .B1(ram[1749]), .B2(n530), .ZN(
        n5990) );
  MOAI22 U14920 ( .A1(n27694), .A2(n529), .B1(ram[1750]), .B2(n530), .ZN(
        n5991) );
  MOAI22 U14921 ( .A1(n27459), .A2(n529), .B1(ram[1751]), .B2(n530), .ZN(
        n5992) );
  MOAI22 U14922 ( .A1(n29104), .A2(n531), .B1(ram[1752]), .B2(n532), .ZN(
        n5993) );
  MOAI22 U14923 ( .A1(n28869), .A2(n531), .B1(ram[1753]), .B2(n532), .ZN(
        n5994) );
  MOAI22 U14924 ( .A1(n28634), .A2(n531), .B1(ram[1754]), .B2(n532), .ZN(
        n5995) );
  MOAI22 U14925 ( .A1(n28399), .A2(n531), .B1(ram[1755]), .B2(n532), .ZN(
        n5996) );
  MOAI22 U14926 ( .A1(n28164), .A2(n531), .B1(ram[1756]), .B2(n532), .ZN(
        n5997) );
  MOAI22 U14927 ( .A1(n27929), .A2(n531), .B1(ram[1757]), .B2(n532), .ZN(
        n5998) );
  MOAI22 U14928 ( .A1(n27694), .A2(n531), .B1(ram[1758]), .B2(n532), .ZN(
        n5999) );
  MOAI22 U14929 ( .A1(n27459), .A2(n531), .B1(ram[1759]), .B2(n532), .ZN(
        n6000) );
  MOAI22 U14930 ( .A1(n29104), .A2(n533), .B1(ram[1760]), .B2(n534), .ZN(
        n6001) );
  MOAI22 U14931 ( .A1(n28869), .A2(n533), .B1(ram[1761]), .B2(n534), .ZN(
        n6002) );
  MOAI22 U14932 ( .A1(n28634), .A2(n533), .B1(ram[1762]), .B2(n534), .ZN(
        n6003) );
  MOAI22 U14933 ( .A1(n28399), .A2(n533), .B1(ram[1763]), .B2(n534), .ZN(
        n6004) );
  MOAI22 U14934 ( .A1(n28164), .A2(n533), .B1(ram[1764]), .B2(n534), .ZN(
        n6005) );
  MOAI22 U14935 ( .A1(n27929), .A2(n533), .B1(ram[1765]), .B2(n534), .ZN(
        n6006) );
  MOAI22 U14936 ( .A1(n27694), .A2(n533), .B1(ram[1766]), .B2(n534), .ZN(
        n6007) );
  MOAI22 U14937 ( .A1(n27459), .A2(n533), .B1(ram[1767]), .B2(n534), .ZN(
        n6008) );
  MOAI22 U14938 ( .A1(n29105), .A2(n535), .B1(ram[1768]), .B2(n536), .ZN(
        n6009) );
  MOAI22 U14939 ( .A1(n28870), .A2(n535), .B1(ram[1769]), .B2(n536), .ZN(
        n6010) );
  MOAI22 U14940 ( .A1(n28635), .A2(n535), .B1(ram[1770]), .B2(n536), .ZN(
        n6011) );
  MOAI22 U14941 ( .A1(n28400), .A2(n535), .B1(ram[1771]), .B2(n536), .ZN(
        n6012) );
  MOAI22 U14942 ( .A1(n28165), .A2(n535), .B1(ram[1772]), .B2(n536), .ZN(
        n6013) );
  MOAI22 U14943 ( .A1(n27930), .A2(n535), .B1(ram[1773]), .B2(n536), .ZN(
        n6014) );
  MOAI22 U14944 ( .A1(n27695), .A2(n535), .B1(ram[1774]), .B2(n536), .ZN(
        n6015) );
  MOAI22 U14945 ( .A1(n27460), .A2(n535), .B1(ram[1775]), .B2(n536), .ZN(
        n6016) );
  MOAI22 U14946 ( .A1(n29105), .A2(n537), .B1(ram[1776]), .B2(n538), .ZN(
        n6017) );
  MOAI22 U14947 ( .A1(n28870), .A2(n537), .B1(ram[1777]), .B2(n538), .ZN(
        n6018) );
  MOAI22 U14948 ( .A1(n28635), .A2(n537), .B1(ram[1778]), .B2(n538), .ZN(
        n6019) );
  MOAI22 U14949 ( .A1(n28400), .A2(n537), .B1(ram[1779]), .B2(n538), .ZN(
        n6020) );
  MOAI22 U14950 ( .A1(n28165), .A2(n537), .B1(ram[1780]), .B2(n538), .ZN(
        n6021) );
  MOAI22 U14951 ( .A1(n27930), .A2(n537), .B1(ram[1781]), .B2(n538), .ZN(
        n6022) );
  MOAI22 U14952 ( .A1(n27695), .A2(n537), .B1(ram[1782]), .B2(n538), .ZN(
        n6023) );
  MOAI22 U14953 ( .A1(n27460), .A2(n537), .B1(ram[1783]), .B2(n538), .ZN(
        n6024) );
  MOAI22 U14954 ( .A1(n29105), .A2(n539), .B1(ram[1784]), .B2(n540), .ZN(
        n6025) );
  MOAI22 U14955 ( .A1(n28870), .A2(n539), .B1(ram[1785]), .B2(n540), .ZN(
        n6026) );
  MOAI22 U14956 ( .A1(n28635), .A2(n539), .B1(ram[1786]), .B2(n540), .ZN(
        n6027) );
  MOAI22 U14957 ( .A1(n28400), .A2(n539), .B1(ram[1787]), .B2(n540), .ZN(
        n6028) );
  MOAI22 U14958 ( .A1(n28165), .A2(n539), .B1(ram[1788]), .B2(n540), .ZN(
        n6029) );
  MOAI22 U14959 ( .A1(n27930), .A2(n539), .B1(ram[1789]), .B2(n540), .ZN(
        n6030) );
  MOAI22 U14960 ( .A1(n27695), .A2(n539), .B1(ram[1790]), .B2(n540), .ZN(
        n6031) );
  MOAI22 U14961 ( .A1(n27460), .A2(n539), .B1(ram[1791]), .B2(n540), .ZN(
        n6032) );
  MOAI22 U14962 ( .A1(n29105), .A2(n541), .B1(ram[1792]), .B2(n542), .ZN(
        n6033) );
  MOAI22 U14963 ( .A1(n28870), .A2(n541), .B1(ram[1793]), .B2(n542), .ZN(
        n6034) );
  MOAI22 U14964 ( .A1(n28635), .A2(n541), .B1(ram[1794]), .B2(n542), .ZN(
        n6035) );
  MOAI22 U14965 ( .A1(n28400), .A2(n541), .B1(ram[1795]), .B2(n542), .ZN(
        n6036) );
  MOAI22 U14966 ( .A1(n28165), .A2(n541), .B1(ram[1796]), .B2(n542), .ZN(
        n6037) );
  MOAI22 U14967 ( .A1(n27930), .A2(n541), .B1(ram[1797]), .B2(n542), .ZN(
        n6038) );
  MOAI22 U14968 ( .A1(n27695), .A2(n541), .B1(ram[1798]), .B2(n542), .ZN(
        n6039) );
  MOAI22 U14969 ( .A1(n27460), .A2(n541), .B1(ram[1799]), .B2(n542), .ZN(
        n6040) );
  MOAI22 U14970 ( .A1(n29105), .A2(n543), .B1(ram[1800]), .B2(n544), .ZN(
        n6041) );
  MOAI22 U14971 ( .A1(n28870), .A2(n543), .B1(ram[1801]), .B2(n544), .ZN(
        n6042) );
  MOAI22 U14972 ( .A1(n28635), .A2(n543), .B1(ram[1802]), .B2(n544), .ZN(
        n6043) );
  MOAI22 U14973 ( .A1(n28400), .A2(n543), .B1(ram[1803]), .B2(n544), .ZN(
        n6044) );
  MOAI22 U14974 ( .A1(n28165), .A2(n543), .B1(ram[1804]), .B2(n544), .ZN(
        n6045) );
  MOAI22 U14975 ( .A1(n27930), .A2(n543), .B1(ram[1805]), .B2(n544), .ZN(
        n6046) );
  MOAI22 U14976 ( .A1(n27695), .A2(n543), .B1(ram[1806]), .B2(n544), .ZN(
        n6047) );
  MOAI22 U14977 ( .A1(n27460), .A2(n543), .B1(ram[1807]), .B2(n544), .ZN(
        n6048) );
  MOAI22 U14978 ( .A1(n29105), .A2(n545), .B1(ram[1808]), .B2(n546), .ZN(
        n6049) );
  MOAI22 U14979 ( .A1(n28870), .A2(n545), .B1(ram[1809]), .B2(n546), .ZN(
        n6050) );
  MOAI22 U14980 ( .A1(n28635), .A2(n545), .B1(ram[1810]), .B2(n546), .ZN(
        n6051) );
  MOAI22 U14981 ( .A1(n28400), .A2(n545), .B1(ram[1811]), .B2(n546), .ZN(
        n6052) );
  MOAI22 U14982 ( .A1(n28165), .A2(n545), .B1(ram[1812]), .B2(n546), .ZN(
        n6053) );
  MOAI22 U14983 ( .A1(n27930), .A2(n545), .B1(ram[1813]), .B2(n546), .ZN(
        n6054) );
  MOAI22 U14984 ( .A1(n27695), .A2(n545), .B1(ram[1814]), .B2(n546), .ZN(
        n6055) );
  MOAI22 U14985 ( .A1(n27460), .A2(n545), .B1(ram[1815]), .B2(n546), .ZN(
        n6056) );
  MOAI22 U14986 ( .A1(n29105), .A2(n547), .B1(ram[1816]), .B2(n548), .ZN(
        n6057) );
  MOAI22 U14987 ( .A1(n28870), .A2(n547), .B1(ram[1817]), .B2(n548), .ZN(
        n6058) );
  MOAI22 U14988 ( .A1(n28635), .A2(n547), .B1(ram[1818]), .B2(n548), .ZN(
        n6059) );
  MOAI22 U14989 ( .A1(n28400), .A2(n547), .B1(ram[1819]), .B2(n548), .ZN(
        n6060) );
  MOAI22 U14990 ( .A1(n28165), .A2(n547), .B1(ram[1820]), .B2(n548), .ZN(
        n6061) );
  MOAI22 U14991 ( .A1(n27930), .A2(n547), .B1(ram[1821]), .B2(n548), .ZN(
        n6062) );
  MOAI22 U14992 ( .A1(n27695), .A2(n547), .B1(ram[1822]), .B2(n548), .ZN(
        n6063) );
  MOAI22 U14993 ( .A1(n27460), .A2(n547), .B1(ram[1823]), .B2(n548), .ZN(
        n6064) );
  MOAI22 U14994 ( .A1(n29105), .A2(n549), .B1(ram[1824]), .B2(n550), .ZN(
        n6065) );
  MOAI22 U14995 ( .A1(n28870), .A2(n549), .B1(ram[1825]), .B2(n550), .ZN(
        n6066) );
  MOAI22 U14996 ( .A1(n28635), .A2(n549), .B1(ram[1826]), .B2(n550), .ZN(
        n6067) );
  MOAI22 U14997 ( .A1(n28400), .A2(n549), .B1(ram[1827]), .B2(n550), .ZN(
        n6068) );
  MOAI22 U14998 ( .A1(n28165), .A2(n549), .B1(ram[1828]), .B2(n550), .ZN(
        n6069) );
  MOAI22 U14999 ( .A1(n27930), .A2(n549), .B1(ram[1829]), .B2(n550), .ZN(
        n6070) );
  MOAI22 U15000 ( .A1(n27695), .A2(n549), .B1(ram[1830]), .B2(n550), .ZN(
        n6071) );
  MOAI22 U15001 ( .A1(n27460), .A2(n549), .B1(ram[1831]), .B2(n550), .ZN(
        n6072) );
  MOAI22 U15002 ( .A1(n29105), .A2(n551), .B1(ram[1832]), .B2(n552), .ZN(
        n6073) );
  MOAI22 U15003 ( .A1(n28870), .A2(n551), .B1(ram[1833]), .B2(n552), .ZN(
        n6074) );
  MOAI22 U15004 ( .A1(n28635), .A2(n551), .B1(ram[1834]), .B2(n552), .ZN(
        n6075) );
  MOAI22 U15005 ( .A1(n28400), .A2(n551), .B1(ram[1835]), .B2(n552), .ZN(
        n6076) );
  MOAI22 U15006 ( .A1(n28165), .A2(n551), .B1(ram[1836]), .B2(n552), .ZN(
        n6077) );
  MOAI22 U15007 ( .A1(n27930), .A2(n551), .B1(ram[1837]), .B2(n552), .ZN(
        n6078) );
  MOAI22 U15008 ( .A1(n27695), .A2(n551), .B1(ram[1838]), .B2(n552), .ZN(
        n6079) );
  MOAI22 U15009 ( .A1(n27460), .A2(n551), .B1(ram[1839]), .B2(n552), .ZN(
        n6080) );
  MOAI22 U15010 ( .A1(n29105), .A2(n553), .B1(ram[1840]), .B2(n554), .ZN(
        n6081) );
  MOAI22 U15011 ( .A1(n28870), .A2(n553), .B1(ram[1841]), .B2(n554), .ZN(
        n6082) );
  MOAI22 U15012 ( .A1(n28635), .A2(n553), .B1(ram[1842]), .B2(n554), .ZN(
        n6083) );
  MOAI22 U15013 ( .A1(n28400), .A2(n553), .B1(ram[1843]), .B2(n554), .ZN(
        n6084) );
  MOAI22 U15014 ( .A1(n28165), .A2(n553), .B1(ram[1844]), .B2(n554), .ZN(
        n6085) );
  MOAI22 U15015 ( .A1(n27930), .A2(n553), .B1(ram[1845]), .B2(n554), .ZN(
        n6086) );
  MOAI22 U15016 ( .A1(n27695), .A2(n553), .B1(ram[1846]), .B2(n554), .ZN(
        n6087) );
  MOAI22 U15017 ( .A1(n27460), .A2(n553), .B1(ram[1847]), .B2(n554), .ZN(
        n6088) );
  MOAI22 U15018 ( .A1(n29105), .A2(n555), .B1(ram[1848]), .B2(n556), .ZN(
        n6089) );
  MOAI22 U15019 ( .A1(n28870), .A2(n555), .B1(ram[1849]), .B2(n556), .ZN(
        n6090) );
  MOAI22 U15020 ( .A1(n28635), .A2(n555), .B1(ram[1850]), .B2(n556), .ZN(
        n6091) );
  MOAI22 U15021 ( .A1(n28400), .A2(n555), .B1(ram[1851]), .B2(n556), .ZN(
        n6092) );
  MOAI22 U15022 ( .A1(n28165), .A2(n555), .B1(ram[1852]), .B2(n556), .ZN(
        n6093) );
  MOAI22 U15023 ( .A1(n27930), .A2(n555), .B1(ram[1853]), .B2(n556), .ZN(
        n6094) );
  MOAI22 U15024 ( .A1(n27695), .A2(n555), .B1(ram[1854]), .B2(n556), .ZN(
        n6095) );
  MOAI22 U15025 ( .A1(n27460), .A2(n555), .B1(ram[1855]), .B2(n556), .ZN(
        n6096) );
  MOAI22 U15026 ( .A1(n29105), .A2(n557), .B1(ram[1856]), .B2(n558), .ZN(
        n6097) );
  MOAI22 U15027 ( .A1(n28870), .A2(n557), .B1(ram[1857]), .B2(n558), .ZN(
        n6098) );
  MOAI22 U15028 ( .A1(n28635), .A2(n557), .B1(ram[1858]), .B2(n558), .ZN(
        n6099) );
  MOAI22 U15029 ( .A1(n28400), .A2(n557), .B1(ram[1859]), .B2(n558), .ZN(
        n6100) );
  MOAI22 U15030 ( .A1(n28165), .A2(n557), .B1(ram[1860]), .B2(n558), .ZN(
        n6101) );
  MOAI22 U15031 ( .A1(n27930), .A2(n557), .B1(ram[1861]), .B2(n558), .ZN(
        n6102) );
  MOAI22 U15032 ( .A1(n27695), .A2(n557), .B1(ram[1862]), .B2(n558), .ZN(
        n6103) );
  MOAI22 U15033 ( .A1(n27460), .A2(n557), .B1(ram[1863]), .B2(n558), .ZN(
        n6104) );
  MOAI22 U15034 ( .A1(n29105), .A2(n559), .B1(ram[1864]), .B2(n560), .ZN(
        n6105) );
  MOAI22 U15035 ( .A1(n28870), .A2(n559), .B1(ram[1865]), .B2(n560), .ZN(
        n6106) );
  MOAI22 U15036 ( .A1(n28635), .A2(n559), .B1(ram[1866]), .B2(n560), .ZN(
        n6107) );
  MOAI22 U15037 ( .A1(n28400), .A2(n559), .B1(ram[1867]), .B2(n560), .ZN(
        n6108) );
  MOAI22 U15038 ( .A1(n28165), .A2(n559), .B1(ram[1868]), .B2(n560), .ZN(
        n6109) );
  MOAI22 U15039 ( .A1(n27930), .A2(n559), .B1(ram[1869]), .B2(n560), .ZN(
        n6110) );
  MOAI22 U15040 ( .A1(n27695), .A2(n559), .B1(ram[1870]), .B2(n560), .ZN(
        n6111) );
  MOAI22 U15041 ( .A1(n27460), .A2(n559), .B1(ram[1871]), .B2(n560), .ZN(
        n6112) );
  MOAI22 U15042 ( .A1(n29106), .A2(n561), .B1(ram[1872]), .B2(n562), .ZN(
        n6113) );
  MOAI22 U15043 ( .A1(n28871), .A2(n561), .B1(ram[1873]), .B2(n562), .ZN(
        n6114) );
  MOAI22 U15044 ( .A1(n28636), .A2(n561), .B1(ram[1874]), .B2(n562), .ZN(
        n6115) );
  MOAI22 U15045 ( .A1(n28401), .A2(n561), .B1(ram[1875]), .B2(n562), .ZN(
        n6116) );
  MOAI22 U15046 ( .A1(n28166), .A2(n561), .B1(ram[1876]), .B2(n562), .ZN(
        n6117) );
  MOAI22 U15047 ( .A1(n27931), .A2(n561), .B1(ram[1877]), .B2(n562), .ZN(
        n6118) );
  MOAI22 U15048 ( .A1(n27696), .A2(n561), .B1(ram[1878]), .B2(n562), .ZN(
        n6119) );
  MOAI22 U15049 ( .A1(n27461), .A2(n561), .B1(ram[1879]), .B2(n562), .ZN(
        n6120) );
  MOAI22 U15050 ( .A1(n29106), .A2(n563), .B1(ram[1880]), .B2(n564), .ZN(
        n6121) );
  MOAI22 U15051 ( .A1(n28871), .A2(n563), .B1(ram[1881]), .B2(n564), .ZN(
        n6122) );
  MOAI22 U15052 ( .A1(n28636), .A2(n563), .B1(ram[1882]), .B2(n564), .ZN(
        n6123) );
  MOAI22 U15053 ( .A1(n28401), .A2(n563), .B1(ram[1883]), .B2(n564), .ZN(
        n6124) );
  MOAI22 U15054 ( .A1(n28166), .A2(n563), .B1(ram[1884]), .B2(n564), .ZN(
        n6125) );
  MOAI22 U15055 ( .A1(n27931), .A2(n563), .B1(ram[1885]), .B2(n564), .ZN(
        n6126) );
  MOAI22 U15056 ( .A1(n27696), .A2(n563), .B1(ram[1886]), .B2(n564), .ZN(
        n6127) );
  MOAI22 U15057 ( .A1(n27461), .A2(n563), .B1(ram[1887]), .B2(n564), .ZN(
        n6128) );
  MOAI22 U15058 ( .A1(n29106), .A2(n565), .B1(ram[1888]), .B2(n566), .ZN(
        n6129) );
  MOAI22 U15059 ( .A1(n28871), .A2(n565), .B1(ram[1889]), .B2(n566), .ZN(
        n6130) );
  MOAI22 U15060 ( .A1(n28636), .A2(n565), .B1(ram[1890]), .B2(n566), .ZN(
        n6131) );
  MOAI22 U15061 ( .A1(n28401), .A2(n565), .B1(ram[1891]), .B2(n566), .ZN(
        n6132) );
  MOAI22 U15062 ( .A1(n28166), .A2(n565), .B1(ram[1892]), .B2(n566), .ZN(
        n6133) );
  MOAI22 U15063 ( .A1(n27931), .A2(n565), .B1(ram[1893]), .B2(n566), .ZN(
        n6134) );
  MOAI22 U15064 ( .A1(n27696), .A2(n565), .B1(ram[1894]), .B2(n566), .ZN(
        n6135) );
  MOAI22 U15065 ( .A1(n27461), .A2(n565), .B1(ram[1895]), .B2(n566), .ZN(
        n6136) );
  MOAI22 U15066 ( .A1(n29106), .A2(n567), .B1(ram[1896]), .B2(n568), .ZN(
        n6137) );
  MOAI22 U15067 ( .A1(n28871), .A2(n567), .B1(ram[1897]), .B2(n568), .ZN(
        n6138) );
  MOAI22 U15068 ( .A1(n28636), .A2(n567), .B1(ram[1898]), .B2(n568), .ZN(
        n6139) );
  MOAI22 U15069 ( .A1(n28401), .A2(n567), .B1(ram[1899]), .B2(n568), .ZN(
        n6140) );
  MOAI22 U15070 ( .A1(n28166), .A2(n567), .B1(ram[1900]), .B2(n568), .ZN(
        n6141) );
  MOAI22 U15071 ( .A1(n27931), .A2(n567), .B1(ram[1901]), .B2(n568), .ZN(
        n6142) );
  MOAI22 U15072 ( .A1(n27696), .A2(n567), .B1(ram[1902]), .B2(n568), .ZN(
        n6143) );
  MOAI22 U15073 ( .A1(n27461), .A2(n567), .B1(ram[1903]), .B2(n568), .ZN(
        n6144) );
  MOAI22 U15074 ( .A1(n29106), .A2(n569), .B1(ram[1904]), .B2(n570), .ZN(
        n6145) );
  MOAI22 U15075 ( .A1(n28871), .A2(n569), .B1(ram[1905]), .B2(n570), .ZN(
        n6146) );
  MOAI22 U15076 ( .A1(n28636), .A2(n569), .B1(ram[1906]), .B2(n570), .ZN(
        n6147) );
  MOAI22 U15077 ( .A1(n28401), .A2(n569), .B1(ram[1907]), .B2(n570), .ZN(
        n6148) );
  MOAI22 U15078 ( .A1(n28166), .A2(n569), .B1(ram[1908]), .B2(n570), .ZN(
        n6149) );
  MOAI22 U15079 ( .A1(n27931), .A2(n569), .B1(ram[1909]), .B2(n570), .ZN(
        n6150) );
  MOAI22 U15080 ( .A1(n27696), .A2(n569), .B1(ram[1910]), .B2(n570), .ZN(
        n6151) );
  MOAI22 U15081 ( .A1(n27461), .A2(n569), .B1(ram[1911]), .B2(n570), .ZN(
        n6152) );
  MOAI22 U15082 ( .A1(n29106), .A2(n571), .B1(ram[1912]), .B2(n572), .ZN(
        n6153) );
  MOAI22 U15083 ( .A1(n28871), .A2(n571), .B1(ram[1913]), .B2(n572), .ZN(
        n6154) );
  MOAI22 U15084 ( .A1(n28636), .A2(n571), .B1(ram[1914]), .B2(n572), .ZN(
        n6155) );
  MOAI22 U15085 ( .A1(n28401), .A2(n571), .B1(ram[1915]), .B2(n572), .ZN(
        n6156) );
  MOAI22 U15086 ( .A1(n28166), .A2(n571), .B1(ram[1916]), .B2(n572), .ZN(
        n6157) );
  MOAI22 U15087 ( .A1(n27931), .A2(n571), .B1(ram[1917]), .B2(n572), .ZN(
        n6158) );
  MOAI22 U15088 ( .A1(n27696), .A2(n571), .B1(ram[1918]), .B2(n572), .ZN(
        n6159) );
  MOAI22 U15089 ( .A1(n27461), .A2(n571), .B1(ram[1919]), .B2(n572), .ZN(
        n6160) );
  MOAI22 U15090 ( .A1(n29106), .A2(n573), .B1(ram[1920]), .B2(n574), .ZN(
        n6161) );
  MOAI22 U15091 ( .A1(n28871), .A2(n573), .B1(ram[1921]), .B2(n574), .ZN(
        n6162) );
  MOAI22 U15092 ( .A1(n28636), .A2(n573), .B1(ram[1922]), .B2(n574), .ZN(
        n6163) );
  MOAI22 U15093 ( .A1(n28401), .A2(n573), .B1(ram[1923]), .B2(n574), .ZN(
        n6164) );
  MOAI22 U15094 ( .A1(n28166), .A2(n573), .B1(ram[1924]), .B2(n574), .ZN(
        n6165) );
  MOAI22 U15095 ( .A1(n27931), .A2(n573), .B1(ram[1925]), .B2(n574), .ZN(
        n6166) );
  MOAI22 U15096 ( .A1(n27696), .A2(n573), .B1(ram[1926]), .B2(n574), .ZN(
        n6167) );
  MOAI22 U15097 ( .A1(n27461), .A2(n573), .B1(ram[1927]), .B2(n574), .ZN(
        n6168) );
  MOAI22 U15098 ( .A1(n29106), .A2(n575), .B1(ram[1928]), .B2(n576), .ZN(
        n6169) );
  MOAI22 U15099 ( .A1(n28871), .A2(n575), .B1(ram[1929]), .B2(n576), .ZN(
        n6170) );
  MOAI22 U15100 ( .A1(n28636), .A2(n575), .B1(ram[1930]), .B2(n576), .ZN(
        n6171) );
  MOAI22 U15101 ( .A1(n28401), .A2(n575), .B1(ram[1931]), .B2(n576), .ZN(
        n6172) );
  MOAI22 U15102 ( .A1(n28166), .A2(n575), .B1(ram[1932]), .B2(n576), .ZN(
        n6173) );
  MOAI22 U15103 ( .A1(n27931), .A2(n575), .B1(ram[1933]), .B2(n576), .ZN(
        n6174) );
  MOAI22 U15104 ( .A1(n27696), .A2(n575), .B1(ram[1934]), .B2(n576), .ZN(
        n6175) );
  MOAI22 U15105 ( .A1(n27461), .A2(n575), .B1(ram[1935]), .B2(n576), .ZN(
        n6176) );
  MOAI22 U15106 ( .A1(n29106), .A2(n577), .B1(ram[1936]), .B2(n578), .ZN(
        n6177) );
  MOAI22 U15107 ( .A1(n28871), .A2(n577), .B1(ram[1937]), .B2(n578), .ZN(
        n6178) );
  MOAI22 U15108 ( .A1(n28636), .A2(n577), .B1(ram[1938]), .B2(n578), .ZN(
        n6179) );
  MOAI22 U15109 ( .A1(n28401), .A2(n577), .B1(ram[1939]), .B2(n578), .ZN(
        n6180) );
  MOAI22 U15110 ( .A1(n28166), .A2(n577), .B1(ram[1940]), .B2(n578), .ZN(
        n6181) );
  MOAI22 U15111 ( .A1(n27931), .A2(n577), .B1(ram[1941]), .B2(n578), .ZN(
        n6182) );
  MOAI22 U15112 ( .A1(n27696), .A2(n577), .B1(ram[1942]), .B2(n578), .ZN(
        n6183) );
  MOAI22 U15113 ( .A1(n27461), .A2(n577), .B1(ram[1943]), .B2(n578), .ZN(
        n6184) );
  MOAI22 U15114 ( .A1(n29106), .A2(n579), .B1(ram[1944]), .B2(n580), .ZN(
        n6185) );
  MOAI22 U15115 ( .A1(n28871), .A2(n579), .B1(ram[1945]), .B2(n580), .ZN(
        n6186) );
  MOAI22 U15116 ( .A1(n28636), .A2(n579), .B1(ram[1946]), .B2(n580), .ZN(
        n6187) );
  MOAI22 U15117 ( .A1(n28401), .A2(n579), .B1(ram[1947]), .B2(n580), .ZN(
        n6188) );
  MOAI22 U15118 ( .A1(n28166), .A2(n579), .B1(ram[1948]), .B2(n580), .ZN(
        n6189) );
  MOAI22 U15119 ( .A1(n27931), .A2(n579), .B1(ram[1949]), .B2(n580), .ZN(
        n6190) );
  MOAI22 U15120 ( .A1(n27696), .A2(n579), .B1(ram[1950]), .B2(n580), .ZN(
        n6191) );
  MOAI22 U15121 ( .A1(n27461), .A2(n579), .B1(ram[1951]), .B2(n580), .ZN(
        n6192) );
  MOAI22 U15122 ( .A1(n29106), .A2(n581), .B1(ram[1952]), .B2(n582), .ZN(
        n6193) );
  MOAI22 U15123 ( .A1(n28871), .A2(n581), .B1(ram[1953]), .B2(n582), .ZN(
        n6194) );
  MOAI22 U15124 ( .A1(n28636), .A2(n581), .B1(ram[1954]), .B2(n582), .ZN(
        n6195) );
  MOAI22 U15125 ( .A1(n28401), .A2(n581), .B1(ram[1955]), .B2(n582), .ZN(
        n6196) );
  MOAI22 U15126 ( .A1(n28166), .A2(n581), .B1(ram[1956]), .B2(n582), .ZN(
        n6197) );
  MOAI22 U15127 ( .A1(n27931), .A2(n581), .B1(ram[1957]), .B2(n582), .ZN(
        n6198) );
  MOAI22 U15128 ( .A1(n27696), .A2(n581), .B1(ram[1958]), .B2(n582), .ZN(
        n6199) );
  MOAI22 U15129 ( .A1(n27461), .A2(n581), .B1(ram[1959]), .B2(n582), .ZN(
        n6200) );
  MOAI22 U15130 ( .A1(n29106), .A2(n583), .B1(ram[1960]), .B2(n584), .ZN(
        n6201) );
  MOAI22 U15131 ( .A1(n28871), .A2(n583), .B1(ram[1961]), .B2(n584), .ZN(
        n6202) );
  MOAI22 U15132 ( .A1(n28636), .A2(n583), .B1(ram[1962]), .B2(n584), .ZN(
        n6203) );
  MOAI22 U15133 ( .A1(n28401), .A2(n583), .B1(ram[1963]), .B2(n584), .ZN(
        n6204) );
  MOAI22 U15134 ( .A1(n28166), .A2(n583), .B1(ram[1964]), .B2(n584), .ZN(
        n6205) );
  MOAI22 U15135 ( .A1(n27931), .A2(n583), .B1(ram[1965]), .B2(n584), .ZN(
        n6206) );
  MOAI22 U15136 ( .A1(n27696), .A2(n583), .B1(ram[1966]), .B2(n584), .ZN(
        n6207) );
  MOAI22 U15137 ( .A1(n27461), .A2(n583), .B1(ram[1967]), .B2(n584), .ZN(
        n6208) );
  MOAI22 U15138 ( .A1(n29106), .A2(n585), .B1(ram[1968]), .B2(n586), .ZN(
        n6209) );
  MOAI22 U15139 ( .A1(n28871), .A2(n585), .B1(ram[1969]), .B2(n586), .ZN(
        n6210) );
  MOAI22 U15140 ( .A1(n28636), .A2(n585), .B1(ram[1970]), .B2(n586), .ZN(
        n6211) );
  MOAI22 U15141 ( .A1(n28401), .A2(n585), .B1(ram[1971]), .B2(n586), .ZN(
        n6212) );
  MOAI22 U15142 ( .A1(n28166), .A2(n585), .B1(ram[1972]), .B2(n586), .ZN(
        n6213) );
  MOAI22 U15143 ( .A1(n27931), .A2(n585), .B1(ram[1973]), .B2(n586), .ZN(
        n6214) );
  MOAI22 U15144 ( .A1(n27696), .A2(n585), .B1(ram[1974]), .B2(n586), .ZN(
        n6215) );
  MOAI22 U15145 ( .A1(n27461), .A2(n585), .B1(ram[1975]), .B2(n586), .ZN(
        n6216) );
  MOAI22 U15146 ( .A1(n29107), .A2(n587), .B1(ram[1976]), .B2(n588), .ZN(
        n6217) );
  MOAI22 U15147 ( .A1(n28872), .A2(n587), .B1(ram[1977]), .B2(n588), .ZN(
        n6218) );
  MOAI22 U15148 ( .A1(n28637), .A2(n587), .B1(ram[1978]), .B2(n588), .ZN(
        n6219) );
  MOAI22 U15149 ( .A1(n28402), .A2(n587), .B1(ram[1979]), .B2(n588), .ZN(
        n6220) );
  MOAI22 U15150 ( .A1(n28167), .A2(n587), .B1(ram[1980]), .B2(n588), .ZN(
        n6221) );
  MOAI22 U15151 ( .A1(n27932), .A2(n587), .B1(ram[1981]), .B2(n588), .ZN(
        n6222) );
  MOAI22 U15152 ( .A1(n27697), .A2(n587), .B1(ram[1982]), .B2(n588), .ZN(
        n6223) );
  MOAI22 U15153 ( .A1(n27462), .A2(n587), .B1(ram[1983]), .B2(n588), .ZN(
        n6224) );
  MOAI22 U15154 ( .A1(n29107), .A2(n589), .B1(ram[1984]), .B2(n590), .ZN(
        n6225) );
  MOAI22 U15155 ( .A1(n28872), .A2(n589), .B1(ram[1985]), .B2(n590), .ZN(
        n6226) );
  MOAI22 U15156 ( .A1(n28637), .A2(n589), .B1(ram[1986]), .B2(n590), .ZN(
        n6227) );
  MOAI22 U15157 ( .A1(n28402), .A2(n589), .B1(ram[1987]), .B2(n590), .ZN(
        n6228) );
  MOAI22 U15158 ( .A1(n28167), .A2(n589), .B1(ram[1988]), .B2(n590), .ZN(
        n6229) );
  MOAI22 U15159 ( .A1(n27932), .A2(n589), .B1(ram[1989]), .B2(n590), .ZN(
        n6230) );
  MOAI22 U15160 ( .A1(n27697), .A2(n589), .B1(ram[1990]), .B2(n590), .ZN(
        n6231) );
  MOAI22 U15161 ( .A1(n27462), .A2(n589), .B1(ram[1991]), .B2(n590), .ZN(
        n6232) );
  MOAI22 U15162 ( .A1(n29107), .A2(n591), .B1(ram[1992]), .B2(n592), .ZN(
        n6233) );
  MOAI22 U15163 ( .A1(n28872), .A2(n591), .B1(ram[1993]), .B2(n592), .ZN(
        n6234) );
  MOAI22 U15164 ( .A1(n28637), .A2(n591), .B1(ram[1994]), .B2(n592), .ZN(
        n6235) );
  MOAI22 U15165 ( .A1(n28402), .A2(n591), .B1(ram[1995]), .B2(n592), .ZN(
        n6236) );
  MOAI22 U15166 ( .A1(n28167), .A2(n591), .B1(ram[1996]), .B2(n592), .ZN(
        n6237) );
  MOAI22 U15167 ( .A1(n27932), .A2(n591), .B1(ram[1997]), .B2(n592), .ZN(
        n6238) );
  MOAI22 U15168 ( .A1(n27697), .A2(n591), .B1(ram[1998]), .B2(n592), .ZN(
        n6239) );
  MOAI22 U15169 ( .A1(n27462), .A2(n591), .B1(ram[1999]), .B2(n592), .ZN(
        n6240) );
  MOAI22 U15170 ( .A1(n29107), .A2(n593), .B1(ram[2000]), .B2(n594), .ZN(
        n6241) );
  MOAI22 U15171 ( .A1(n28872), .A2(n593), .B1(ram[2001]), .B2(n594), .ZN(
        n6242) );
  MOAI22 U15172 ( .A1(n28637), .A2(n593), .B1(ram[2002]), .B2(n594), .ZN(
        n6243) );
  MOAI22 U15173 ( .A1(n28402), .A2(n593), .B1(ram[2003]), .B2(n594), .ZN(
        n6244) );
  MOAI22 U15174 ( .A1(n28167), .A2(n593), .B1(ram[2004]), .B2(n594), .ZN(
        n6245) );
  MOAI22 U15175 ( .A1(n27932), .A2(n593), .B1(ram[2005]), .B2(n594), .ZN(
        n6246) );
  MOAI22 U15176 ( .A1(n27697), .A2(n593), .B1(ram[2006]), .B2(n594), .ZN(
        n6247) );
  MOAI22 U15177 ( .A1(n27462), .A2(n593), .B1(ram[2007]), .B2(n594), .ZN(
        n6248) );
  MOAI22 U15178 ( .A1(n29107), .A2(n595), .B1(ram[2008]), .B2(n596), .ZN(
        n6249) );
  MOAI22 U15179 ( .A1(n28872), .A2(n595), .B1(ram[2009]), .B2(n596), .ZN(
        n6250) );
  MOAI22 U15180 ( .A1(n28637), .A2(n595), .B1(ram[2010]), .B2(n596), .ZN(
        n6251) );
  MOAI22 U15181 ( .A1(n28402), .A2(n595), .B1(ram[2011]), .B2(n596), .ZN(
        n6252) );
  MOAI22 U15182 ( .A1(n28167), .A2(n595), .B1(ram[2012]), .B2(n596), .ZN(
        n6253) );
  MOAI22 U15183 ( .A1(n27932), .A2(n595), .B1(ram[2013]), .B2(n596), .ZN(
        n6254) );
  MOAI22 U15184 ( .A1(n27697), .A2(n595), .B1(ram[2014]), .B2(n596), .ZN(
        n6255) );
  MOAI22 U15185 ( .A1(n27462), .A2(n595), .B1(ram[2015]), .B2(n596), .ZN(
        n6256) );
  MOAI22 U15186 ( .A1(n29107), .A2(n597), .B1(ram[2016]), .B2(n598), .ZN(
        n6257) );
  MOAI22 U15187 ( .A1(n28872), .A2(n597), .B1(ram[2017]), .B2(n598), .ZN(
        n6258) );
  MOAI22 U15188 ( .A1(n28637), .A2(n597), .B1(ram[2018]), .B2(n598), .ZN(
        n6259) );
  MOAI22 U15189 ( .A1(n28402), .A2(n597), .B1(ram[2019]), .B2(n598), .ZN(
        n6260) );
  MOAI22 U15190 ( .A1(n28167), .A2(n597), .B1(ram[2020]), .B2(n598), .ZN(
        n6261) );
  MOAI22 U15191 ( .A1(n27932), .A2(n597), .B1(ram[2021]), .B2(n598), .ZN(
        n6262) );
  MOAI22 U15192 ( .A1(n27697), .A2(n597), .B1(ram[2022]), .B2(n598), .ZN(
        n6263) );
  MOAI22 U15193 ( .A1(n27462), .A2(n597), .B1(ram[2023]), .B2(n598), .ZN(
        n6264) );
  MOAI22 U15194 ( .A1(n29107), .A2(n599), .B1(ram[2024]), .B2(n600), .ZN(
        n6265) );
  MOAI22 U15195 ( .A1(n28872), .A2(n599), .B1(ram[2025]), .B2(n600), .ZN(
        n6266) );
  MOAI22 U15196 ( .A1(n28637), .A2(n599), .B1(ram[2026]), .B2(n600), .ZN(
        n6267) );
  MOAI22 U15197 ( .A1(n28402), .A2(n599), .B1(ram[2027]), .B2(n600), .ZN(
        n6268) );
  MOAI22 U15198 ( .A1(n28167), .A2(n599), .B1(ram[2028]), .B2(n600), .ZN(
        n6269) );
  MOAI22 U15199 ( .A1(n27932), .A2(n599), .B1(ram[2029]), .B2(n600), .ZN(
        n6270) );
  MOAI22 U15200 ( .A1(n27697), .A2(n599), .B1(ram[2030]), .B2(n600), .ZN(
        n6271) );
  MOAI22 U15201 ( .A1(n27462), .A2(n599), .B1(ram[2031]), .B2(n600), .ZN(
        n6272) );
  MOAI22 U15202 ( .A1(n29107), .A2(n601), .B1(ram[2032]), .B2(n602), .ZN(
        n6273) );
  MOAI22 U15203 ( .A1(n28872), .A2(n601), .B1(ram[2033]), .B2(n602), .ZN(
        n6274) );
  MOAI22 U15204 ( .A1(n28637), .A2(n601), .B1(ram[2034]), .B2(n602), .ZN(
        n6275) );
  MOAI22 U15205 ( .A1(n28402), .A2(n601), .B1(ram[2035]), .B2(n602), .ZN(
        n6276) );
  MOAI22 U15206 ( .A1(n28167), .A2(n601), .B1(ram[2036]), .B2(n602), .ZN(
        n6277) );
  MOAI22 U15207 ( .A1(n27932), .A2(n601), .B1(ram[2037]), .B2(n602), .ZN(
        n6278) );
  MOAI22 U15208 ( .A1(n27697), .A2(n601), .B1(ram[2038]), .B2(n602), .ZN(
        n6279) );
  MOAI22 U15209 ( .A1(n27462), .A2(n601), .B1(ram[2039]), .B2(n602), .ZN(
        n6280) );
  MOAI22 U15210 ( .A1(n29107), .A2(n603), .B1(ram[2040]), .B2(n604), .ZN(
        n6281) );
  MOAI22 U15211 ( .A1(n28872), .A2(n603), .B1(ram[2041]), .B2(n604), .ZN(
        n6282) );
  MOAI22 U15212 ( .A1(n28637), .A2(n603), .B1(ram[2042]), .B2(n604), .ZN(
        n6283) );
  MOAI22 U15213 ( .A1(n28402), .A2(n603), .B1(ram[2043]), .B2(n604), .ZN(
        n6284) );
  MOAI22 U15214 ( .A1(n28167), .A2(n603), .B1(ram[2044]), .B2(n604), .ZN(
        n6285) );
  MOAI22 U15215 ( .A1(n27932), .A2(n603), .B1(ram[2045]), .B2(n604), .ZN(
        n6286) );
  MOAI22 U15216 ( .A1(n27697), .A2(n603), .B1(ram[2046]), .B2(n604), .ZN(
        n6287) );
  MOAI22 U15217 ( .A1(n27462), .A2(n603), .B1(ram[2047]), .B2(n604), .ZN(
        n6288) );
  MOAI22 U15218 ( .A1(n29107), .A2(n606), .B1(ram[2048]), .B2(n607), .ZN(
        n6289) );
  MOAI22 U15219 ( .A1(n28872), .A2(n606), .B1(ram[2049]), .B2(n607), .ZN(
        n6290) );
  MOAI22 U15220 ( .A1(n28637), .A2(n606), .B1(ram[2050]), .B2(n607), .ZN(
        n6291) );
  MOAI22 U15221 ( .A1(n28402), .A2(n606), .B1(ram[2051]), .B2(n607), .ZN(
        n6292) );
  MOAI22 U15222 ( .A1(n28167), .A2(n606), .B1(ram[2052]), .B2(n607), .ZN(
        n6293) );
  MOAI22 U15223 ( .A1(n27932), .A2(n606), .B1(ram[2053]), .B2(n607), .ZN(
        n6294) );
  MOAI22 U15224 ( .A1(n27697), .A2(n606), .B1(ram[2054]), .B2(n607), .ZN(
        n6295) );
  MOAI22 U15225 ( .A1(n27462), .A2(n606), .B1(ram[2055]), .B2(n607), .ZN(
        n6296) );
  MOAI22 U15226 ( .A1(n29107), .A2(n609), .B1(ram[2056]), .B2(n610), .ZN(
        n6297) );
  MOAI22 U15227 ( .A1(n28872), .A2(n609), .B1(ram[2057]), .B2(n610), .ZN(
        n6298) );
  MOAI22 U15228 ( .A1(n28637), .A2(n609), .B1(ram[2058]), .B2(n610), .ZN(
        n6299) );
  MOAI22 U15229 ( .A1(n28402), .A2(n609), .B1(ram[2059]), .B2(n610), .ZN(
        n6300) );
  MOAI22 U15230 ( .A1(n28167), .A2(n609), .B1(ram[2060]), .B2(n610), .ZN(
        n6301) );
  MOAI22 U15231 ( .A1(n27932), .A2(n609), .B1(ram[2061]), .B2(n610), .ZN(
        n6302) );
  MOAI22 U15232 ( .A1(n27697), .A2(n609), .B1(ram[2062]), .B2(n610), .ZN(
        n6303) );
  MOAI22 U15233 ( .A1(n27462), .A2(n609), .B1(ram[2063]), .B2(n610), .ZN(
        n6304) );
  MOAI22 U15234 ( .A1(n29107), .A2(n611), .B1(ram[2064]), .B2(n612), .ZN(
        n6305) );
  MOAI22 U15235 ( .A1(n28872), .A2(n611), .B1(ram[2065]), .B2(n612), .ZN(
        n6306) );
  MOAI22 U15236 ( .A1(n28637), .A2(n611), .B1(ram[2066]), .B2(n612), .ZN(
        n6307) );
  MOAI22 U15237 ( .A1(n28402), .A2(n611), .B1(ram[2067]), .B2(n612), .ZN(
        n6308) );
  MOAI22 U15238 ( .A1(n28167), .A2(n611), .B1(ram[2068]), .B2(n612), .ZN(
        n6309) );
  MOAI22 U15239 ( .A1(n27932), .A2(n611), .B1(ram[2069]), .B2(n612), .ZN(
        n6310) );
  MOAI22 U15240 ( .A1(n27697), .A2(n611), .B1(ram[2070]), .B2(n612), .ZN(
        n6311) );
  MOAI22 U15241 ( .A1(n27462), .A2(n611), .B1(ram[2071]), .B2(n612), .ZN(
        n6312) );
  MOAI22 U15242 ( .A1(n29107), .A2(n613), .B1(ram[2072]), .B2(n614), .ZN(
        n6313) );
  MOAI22 U15243 ( .A1(n28872), .A2(n613), .B1(ram[2073]), .B2(n614), .ZN(
        n6314) );
  MOAI22 U15244 ( .A1(n28637), .A2(n613), .B1(ram[2074]), .B2(n614), .ZN(
        n6315) );
  MOAI22 U15245 ( .A1(n28402), .A2(n613), .B1(ram[2075]), .B2(n614), .ZN(
        n6316) );
  MOAI22 U15246 ( .A1(n28167), .A2(n613), .B1(ram[2076]), .B2(n614), .ZN(
        n6317) );
  MOAI22 U15247 ( .A1(n27932), .A2(n613), .B1(ram[2077]), .B2(n614), .ZN(
        n6318) );
  MOAI22 U15248 ( .A1(n27697), .A2(n613), .B1(ram[2078]), .B2(n614), .ZN(
        n6319) );
  MOAI22 U15249 ( .A1(n27462), .A2(n613), .B1(ram[2079]), .B2(n614), .ZN(
        n6320) );
  MOAI22 U15250 ( .A1(n29108), .A2(n615), .B1(ram[2080]), .B2(n616), .ZN(
        n6321) );
  MOAI22 U15251 ( .A1(n28873), .A2(n615), .B1(ram[2081]), .B2(n616), .ZN(
        n6322) );
  MOAI22 U15252 ( .A1(n28638), .A2(n615), .B1(ram[2082]), .B2(n616), .ZN(
        n6323) );
  MOAI22 U15253 ( .A1(n28403), .A2(n615), .B1(ram[2083]), .B2(n616), .ZN(
        n6324) );
  MOAI22 U15254 ( .A1(n28168), .A2(n615), .B1(ram[2084]), .B2(n616), .ZN(
        n6325) );
  MOAI22 U15255 ( .A1(n27933), .A2(n615), .B1(ram[2085]), .B2(n616), .ZN(
        n6326) );
  MOAI22 U15256 ( .A1(n27698), .A2(n615), .B1(ram[2086]), .B2(n616), .ZN(
        n6327) );
  MOAI22 U15257 ( .A1(n27463), .A2(n615), .B1(ram[2087]), .B2(n616), .ZN(
        n6328) );
  MOAI22 U15258 ( .A1(n29108), .A2(n617), .B1(ram[2088]), .B2(n618), .ZN(
        n6329) );
  MOAI22 U15259 ( .A1(n28873), .A2(n617), .B1(ram[2089]), .B2(n618), .ZN(
        n6330) );
  MOAI22 U15260 ( .A1(n28638), .A2(n617), .B1(ram[2090]), .B2(n618), .ZN(
        n6331) );
  MOAI22 U15261 ( .A1(n28403), .A2(n617), .B1(ram[2091]), .B2(n618), .ZN(
        n6332) );
  MOAI22 U15262 ( .A1(n28168), .A2(n617), .B1(ram[2092]), .B2(n618), .ZN(
        n6333) );
  MOAI22 U15263 ( .A1(n27933), .A2(n617), .B1(ram[2093]), .B2(n618), .ZN(
        n6334) );
  MOAI22 U15264 ( .A1(n27698), .A2(n617), .B1(ram[2094]), .B2(n618), .ZN(
        n6335) );
  MOAI22 U15265 ( .A1(n27463), .A2(n617), .B1(ram[2095]), .B2(n618), .ZN(
        n6336) );
  MOAI22 U15266 ( .A1(n29108), .A2(n619), .B1(ram[2096]), .B2(n620), .ZN(
        n6337) );
  MOAI22 U15267 ( .A1(n28873), .A2(n619), .B1(ram[2097]), .B2(n620), .ZN(
        n6338) );
  MOAI22 U15268 ( .A1(n28638), .A2(n619), .B1(ram[2098]), .B2(n620), .ZN(
        n6339) );
  MOAI22 U15269 ( .A1(n28403), .A2(n619), .B1(ram[2099]), .B2(n620), .ZN(
        n6340) );
  MOAI22 U15270 ( .A1(n28168), .A2(n619), .B1(ram[2100]), .B2(n620), .ZN(
        n6341) );
  MOAI22 U15271 ( .A1(n27933), .A2(n619), .B1(ram[2101]), .B2(n620), .ZN(
        n6342) );
  MOAI22 U15272 ( .A1(n27698), .A2(n619), .B1(ram[2102]), .B2(n620), .ZN(
        n6343) );
  MOAI22 U15273 ( .A1(n27463), .A2(n619), .B1(ram[2103]), .B2(n620), .ZN(
        n6344) );
  MOAI22 U15274 ( .A1(n29108), .A2(n621), .B1(ram[2104]), .B2(n622), .ZN(
        n6345) );
  MOAI22 U15275 ( .A1(n28873), .A2(n621), .B1(ram[2105]), .B2(n622), .ZN(
        n6346) );
  MOAI22 U15276 ( .A1(n28638), .A2(n621), .B1(ram[2106]), .B2(n622), .ZN(
        n6347) );
  MOAI22 U15277 ( .A1(n28403), .A2(n621), .B1(ram[2107]), .B2(n622), .ZN(
        n6348) );
  MOAI22 U15278 ( .A1(n28168), .A2(n621), .B1(ram[2108]), .B2(n622), .ZN(
        n6349) );
  MOAI22 U15279 ( .A1(n27933), .A2(n621), .B1(ram[2109]), .B2(n622), .ZN(
        n6350) );
  MOAI22 U15280 ( .A1(n27698), .A2(n621), .B1(ram[2110]), .B2(n622), .ZN(
        n6351) );
  MOAI22 U15281 ( .A1(n27463), .A2(n621), .B1(ram[2111]), .B2(n622), .ZN(
        n6352) );
  MOAI22 U15282 ( .A1(n29108), .A2(n623), .B1(ram[2112]), .B2(n624), .ZN(
        n6353) );
  MOAI22 U15283 ( .A1(n28873), .A2(n623), .B1(ram[2113]), .B2(n624), .ZN(
        n6354) );
  MOAI22 U15284 ( .A1(n28638), .A2(n623), .B1(ram[2114]), .B2(n624), .ZN(
        n6355) );
  MOAI22 U15285 ( .A1(n28403), .A2(n623), .B1(ram[2115]), .B2(n624), .ZN(
        n6356) );
  MOAI22 U15286 ( .A1(n28168), .A2(n623), .B1(ram[2116]), .B2(n624), .ZN(
        n6357) );
  MOAI22 U15287 ( .A1(n27933), .A2(n623), .B1(ram[2117]), .B2(n624), .ZN(
        n6358) );
  MOAI22 U15288 ( .A1(n27698), .A2(n623), .B1(ram[2118]), .B2(n624), .ZN(
        n6359) );
  MOAI22 U15289 ( .A1(n27463), .A2(n623), .B1(ram[2119]), .B2(n624), .ZN(
        n6360) );
  MOAI22 U15290 ( .A1(n29108), .A2(n625), .B1(ram[2120]), .B2(n626), .ZN(
        n6361) );
  MOAI22 U15291 ( .A1(n28873), .A2(n625), .B1(ram[2121]), .B2(n626), .ZN(
        n6362) );
  MOAI22 U15292 ( .A1(n28638), .A2(n625), .B1(ram[2122]), .B2(n626), .ZN(
        n6363) );
  MOAI22 U15293 ( .A1(n28403), .A2(n625), .B1(ram[2123]), .B2(n626), .ZN(
        n6364) );
  MOAI22 U15294 ( .A1(n28168), .A2(n625), .B1(ram[2124]), .B2(n626), .ZN(
        n6365) );
  MOAI22 U15295 ( .A1(n27933), .A2(n625), .B1(ram[2125]), .B2(n626), .ZN(
        n6366) );
  MOAI22 U15296 ( .A1(n27698), .A2(n625), .B1(ram[2126]), .B2(n626), .ZN(
        n6367) );
  MOAI22 U15297 ( .A1(n27463), .A2(n625), .B1(ram[2127]), .B2(n626), .ZN(
        n6368) );
  MOAI22 U15298 ( .A1(n29108), .A2(n627), .B1(ram[2128]), .B2(n628), .ZN(
        n6369) );
  MOAI22 U15299 ( .A1(n28873), .A2(n627), .B1(ram[2129]), .B2(n628), .ZN(
        n6370) );
  MOAI22 U15300 ( .A1(n28638), .A2(n627), .B1(ram[2130]), .B2(n628), .ZN(
        n6371) );
  MOAI22 U15301 ( .A1(n28403), .A2(n627), .B1(ram[2131]), .B2(n628), .ZN(
        n6372) );
  MOAI22 U15302 ( .A1(n28168), .A2(n627), .B1(ram[2132]), .B2(n628), .ZN(
        n6373) );
  MOAI22 U15303 ( .A1(n27933), .A2(n627), .B1(ram[2133]), .B2(n628), .ZN(
        n6374) );
  MOAI22 U15304 ( .A1(n27698), .A2(n627), .B1(ram[2134]), .B2(n628), .ZN(
        n6375) );
  MOAI22 U15305 ( .A1(n27463), .A2(n627), .B1(ram[2135]), .B2(n628), .ZN(
        n6376) );
  MOAI22 U15306 ( .A1(n29108), .A2(n629), .B1(ram[2136]), .B2(n630), .ZN(
        n6377) );
  MOAI22 U15307 ( .A1(n28873), .A2(n629), .B1(ram[2137]), .B2(n630), .ZN(
        n6378) );
  MOAI22 U15308 ( .A1(n28638), .A2(n629), .B1(ram[2138]), .B2(n630), .ZN(
        n6379) );
  MOAI22 U15309 ( .A1(n28403), .A2(n629), .B1(ram[2139]), .B2(n630), .ZN(
        n6380) );
  MOAI22 U15310 ( .A1(n28168), .A2(n629), .B1(ram[2140]), .B2(n630), .ZN(
        n6381) );
  MOAI22 U15311 ( .A1(n27933), .A2(n629), .B1(ram[2141]), .B2(n630), .ZN(
        n6382) );
  MOAI22 U15312 ( .A1(n27698), .A2(n629), .B1(ram[2142]), .B2(n630), .ZN(
        n6383) );
  MOAI22 U15313 ( .A1(n27463), .A2(n629), .B1(ram[2143]), .B2(n630), .ZN(
        n6384) );
  MOAI22 U15314 ( .A1(n29108), .A2(n631), .B1(ram[2144]), .B2(n632), .ZN(
        n6385) );
  MOAI22 U15315 ( .A1(n28873), .A2(n631), .B1(ram[2145]), .B2(n632), .ZN(
        n6386) );
  MOAI22 U15316 ( .A1(n28638), .A2(n631), .B1(ram[2146]), .B2(n632), .ZN(
        n6387) );
  MOAI22 U15317 ( .A1(n28403), .A2(n631), .B1(ram[2147]), .B2(n632), .ZN(
        n6388) );
  MOAI22 U15318 ( .A1(n28168), .A2(n631), .B1(ram[2148]), .B2(n632), .ZN(
        n6389) );
  MOAI22 U15319 ( .A1(n27933), .A2(n631), .B1(ram[2149]), .B2(n632), .ZN(
        n6390) );
  MOAI22 U15320 ( .A1(n27698), .A2(n631), .B1(ram[2150]), .B2(n632), .ZN(
        n6391) );
  MOAI22 U15321 ( .A1(n27463), .A2(n631), .B1(ram[2151]), .B2(n632), .ZN(
        n6392) );
  MOAI22 U15322 ( .A1(n29108), .A2(n633), .B1(ram[2152]), .B2(n634), .ZN(
        n6393) );
  MOAI22 U15323 ( .A1(n28873), .A2(n633), .B1(ram[2153]), .B2(n634), .ZN(
        n6394) );
  MOAI22 U15324 ( .A1(n28638), .A2(n633), .B1(ram[2154]), .B2(n634), .ZN(
        n6395) );
  MOAI22 U15325 ( .A1(n28403), .A2(n633), .B1(ram[2155]), .B2(n634), .ZN(
        n6396) );
  MOAI22 U15326 ( .A1(n28168), .A2(n633), .B1(ram[2156]), .B2(n634), .ZN(
        n6397) );
  MOAI22 U15327 ( .A1(n27933), .A2(n633), .B1(ram[2157]), .B2(n634), .ZN(
        n6398) );
  MOAI22 U15328 ( .A1(n27698), .A2(n633), .B1(ram[2158]), .B2(n634), .ZN(
        n6399) );
  MOAI22 U15329 ( .A1(n27463), .A2(n633), .B1(ram[2159]), .B2(n634), .ZN(
        n6400) );
  MOAI22 U15330 ( .A1(n29108), .A2(n635), .B1(ram[2160]), .B2(n636), .ZN(
        n6401) );
  MOAI22 U15331 ( .A1(n28873), .A2(n635), .B1(ram[2161]), .B2(n636), .ZN(
        n6402) );
  MOAI22 U15332 ( .A1(n28638), .A2(n635), .B1(ram[2162]), .B2(n636), .ZN(
        n6403) );
  MOAI22 U15333 ( .A1(n28403), .A2(n635), .B1(ram[2163]), .B2(n636), .ZN(
        n6404) );
  MOAI22 U15334 ( .A1(n28168), .A2(n635), .B1(ram[2164]), .B2(n636), .ZN(
        n6405) );
  MOAI22 U15335 ( .A1(n27933), .A2(n635), .B1(ram[2165]), .B2(n636), .ZN(
        n6406) );
  MOAI22 U15336 ( .A1(n27698), .A2(n635), .B1(ram[2166]), .B2(n636), .ZN(
        n6407) );
  MOAI22 U15337 ( .A1(n27463), .A2(n635), .B1(ram[2167]), .B2(n636), .ZN(
        n6408) );
  MOAI22 U15338 ( .A1(n29108), .A2(n637), .B1(ram[2168]), .B2(n638), .ZN(
        n6409) );
  MOAI22 U15339 ( .A1(n28873), .A2(n637), .B1(ram[2169]), .B2(n638), .ZN(
        n6410) );
  MOAI22 U15340 ( .A1(n28638), .A2(n637), .B1(ram[2170]), .B2(n638), .ZN(
        n6411) );
  MOAI22 U15341 ( .A1(n28403), .A2(n637), .B1(ram[2171]), .B2(n638), .ZN(
        n6412) );
  MOAI22 U15342 ( .A1(n28168), .A2(n637), .B1(ram[2172]), .B2(n638), .ZN(
        n6413) );
  MOAI22 U15343 ( .A1(n27933), .A2(n637), .B1(ram[2173]), .B2(n638), .ZN(
        n6414) );
  MOAI22 U15344 ( .A1(n27698), .A2(n637), .B1(ram[2174]), .B2(n638), .ZN(
        n6415) );
  MOAI22 U15345 ( .A1(n27463), .A2(n637), .B1(ram[2175]), .B2(n638), .ZN(
        n6416) );
  MOAI22 U15346 ( .A1(n29108), .A2(n639), .B1(ram[2176]), .B2(n640), .ZN(
        n6417) );
  MOAI22 U15347 ( .A1(n28873), .A2(n639), .B1(ram[2177]), .B2(n640), .ZN(
        n6418) );
  MOAI22 U15348 ( .A1(n28638), .A2(n639), .B1(ram[2178]), .B2(n640), .ZN(
        n6419) );
  MOAI22 U15349 ( .A1(n28403), .A2(n639), .B1(ram[2179]), .B2(n640), .ZN(
        n6420) );
  MOAI22 U15350 ( .A1(n28168), .A2(n639), .B1(ram[2180]), .B2(n640), .ZN(
        n6421) );
  MOAI22 U15351 ( .A1(n27933), .A2(n639), .B1(ram[2181]), .B2(n640), .ZN(
        n6422) );
  MOAI22 U15352 ( .A1(n27698), .A2(n639), .B1(ram[2182]), .B2(n640), .ZN(
        n6423) );
  MOAI22 U15353 ( .A1(n27463), .A2(n639), .B1(ram[2183]), .B2(n640), .ZN(
        n6424) );
  MOAI22 U15354 ( .A1(n29109), .A2(n641), .B1(ram[2184]), .B2(n642), .ZN(
        n6425) );
  MOAI22 U15355 ( .A1(n28874), .A2(n641), .B1(ram[2185]), .B2(n642), .ZN(
        n6426) );
  MOAI22 U15356 ( .A1(n28639), .A2(n641), .B1(ram[2186]), .B2(n642), .ZN(
        n6427) );
  MOAI22 U15357 ( .A1(n28404), .A2(n641), .B1(ram[2187]), .B2(n642), .ZN(
        n6428) );
  MOAI22 U15358 ( .A1(n28169), .A2(n641), .B1(ram[2188]), .B2(n642), .ZN(
        n6429) );
  MOAI22 U15359 ( .A1(n27934), .A2(n641), .B1(ram[2189]), .B2(n642), .ZN(
        n6430) );
  MOAI22 U15360 ( .A1(n27699), .A2(n641), .B1(ram[2190]), .B2(n642), .ZN(
        n6431) );
  MOAI22 U15361 ( .A1(n27464), .A2(n641), .B1(ram[2191]), .B2(n642), .ZN(
        n6432) );
  MOAI22 U15362 ( .A1(n29109), .A2(n643), .B1(ram[2192]), .B2(n644), .ZN(
        n6433) );
  MOAI22 U15363 ( .A1(n28874), .A2(n643), .B1(ram[2193]), .B2(n644), .ZN(
        n6434) );
  MOAI22 U15364 ( .A1(n28639), .A2(n643), .B1(ram[2194]), .B2(n644), .ZN(
        n6435) );
  MOAI22 U15365 ( .A1(n28404), .A2(n643), .B1(ram[2195]), .B2(n644), .ZN(
        n6436) );
  MOAI22 U15366 ( .A1(n28169), .A2(n643), .B1(ram[2196]), .B2(n644), .ZN(
        n6437) );
  MOAI22 U15367 ( .A1(n27934), .A2(n643), .B1(ram[2197]), .B2(n644), .ZN(
        n6438) );
  MOAI22 U15368 ( .A1(n27699), .A2(n643), .B1(ram[2198]), .B2(n644), .ZN(
        n6439) );
  MOAI22 U15369 ( .A1(n27464), .A2(n643), .B1(ram[2199]), .B2(n644), .ZN(
        n6440) );
  MOAI22 U15370 ( .A1(n29109), .A2(n645), .B1(ram[2200]), .B2(n646), .ZN(
        n6441) );
  MOAI22 U15371 ( .A1(n28874), .A2(n645), .B1(ram[2201]), .B2(n646), .ZN(
        n6442) );
  MOAI22 U15372 ( .A1(n28639), .A2(n645), .B1(ram[2202]), .B2(n646), .ZN(
        n6443) );
  MOAI22 U15373 ( .A1(n28404), .A2(n645), .B1(ram[2203]), .B2(n646), .ZN(
        n6444) );
  MOAI22 U15374 ( .A1(n28169), .A2(n645), .B1(ram[2204]), .B2(n646), .ZN(
        n6445) );
  MOAI22 U15375 ( .A1(n27934), .A2(n645), .B1(ram[2205]), .B2(n646), .ZN(
        n6446) );
  MOAI22 U15376 ( .A1(n27699), .A2(n645), .B1(ram[2206]), .B2(n646), .ZN(
        n6447) );
  MOAI22 U15377 ( .A1(n27464), .A2(n645), .B1(ram[2207]), .B2(n646), .ZN(
        n6448) );
  MOAI22 U15378 ( .A1(n29109), .A2(n647), .B1(ram[2208]), .B2(n648), .ZN(
        n6449) );
  MOAI22 U15379 ( .A1(n28874), .A2(n647), .B1(ram[2209]), .B2(n648), .ZN(
        n6450) );
  MOAI22 U15380 ( .A1(n28639), .A2(n647), .B1(ram[2210]), .B2(n648), .ZN(
        n6451) );
  MOAI22 U15381 ( .A1(n28404), .A2(n647), .B1(ram[2211]), .B2(n648), .ZN(
        n6452) );
  MOAI22 U15382 ( .A1(n28169), .A2(n647), .B1(ram[2212]), .B2(n648), .ZN(
        n6453) );
  MOAI22 U15383 ( .A1(n27934), .A2(n647), .B1(ram[2213]), .B2(n648), .ZN(
        n6454) );
  MOAI22 U15384 ( .A1(n27699), .A2(n647), .B1(ram[2214]), .B2(n648), .ZN(
        n6455) );
  MOAI22 U15385 ( .A1(n27464), .A2(n647), .B1(ram[2215]), .B2(n648), .ZN(
        n6456) );
  MOAI22 U15386 ( .A1(n29109), .A2(n649), .B1(ram[2216]), .B2(n650), .ZN(
        n6457) );
  MOAI22 U15387 ( .A1(n28874), .A2(n649), .B1(ram[2217]), .B2(n650), .ZN(
        n6458) );
  MOAI22 U15388 ( .A1(n28639), .A2(n649), .B1(ram[2218]), .B2(n650), .ZN(
        n6459) );
  MOAI22 U15389 ( .A1(n28404), .A2(n649), .B1(ram[2219]), .B2(n650), .ZN(
        n6460) );
  MOAI22 U15390 ( .A1(n28169), .A2(n649), .B1(ram[2220]), .B2(n650), .ZN(
        n6461) );
  MOAI22 U15391 ( .A1(n27934), .A2(n649), .B1(ram[2221]), .B2(n650), .ZN(
        n6462) );
  MOAI22 U15392 ( .A1(n27699), .A2(n649), .B1(ram[2222]), .B2(n650), .ZN(
        n6463) );
  MOAI22 U15393 ( .A1(n27464), .A2(n649), .B1(ram[2223]), .B2(n650), .ZN(
        n6464) );
  MOAI22 U15394 ( .A1(n29109), .A2(n651), .B1(ram[2224]), .B2(n652), .ZN(
        n6465) );
  MOAI22 U15395 ( .A1(n28874), .A2(n651), .B1(ram[2225]), .B2(n652), .ZN(
        n6466) );
  MOAI22 U15396 ( .A1(n28639), .A2(n651), .B1(ram[2226]), .B2(n652), .ZN(
        n6467) );
  MOAI22 U15397 ( .A1(n28404), .A2(n651), .B1(ram[2227]), .B2(n652), .ZN(
        n6468) );
  MOAI22 U15398 ( .A1(n28169), .A2(n651), .B1(ram[2228]), .B2(n652), .ZN(
        n6469) );
  MOAI22 U15399 ( .A1(n27934), .A2(n651), .B1(ram[2229]), .B2(n652), .ZN(
        n6470) );
  MOAI22 U15400 ( .A1(n27699), .A2(n651), .B1(ram[2230]), .B2(n652), .ZN(
        n6471) );
  MOAI22 U15401 ( .A1(n27464), .A2(n651), .B1(ram[2231]), .B2(n652), .ZN(
        n6472) );
  MOAI22 U15402 ( .A1(n29109), .A2(n653), .B1(ram[2232]), .B2(n654), .ZN(
        n6473) );
  MOAI22 U15403 ( .A1(n28874), .A2(n653), .B1(ram[2233]), .B2(n654), .ZN(
        n6474) );
  MOAI22 U15404 ( .A1(n28639), .A2(n653), .B1(ram[2234]), .B2(n654), .ZN(
        n6475) );
  MOAI22 U15405 ( .A1(n28404), .A2(n653), .B1(ram[2235]), .B2(n654), .ZN(
        n6476) );
  MOAI22 U15406 ( .A1(n28169), .A2(n653), .B1(ram[2236]), .B2(n654), .ZN(
        n6477) );
  MOAI22 U15407 ( .A1(n27934), .A2(n653), .B1(ram[2237]), .B2(n654), .ZN(
        n6478) );
  MOAI22 U15408 ( .A1(n27699), .A2(n653), .B1(ram[2238]), .B2(n654), .ZN(
        n6479) );
  MOAI22 U15409 ( .A1(n27464), .A2(n653), .B1(ram[2239]), .B2(n654), .ZN(
        n6480) );
  MOAI22 U15410 ( .A1(n29109), .A2(n655), .B1(ram[2240]), .B2(n656), .ZN(
        n6481) );
  MOAI22 U15411 ( .A1(n28874), .A2(n655), .B1(ram[2241]), .B2(n656), .ZN(
        n6482) );
  MOAI22 U15412 ( .A1(n28639), .A2(n655), .B1(ram[2242]), .B2(n656), .ZN(
        n6483) );
  MOAI22 U15413 ( .A1(n28404), .A2(n655), .B1(ram[2243]), .B2(n656), .ZN(
        n6484) );
  MOAI22 U15414 ( .A1(n28169), .A2(n655), .B1(ram[2244]), .B2(n656), .ZN(
        n6485) );
  MOAI22 U15415 ( .A1(n27934), .A2(n655), .B1(ram[2245]), .B2(n656), .ZN(
        n6486) );
  MOAI22 U15416 ( .A1(n27699), .A2(n655), .B1(ram[2246]), .B2(n656), .ZN(
        n6487) );
  MOAI22 U15417 ( .A1(n27464), .A2(n655), .B1(ram[2247]), .B2(n656), .ZN(
        n6488) );
  MOAI22 U15418 ( .A1(n29109), .A2(n657), .B1(ram[2248]), .B2(n658), .ZN(
        n6489) );
  MOAI22 U15419 ( .A1(n28874), .A2(n657), .B1(ram[2249]), .B2(n658), .ZN(
        n6490) );
  MOAI22 U15420 ( .A1(n28639), .A2(n657), .B1(ram[2250]), .B2(n658), .ZN(
        n6491) );
  MOAI22 U15421 ( .A1(n28404), .A2(n657), .B1(ram[2251]), .B2(n658), .ZN(
        n6492) );
  MOAI22 U15422 ( .A1(n28169), .A2(n657), .B1(ram[2252]), .B2(n658), .ZN(
        n6493) );
  MOAI22 U15423 ( .A1(n27934), .A2(n657), .B1(ram[2253]), .B2(n658), .ZN(
        n6494) );
  MOAI22 U15424 ( .A1(n27699), .A2(n657), .B1(ram[2254]), .B2(n658), .ZN(
        n6495) );
  MOAI22 U15425 ( .A1(n27464), .A2(n657), .B1(ram[2255]), .B2(n658), .ZN(
        n6496) );
  MOAI22 U15426 ( .A1(n29109), .A2(n659), .B1(ram[2256]), .B2(n660), .ZN(
        n6497) );
  MOAI22 U15427 ( .A1(n28874), .A2(n659), .B1(ram[2257]), .B2(n660), .ZN(
        n6498) );
  MOAI22 U15428 ( .A1(n28639), .A2(n659), .B1(ram[2258]), .B2(n660), .ZN(
        n6499) );
  MOAI22 U15429 ( .A1(n28404), .A2(n659), .B1(ram[2259]), .B2(n660), .ZN(
        n6500) );
  MOAI22 U15430 ( .A1(n28169), .A2(n659), .B1(ram[2260]), .B2(n660), .ZN(
        n6501) );
  MOAI22 U15431 ( .A1(n27934), .A2(n659), .B1(ram[2261]), .B2(n660), .ZN(
        n6502) );
  MOAI22 U15432 ( .A1(n27699), .A2(n659), .B1(ram[2262]), .B2(n660), .ZN(
        n6503) );
  MOAI22 U15433 ( .A1(n27464), .A2(n659), .B1(ram[2263]), .B2(n660), .ZN(
        n6504) );
  MOAI22 U15434 ( .A1(n29109), .A2(n661), .B1(ram[2264]), .B2(n662), .ZN(
        n6505) );
  MOAI22 U15435 ( .A1(n28874), .A2(n661), .B1(ram[2265]), .B2(n662), .ZN(
        n6506) );
  MOAI22 U15436 ( .A1(n28639), .A2(n661), .B1(ram[2266]), .B2(n662), .ZN(
        n6507) );
  MOAI22 U15437 ( .A1(n28404), .A2(n661), .B1(ram[2267]), .B2(n662), .ZN(
        n6508) );
  MOAI22 U15438 ( .A1(n28169), .A2(n661), .B1(ram[2268]), .B2(n662), .ZN(
        n6509) );
  MOAI22 U15439 ( .A1(n27934), .A2(n661), .B1(ram[2269]), .B2(n662), .ZN(
        n6510) );
  MOAI22 U15440 ( .A1(n27699), .A2(n661), .B1(ram[2270]), .B2(n662), .ZN(
        n6511) );
  MOAI22 U15441 ( .A1(n27464), .A2(n661), .B1(ram[2271]), .B2(n662), .ZN(
        n6512) );
  MOAI22 U15442 ( .A1(n29109), .A2(n663), .B1(ram[2272]), .B2(n664), .ZN(
        n6513) );
  MOAI22 U15443 ( .A1(n28874), .A2(n663), .B1(ram[2273]), .B2(n664), .ZN(
        n6514) );
  MOAI22 U15444 ( .A1(n28639), .A2(n663), .B1(ram[2274]), .B2(n664), .ZN(
        n6515) );
  MOAI22 U15445 ( .A1(n28404), .A2(n663), .B1(ram[2275]), .B2(n664), .ZN(
        n6516) );
  MOAI22 U15446 ( .A1(n28169), .A2(n663), .B1(ram[2276]), .B2(n664), .ZN(
        n6517) );
  MOAI22 U15447 ( .A1(n27934), .A2(n663), .B1(ram[2277]), .B2(n664), .ZN(
        n6518) );
  MOAI22 U15448 ( .A1(n27699), .A2(n663), .B1(ram[2278]), .B2(n664), .ZN(
        n6519) );
  MOAI22 U15449 ( .A1(n27464), .A2(n663), .B1(ram[2279]), .B2(n664), .ZN(
        n6520) );
  MOAI22 U15450 ( .A1(n29109), .A2(n665), .B1(ram[2280]), .B2(n666), .ZN(
        n6521) );
  MOAI22 U15451 ( .A1(n28874), .A2(n665), .B1(ram[2281]), .B2(n666), .ZN(
        n6522) );
  MOAI22 U15452 ( .A1(n28639), .A2(n665), .B1(ram[2282]), .B2(n666), .ZN(
        n6523) );
  MOAI22 U15453 ( .A1(n28404), .A2(n665), .B1(ram[2283]), .B2(n666), .ZN(
        n6524) );
  MOAI22 U15454 ( .A1(n28169), .A2(n665), .B1(ram[2284]), .B2(n666), .ZN(
        n6525) );
  MOAI22 U15455 ( .A1(n27934), .A2(n665), .B1(ram[2285]), .B2(n666), .ZN(
        n6526) );
  MOAI22 U15456 ( .A1(n27699), .A2(n665), .B1(ram[2286]), .B2(n666), .ZN(
        n6527) );
  MOAI22 U15457 ( .A1(n27464), .A2(n665), .B1(ram[2287]), .B2(n666), .ZN(
        n6528) );
  MOAI22 U15458 ( .A1(n29110), .A2(n667), .B1(ram[2288]), .B2(n668), .ZN(
        n6529) );
  MOAI22 U15459 ( .A1(n28875), .A2(n667), .B1(ram[2289]), .B2(n668), .ZN(
        n6530) );
  MOAI22 U15460 ( .A1(n28640), .A2(n667), .B1(ram[2290]), .B2(n668), .ZN(
        n6531) );
  MOAI22 U15461 ( .A1(n28405), .A2(n667), .B1(ram[2291]), .B2(n668), .ZN(
        n6532) );
  MOAI22 U15462 ( .A1(n28170), .A2(n667), .B1(ram[2292]), .B2(n668), .ZN(
        n6533) );
  MOAI22 U15463 ( .A1(n27935), .A2(n667), .B1(ram[2293]), .B2(n668), .ZN(
        n6534) );
  MOAI22 U15464 ( .A1(n27700), .A2(n667), .B1(ram[2294]), .B2(n668), .ZN(
        n6535) );
  MOAI22 U15465 ( .A1(n27465), .A2(n667), .B1(ram[2295]), .B2(n668), .ZN(
        n6536) );
  MOAI22 U15466 ( .A1(n29110), .A2(n669), .B1(ram[2296]), .B2(n670), .ZN(
        n6537) );
  MOAI22 U15467 ( .A1(n28875), .A2(n669), .B1(ram[2297]), .B2(n670), .ZN(
        n6538) );
  MOAI22 U15468 ( .A1(n28640), .A2(n669), .B1(ram[2298]), .B2(n670), .ZN(
        n6539) );
  MOAI22 U15469 ( .A1(n28405), .A2(n669), .B1(ram[2299]), .B2(n670), .ZN(
        n6540) );
  MOAI22 U15470 ( .A1(n28170), .A2(n669), .B1(ram[2300]), .B2(n670), .ZN(
        n6541) );
  MOAI22 U15471 ( .A1(n27935), .A2(n669), .B1(ram[2301]), .B2(n670), .ZN(
        n6542) );
  MOAI22 U15472 ( .A1(n27700), .A2(n669), .B1(ram[2302]), .B2(n670), .ZN(
        n6543) );
  MOAI22 U15473 ( .A1(n27465), .A2(n669), .B1(ram[2303]), .B2(n670), .ZN(
        n6544) );
  MOAI22 U15474 ( .A1(n29110), .A2(n671), .B1(ram[2304]), .B2(n672), .ZN(
        n6545) );
  MOAI22 U15475 ( .A1(n28875), .A2(n671), .B1(ram[2305]), .B2(n672), .ZN(
        n6546) );
  MOAI22 U15476 ( .A1(n28640), .A2(n671), .B1(ram[2306]), .B2(n672), .ZN(
        n6547) );
  MOAI22 U15477 ( .A1(n28405), .A2(n671), .B1(ram[2307]), .B2(n672), .ZN(
        n6548) );
  MOAI22 U15478 ( .A1(n28170), .A2(n671), .B1(ram[2308]), .B2(n672), .ZN(
        n6549) );
  MOAI22 U15479 ( .A1(n27935), .A2(n671), .B1(ram[2309]), .B2(n672), .ZN(
        n6550) );
  MOAI22 U15480 ( .A1(n27700), .A2(n671), .B1(ram[2310]), .B2(n672), .ZN(
        n6551) );
  MOAI22 U15481 ( .A1(n27465), .A2(n671), .B1(ram[2311]), .B2(n672), .ZN(
        n6552) );
  MOAI22 U15482 ( .A1(n29110), .A2(n673), .B1(ram[2312]), .B2(n674), .ZN(
        n6553) );
  MOAI22 U15483 ( .A1(n28875), .A2(n673), .B1(ram[2313]), .B2(n674), .ZN(
        n6554) );
  MOAI22 U15484 ( .A1(n28640), .A2(n673), .B1(ram[2314]), .B2(n674), .ZN(
        n6555) );
  MOAI22 U15485 ( .A1(n28405), .A2(n673), .B1(ram[2315]), .B2(n674), .ZN(
        n6556) );
  MOAI22 U15486 ( .A1(n28170), .A2(n673), .B1(ram[2316]), .B2(n674), .ZN(
        n6557) );
  MOAI22 U15487 ( .A1(n27935), .A2(n673), .B1(ram[2317]), .B2(n674), .ZN(
        n6558) );
  MOAI22 U15488 ( .A1(n27700), .A2(n673), .B1(ram[2318]), .B2(n674), .ZN(
        n6559) );
  MOAI22 U15489 ( .A1(n27465), .A2(n673), .B1(ram[2319]), .B2(n674), .ZN(
        n6560) );
  MOAI22 U15490 ( .A1(n29110), .A2(n675), .B1(ram[2320]), .B2(n676), .ZN(
        n6561) );
  MOAI22 U15491 ( .A1(n28875), .A2(n675), .B1(ram[2321]), .B2(n676), .ZN(
        n6562) );
  MOAI22 U15492 ( .A1(n28640), .A2(n675), .B1(ram[2322]), .B2(n676), .ZN(
        n6563) );
  MOAI22 U15493 ( .A1(n28405), .A2(n675), .B1(ram[2323]), .B2(n676), .ZN(
        n6564) );
  MOAI22 U15494 ( .A1(n28170), .A2(n675), .B1(ram[2324]), .B2(n676), .ZN(
        n6565) );
  MOAI22 U15495 ( .A1(n27935), .A2(n675), .B1(ram[2325]), .B2(n676), .ZN(
        n6566) );
  MOAI22 U15496 ( .A1(n27700), .A2(n675), .B1(ram[2326]), .B2(n676), .ZN(
        n6567) );
  MOAI22 U15497 ( .A1(n27465), .A2(n675), .B1(ram[2327]), .B2(n676), .ZN(
        n6568) );
  MOAI22 U15498 ( .A1(n29110), .A2(n677), .B1(ram[2328]), .B2(n678), .ZN(
        n6569) );
  MOAI22 U15499 ( .A1(n28875), .A2(n677), .B1(ram[2329]), .B2(n678), .ZN(
        n6570) );
  MOAI22 U15500 ( .A1(n28640), .A2(n677), .B1(ram[2330]), .B2(n678), .ZN(
        n6571) );
  MOAI22 U15501 ( .A1(n28405), .A2(n677), .B1(ram[2331]), .B2(n678), .ZN(
        n6572) );
  MOAI22 U15502 ( .A1(n28170), .A2(n677), .B1(ram[2332]), .B2(n678), .ZN(
        n6573) );
  MOAI22 U15503 ( .A1(n27935), .A2(n677), .B1(ram[2333]), .B2(n678), .ZN(
        n6574) );
  MOAI22 U15504 ( .A1(n27700), .A2(n677), .B1(ram[2334]), .B2(n678), .ZN(
        n6575) );
  MOAI22 U15505 ( .A1(n27465), .A2(n677), .B1(ram[2335]), .B2(n678), .ZN(
        n6576) );
  MOAI22 U15506 ( .A1(n29110), .A2(n679), .B1(ram[2336]), .B2(n680), .ZN(
        n6577) );
  MOAI22 U15507 ( .A1(n28875), .A2(n679), .B1(ram[2337]), .B2(n680), .ZN(
        n6578) );
  MOAI22 U15508 ( .A1(n28640), .A2(n679), .B1(ram[2338]), .B2(n680), .ZN(
        n6579) );
  MOAI22 U15509 ( .A1(n28405), .A2(n679), .B1(ram[2339]), .B2(n680), .ZN(
        n6580) );
  MOAI22 U15510 ( .A1(n28170), .A2(n679), .B1(ram[2340]), .B2(n680), .ZN(
        n6581) );
  MOAI22 U15511 ( .A1(n27935), .A2(n679), .B1(ram[2341]), .B2(n680), .ZN(
        n6582) );
  MOAI22 U15512 ( .A1(n27700), .A2(n679), .B1(ram[2342]), .B2(n680), .ZN(
        n6583) );
  MOAI22 U15513 ( .A1(n27465), .A2(n679), .B1(ram[2343]), .B2(n680), .ZN(
        n6584) );
  MOAI22 U15514 ( .A1(n29110), .A2(n681), .B1(ram[2344]), .B2(n682), .ZN(
        n6585) );
  MOAI22 U15515 ( .A1(n28875), .A2(n681), .B1(ram[2345]), .B2(n682), .ZN(
        n6586) );
  MOAI22 U15516 ( .A1(n28640), .A2(n681), .B1(ram[2346]), .B2(n682), .ZN(
        n6587) );
  MOAI22 U15517 ( .A1(n28405), .A2(n681), .B1(ram[2347]), .B2(n682), .ZN(
        n6588) );
  MOAI22 U15518 ( .A1(n28170), .A2(n681), .B1(ram[2348]), .B2(n682), .ZN(
        n6589) );
  MOAI22 U15519 ( .A1(n27935), .A2(n681), .B1(ram[2349]), .B2(n682), .ZN(
        n6590) );
  MOAI22 U15520 ( .A1(n27700), .A2(n681), .B1(ram[2350]), .B2(n682), .ZN(
        n6591) );
  MOAI22 U15521 ( .A1(n27465), .A2(n681), .B1(ram[2351]), .B2(n682), .ZN(
        n6592) );
  MOAI22 U15522 ( .A1(n29110), .A2(n683), .B1(ram[2352]), .B2(n684), .ZN(
        n6593) );
  MOAI22 U15523 ( .A1(n28875), .A2(n683), .B1(ram[2353]), .B2(n684), .ZN(
        n6594) );
  MOAI22 U15524 ( .A1(n28640), .A2(n683), .B1(ram[2354]), .B2(n684), .ZN(
        n6595) );
  MOAI22 U15525 ( .A1(n28405), .A2(n683), .B1(ram[2355]), .B2(n684), .ZN(
        n6596) );
  MOAI22 U15526 ( .A1(n28170), .A2(n683), .B1(ram[2356]), .B2(n684), .ZN(
        n6597) );
  MOAI22 U15527 ( .A1(n27935), .A2(n683), .B1(ram[2357]), .B2(n684), .ZN(
        n6598) );
  MOAI22 U15528 ( .A1(n27700), .A2(n683), .B1(ram[2358]), .B2(n684), .ZN(
        n6599) );
  MOAI22 U15529 ( .A1(n27465), .A2(n683), .B1(ram[2359]), .B2(n684), .ZN(
        n6600) );
  MOAI22 U15530 ( .A1(n29110), .A2(n685), .B1(ram[2360]), .B2(n686), .ZN(
        n6601) );
  MOAI22 U15531 ( .A1(n28875), .A2(n685), .B1(ram[2361]), .B2(n686), .ZN(
        n6602) );
  MOAI22 U15532 ( .A1(n28640), .A2(n685), .B1(ram[2362]), .B2(n686), .ZN(
        n6603) );
  MOAI22 U15533 ( .A1(n28405), .A2(n685), .B1(ram[2363]), .B2(n686), .ZN(
        n6604) );
  MOAI22 U15534 ( .A1(n28170), .A2(n685), .B1(ram[2364]), .B2(n686), .ZN(
        n6605) );
  MOAI22 U15535 ( .A1(n27935), .A2(n685), .B1(ram[2365]), .B2(n686), .ZN(
        n6606) );
  MOAI22 U15536 ( .A1(n27700), .A2(n685), .B1(ram[2366]), .B2(n686), .ZN(
        n6607) );
  MOAI22 U15537 ( .A1(n27465), .A2(n685), .B1(ram[2367]), .B2(n686), .ZN(
        n6608) );
  MOAI22 U15538 ( .A1(n29110), .A2(n687), .B1(ram[2368]), .B2(n688), .ZN(
        n6609) );
  MOAI22 U15539 ( .A1(n28875), .A2(n687), .B1(ram[2369]), .B2(n688), .ZN(
        n6610) );
  MOAI22 U15540 ( .A1(n28640), .A2(n687), .B1(ram[2370]), .B2(n688), .ZN(
        n6611) );
  MOAI22 U15541 ( .A1(n28405), .A2(n687), .B1(ram[2371]), .B2(n688), .ZN(
        n6612) );
  MOAI22 U15542 ( .A1(n28170), .A2(n687), .B1(ram[2372]), .B2(n688), .ZN(
        n6613) );
  MOAI22 U15543 ( .A1(n27935), .A2(n687), .B1(ram[2373]), .B2(n688), .ZN(
        n6614) );
  MOAI22 U15544 ( .A1(n27700), .A2(n687), .B1(ram[2374]), .B2(n688), .ZN(
        n6615) );
  MOAI22 U15545 ( .A1(n27465), .A2(n687), .B1(ram[2375]), .B2(n688), .ZN(
        n6616) );
  MOAI22 U15546 ( .A1(n29110), .A2(n689), .B1(ram[2376]), .B2(n690), .ZN(
        n6617) );
  MOAI22 U15547 ( .A1(n28875), .A2(n689), .B1(ram[2377]), .B2(n690), .ZN(
        n6618) );
  MOAI22 U15548 ( .A1(n28640), .A2(n689), .B1(ram[2378]), .B2(n690), .ZN(
        n6619) );
  MOAI22 U15549 ( .A1(n28405), .A2(n689), .B1(ram[2379]), .B2(n690), .ZN(
        n6620) );
  MOAI22 U15550 ( .A1(n28170), .A2(n689), .B1(ram[2380]), .B2(n690), .ZN(
        n6621) );
  MOAI22 U15551 ( .A1(n27935), .A2(n689), .B1(ram[2381]), .B2(n690), .ZN(
        n6622) );
  MOAI22 U15552 ( .A1(n27700), .A2(n689), .B1(ram[2382]), .B2(n690), .ZN(
        n6623) );
  MOAI22 U15553 ( .A1(n27465), .A2(n689), .B1(ram[2383]), .B2(n690), .ZN(
        n6624) );
  MOAI22 U15554 ( .A1(n29110), .A2(n691), .B1(ram[2384]), .B2(n692), .ZN(
        n6625) );
  MOAI22 U15555 ( .A1(n28875), .A2(n691), .B1(ram[2385]), .B2(n692), .ZN(
        n6626) );
  MOAI22 U15556 ( .A1(n28640), .A2(n691), .B1(ram[2386]), .B2(n692), .ZN(
        n6627) );
  MOAI22 U15557 ( .A1(n28405), .A2(n691), .B1(ram[2387]), .B2(n692), .ZN(
        n6628) );
  MOAI22 U15558 ( .A1(n28170), .A2(n691), .B1(ram[2388]), .B2(n692), .ZN(
        n6629) );
  MOAI22 U15559 ( .A1(n27935), .A2(n691), .B1(ram[2389]), .B2(n692), .ZN(
        n6630) );
  MOAI22 U15560 ( .A1(n27700), .A2(n691), .B1(ram[2390]), .B2(n692), .ZN(
        n6631) );
  MOAI22 U15561 ( .A1(n27465), .A2(n691), .B1(ram[2391]), .B2(n692), .ZN(
        n6632) );
  MOAI22 U15562 ( .A1(n29111), .A2(n693), .B1(ram[2392]), .B2(n694), .ZN(
        n6633) );
  MOAI22 U15563 ( .A1(n28876), .A2(n693), .B1(ram[2393]), .B2(n694), .ZN(
        n6634) );
  MOAI22 U15564 ( .A1(n28641), .A2(n693), .B1(ram[2394]), .B2(n694), .ZN(
        n6635) );
  MOAI22 U15565 ( .A1(n28406), .A2(n693), .B1(ram[2395]), .B2(n694), .ZN(
        n6636) );
  MOAI22 U15566 ( .A1(n28171), .A2(n693), .B1(ram[2396]), .B2(n694), .ZN(
        n6637) );
  MOAI22 U15567 ( .A1(n27936), .A2(n693), .B1(ram[2397]), .B2(n694), .ZN(
        n6638) );
  MOAI22 U15568 ( .A1(n27701), .A2(n693), .B1(ram[2398]), .B2(n694), .ZN(
        n6639) );
  MOAI22 U15569 ( .A1(n27466), .A2(n693), .B1(ram[2399]), .B2(n694), .ZN(
        n6640) );
  MOAI22 U15570 ( .A1(n29111), .A2(n695), .B1(ram[2400]), .B2(n696), .ZN(
        n6641) );
  MOAI22 U15571 ( .A1(n28876), .A2(n695), .B1(ram[2401]), .B2(n696), .ZN(
        n6642) );
  MOAI22 U15572 ( .A1(n28641), .A2(n695), .B1(ram[2402]), .B2(n696), .ZN(
        n6643) );
  MOAI22 U15573 ( .A1(n28406), .A2(n695), .B1(ram[2403]), .B2(n696), .ZN(
        n6644) );
  MOAI22 U15574 ( .A1(n28171), .A2(n695), .B1(ram[2404]), .B2(n696), .ZN(
        n6645) );
  MOAI22 U15575 ( .A1(n27936), .A2(n695), .B1(ram[2405]), .B2(n696), .ZN(
        n6646) );
  MOAI22 U15576 ( .A1(n27701), .A2(n695), .B1(ram[2406]), .B2(n696), .ZN(
        n6647) );
  MOAI22 U15577 ( .A1(n27466), .A2(n695), .B1(ram[2407]), .B2(n696), .ZN(
        n6648) );
  MOAI22 U15578 ( .A1(n29111), .A2(n697), .B1(ram[2408]), .B2(n698), .ZN(
        n6649) );
  MOAI22 U15579 ( .A1(n28876), .A2(n697), .B1(ram[2409]), .B2(n698), .ZN(
        n6650) );
  MOAI22 U15580 ( .A1(n28641), .A2(n697), .B1(ram[2410]), .B2(n698), .ZN(
        n6651) );
  MOAI22 U15581 ( .A1(n28406), .A2(n697), .B1(ram[2411]), .B2(n698), .ZN(
        n6652) );
  MOAI22 U15582 ( .A1(n28171), .A2(n697), .B1(ram[2412]), .B2(n698), .ZN(
        n6653) );
  MOAI22 U15583 ( .A1(n27936), .A2(n697), .B1(ram[2413]), .B2(n698), .ZN(
        n6654) );
  MOAI22 U15584 ( .A1(n27701), .A2(n697), .B1(ram[2414]), .B2(n698), .ZN(
        n6655) );
  MOAI22 U15585 ( .A1(n27466), .A2(n697), .B1(ram[2415]), .B2(n698), .ZN(
        n6656) );
  MOAI22 U15586 ( .A1(n29111), .A2(n699), .B1(ram[2416]), .B2(n700), .ZN(
        n6657) );
  MOAI22 U15587 ( .A1(n28876), .A2(n699), .B1(ram[2417]), .B2(n700), .ZN(
        n6658) );
  MOAI22 U15588 ( .A1(n28641), .A2(n699), .B1(ram[2418]), .B2(n700), .ZN(
        n6659) );
  MOAI22 U15589 ( .A1(n28406), .A2(n699), .B1(ram[2419]), .B2(n700), .ZN(
        n6660) );
  MOAI22 U15590 ( .A1(n28171), .A2(n699), .B1(ram[2420]), .B2(n700), .ZN(
        n6661) );
  MOAI22 U15591 ( .A1(n27936), .A2(n699), .B1(ram[2421]), .B2(n700), .ZN(
        n6662) );
  MOAI22 U15592 ( .A1(n27701), .A2(n699), .B1(ram[2422]), .B2(n700), .ZN(
        n6663) );
  MOAI22 U15593 ( .A1(n27466), .A2(n699), .B1(ram[2423]), .B2(n700), .ZN(
        n6664) );
  MOAI22 U15594 ( .A1(n29111), .A2(n701), .B1(ram[2424]), .B2(n702), .ZN(
        n6665) );
  MOAI22 U15595 ( .A1(n28876), .A2(n701), .B1(ram[2425]), .B2(n702), .ZN(
        n6666) );
  MOAI22 U15596 ( .A1(n28641), .A2(n701), .B1(ram[2426]), .B2(n702), .ZN(
        n6667) );
  MOAI22 U15597 ( .A1(n28406), .A2(n701), .B1(ram[2427]), .B2(n702), .ZN(
        n6668) );
  MOAI22 U15598 ( .A1(n28171), .A2(n701), .B1(ram[2428]), .B2(n702), .ZN(
        n6669) );
  MOAI22 U15599 ( .A1(n27936), .A2(n701), .B1(ram[2429]), .B2(n702), .ZN(
        n6670) );
  MOAI22 U15600 ( .A1(n27701), .A2(n701), .B1(ram[2430]), .B2(n702), .ZN(
        n6671) );
  MOAI22 U15601 ( .A1(n27466), .A2(n701), .B1(ram[2431]), .B2(n702), .ZN(
        n6672) );
  MOAI22 U15602 ( .A1(n29111), .A2(n703), .B1(ram[2432]), .B2(n704), .ZN(
        n6673) );
  MOAI22 U15603 ( .A1(n28876), .A2(n703), .B1(ram[2433]), .B2(n704), .ZN(
        n6674) );
  MOAI22 U15604 ( .A1(n28641), .A2(n703), .B1(ram[2434]), .B2(n704), .ZN(
        n6675) );
  MOAI22 U15605 ( .A1(n28406), .A2(n703), .B1(ram[2435]), .B2(n704), .ZN(
        n6676) );
  MOAI22 U15606 ( .A1(n28171), .A2(n703), .B1(ram[2436]), .B2(n704), .ZN(
        n6677) );
  MOAI22 U15607 ( .A1(n27936), .A2(n703), .B1(ram[2437]), .B2(n704), .ZN(
        n6678) );
  MOAI22 U15608 ( .A1(n27701), .A2(n703), .B1(ram[2438]), .B2(n704), .ZN(
        n6679) );
  MOAI22 U15609 ( .A1(n27466), .A2(n703), .B1(ram[2439]), .B2(n704), .ZN(
        n6680) );
  MOAI22 U15610 ( .A1(n29111), .A2(n705), .B1(ram[2440]), .B2(n706), .ZN(
        n6681) );
  MOAI22 U15611 ( .A1(n28876), .A2(n705), .B1(ram[2441]), .B2(n706), .ZN(
        n6682) );
  MOAI22 U15612 ( .A1(n28641), .A2(n705), .B1(ram[2442]), .B2(n706), .ZN(
        n6683) );
  MOAI22 U15613 ( .A1(n28406), .A2(n705), .B1(ram[2443]), .B2(n706), .ZN(
        n6684) );
  MOAI22 U15614 ( .A1(n28171), .A2(n705), .B1(ram[2444]), .B2(n706), .ZN(
        n6685) );
  MOAI22 U15615 ( .A1(n27936), .A2(n705), .B1(ram[2445]), .B2(n706), .ZN(
        n6686) );
  MOAI22 U15616 ( .A1(n27701), .A2(n705), .B1(ram[2446]), .B2(n706), .ZN(
        n6687) );
  MOAI22 U15617 ( .A1(n27466), .A2(n705), .B1(ram[2447]), .B2(n706), .ZN(
        n6688) );
  MOAI22 U15618 ( .A1(n29111), .A2(n707), .B1(ram[2448]), .B2(n708), .ZN(
        n6689) );
  MOAI22 U15619 ( .A1(n28876), .A2(n707), .B1(ram[2449]), .B2(n708), .ZN(
        n6690) );
  MOAI22 U15620 ( .A1(n28641), .A2(n707), .B1(ram[2450]), .B2(n708), .ZN(
        n6691) );
  MOAI22 U15621 ( .A1(n28406), .A2(n707), .B1(ram[2451]), .B2(n708), .ZN(
        n6692) );
  MOAI22 U15622 ( .A1(n28171), .A2(n707), .B1(ram[2452]), .B2(n708), .ZN(
        n6693) );
  MOAI22 U15623 ( .A1(n27936), .A2(n707), .B1(ram[2453]), .B2(n708), .ZN(
        n6694) );
  MOAI22 U15624 ( .A1(n27701), .A2(n707), .B1(ram[2454]), .B2(n708), .ZN(
        n6695) );
  MOAI22 U15625 ( .A1(n27466), .A2(n707), .B1(ram[2455]), .B2(n708), .ZN(
        n6696) );
  MOAI22 U15626 ( .A1(n29111), .A2(n709), .B1(ram[2456]), .B2(n710), .ZN(
        n6697) );
  MOAI22 U15627 ( .A1(n28876), .A2(n709), .B1(ram[2457]), .B2(n710), .ZN(
        n6698) );
  MOAI22 U15628 ( .A1(n28641), .A2(n709), .B1(ram[2458]), .B2(n710), .ZN(
        n6699) );
  MOAI22 U15629 ( .A1(n28406), .A2(n709), .B1(ram[2459]), .B2(n710), .ZN(
        n6700) );
  MOAI22 U15630 ( .A1(n28171), .A2(n709), .B1(ram[2460]), .B2(n710), .ZN(
        n6701) );
  MOAI22 U15631 ( .A1(n27936), .A2(n709), .B1(ram[2461]), .B2(n710), .ZN(
        n6702) );
  MOAI22 U15632 ( .A1(n27701), .A2(n709), .B1(ram[2462]), .B2(n710), .ZN(
        n6703) );
  MOAI22 U15633 ( .A1(n27466), .A2(n709), .B1(ram[2463]), .B2(n710), .ZN(
        n6704) );
  MOAI22 U15634 ( .A1(n29111), .A2(n711), .B1(ram[2464]), .B2(n712), .ZN(
        n6705) );
  MOAI22 U15635 ( .A1(n28876), .A2(n711), .B1(ram[2465]), .B2(n712), .ZN(
        n6706) );
  MOAI22 U15636 ( .A1(n28641), .A2(n711), .B1(ram[2466]), .B2(n712), .ZN(
        n6707) );
  MOAI22 U15637 ( .A1(n28406), .A2(n711), .B1(ram[2467]), .B2(n712), .ZN(
        n6708) );
  MOAI22 U15638 ( .A1(n28171), .A2(n711), .B1(ram[2468]), .B2(n712), .ZN(
        n6709) );
  MOAI22 U15639 ( .A1(n27936), .A2(n711), .B1(ram[2469]), .B2(n712), .ZN(
        n6710) );
  MOAI22 U15640 ( .A1(n27701), .A2(n711), .B1(ram[2470]), .B2(n712), .ZN(
        n6711) );
  MOAI22 U15641 ( .A1(n27466), .A2(n711), .B1(ram[2471]), .B2(n712), .ZN(
        n6712) );
  MOAI22 U15642 ( .A1(n29111), .A2(n713), .B1(ram[2472]), .B2(n714), .ZN(
        n6713) );
  MOAI22 U15643 ( .A1(n28876), .A2(n713), .B1(ram[2473]), .B2(n714), .ZN(
        n6714) );
  MOAI22 U15644 ( .A1(n28641), .A2(n713), .B1(ram[2474]), .B2(n714), .ZN(
        n6715) );
  MOAI22 U15645 ( .A1(n28406), .A2(n713), .B1(ram[2475]), .B2(n714), .ZN(
        n6716) );
  MOAI22 U15646 ( .A1(n28171), .A2(n713), .B1(ram[2476]), .B2(n714), .ZN(
        n6717) );
  MOAI22 U15647 ( .A1(n27936), .A2(n713), .B1(ram[2477]), .B2(n714), .ZN(
        n6718) );
  MOAI22 U15648 ( .A1(n27701), .A2(n713), .B1(ram[2478]), .B2(n714), .ZN(
        n6719) );
  MOAI22 U15649 ( .A1(n27466), .A2(n713), .B1(ram[2479]), .B2(n714), .ZN(
        n6720) );
  MOAI22 U15650 ( .A1(n29111), .A2(n715), .B1(ram[2480]), .B2(n716), .ZN(
        n6721) );
  MOAI22 U15651 ( .A1(n28876), .A2(n715), .B1(ram[2481]), .B2(n716), .ZN(
        n6722) );
  MOAI22 U15652 ( .A1(n28641), .A2(n715), .B1(ram[2482]), .B2(n716), .ZN(
        n6723) );
  MOAI22 U15653 ( .A1(n28406), .A2(n715), .B1(ram[2483]), .B2(n716), .ZN(
        n6724) );
  MOAI22 U15654 ( .A1(n28171), .A2(n715), .B1(ram[2484]), .B2(n716), .ZN(
        n6725) );
  MOAI22 U15655 ( .A1(n27936), .A2(n715), .B1(ram[2485]), .B2(n716), .ZN(
        n6726) );
  MOAI22 U15656 ( .A1(n27701), .A2(n715), .B1(ram[2486]), .B2(n716), .ZN(
        n6727) );
  MOAI22 U15657 ( .A1(n27466), .A2(n715), .B1(ram[2487]), .B2(n716), .ZN(
        n6728) );
  MOAI22 U15658 ( .A1(n29111), .A2(n717), .B1(ram[2488]), .B2(n718), .ZN(
        n6729) );
  MOAI22 U15659 ( .A1(n28876), .A2(n717), .B1(ram[2489]), .B2(n718), .ZN(
        n6730) );
  MOAI22 U15660 ( .A1(n28641), .A2(n717), .B1(ram[2490]), .B2(n718), .ZN(
        n6731) );
  MOAI22 U15661 ( .A1(n28406), .A2(n717), .B1(ram[2491]), .B2(n718), .ZN(
        n6732) );
  MOAI22 U15662 ( .A1(n28171), .A2(n717), .B1(ram[2492]), .B2(n718), .ZN(
        n6733) );
  MOAI22 U15663 ( .A1(n27936), .A2(n717), .B1(ram[2493]), .B2(n718), .ZN(
        n6734) );
  MOAI22 U15664 ( .A1(n27701), .A2(n717), .B1(ram[2494]), .B2(n718), .ZN(
        n6735) );
  MOAI22 U15665 ( .A1(n27466), .A2(n717), .B1(ram[2495]), .B2(n718), .ZN(
        n6736) );
  MOAI22 U15666 ( .A1(n29112), .A2(n719), .B1(ram[2496]), .B2(n720), .ZN(
        n6737) );
  MOAI22 U15667 ( .A1(n28877), .A2(n719), .B1(ram[2497]), .B2(n720), .ZN(
        n6738) );
  MOAI22 U15668 ( .A1(n28642), .A2(n719), .B1(ram[2498]), .B2(n720), .ZN(
        n6739) );
  MOAI22 U15669 ( .A1(n28407), .A2(n719), .B1(ram[2499]), .B2(n720), .ZN(
        n6740) );
  MOAI22 U15670 ( .A1(n28172), .A2(n719), .B1(ram[2500]), .B2(n720), .ZN(
        n6741) );
  MOAI22 U15671 ( .A1(n27937), .A2(n719), .B1(ram[2501]), .B2(n720), .ZN(
        n6742) );
  MOAI22 U15672 ( .A1(n27702), .A2(n719), .B1(ram[2502]), .B2(n720), .ZN(
        n6743) );
  MOAI22 U15673 ( .A1(n27467), .A2(n719), .B1(ram[2503]), .B2(n720), .ZN(
        n6744) );
  MOAI22 U15674 ( .A1(n29112), .A2(n721), .B1(ram[2504]), .B2(n722), .ZN(
        n6745) );
  MOAI22 U15675 ( .A1(n28877), .A2(n721), .B1(ram[2505]), .B2(n722), .ZN(
        n6746) );
  MOAI22 U15676 ( .A1(n28642), .A2(n721), .B1(ram[2506]), .B2(n722), .ZN(
        n6747) );
  MOAI22 U15677 ( .A1(n28407), .A2(n721), .B1(ram[2507]), .B2(n722), .ZN(
        n6748) );
  MOAI22 U15678 ( .A1(n28172), .A2(n721), .B1(ram[2508]), .B2(n722), .ZN(
        n6749) );
  MOAI22 U15679 ( .A1(n27937), .A2(n721), .B1(ram[2509]), .B2(n722), .ZN(
        n6750) );
  MOAI22 U15680 ( .A1(n27702), .A2(n721), .B1(ram[2510]), .B2(n722), .ZN(
        n6751) );
  MOAI22 U15681 ( .A1(n27467), .A2(n721), .B1(ram[2511]), .B2(n722), .ZN(
        n6752) );
  MOAI22 U15682 ( .A1(n29112), .A2(n723), .B1(ram[2512]), .B2(n724), .ZN(
        n6753) );
  MOAI22 U15683 ( .A1(n28877), .A2(n723), .B1(ram[2513]), .B2(n724), .ZN(
        n6754) );
  MOAI22 U15684 ( .A1(n28642), .A2(n723), .B1(ram[2514]), .B2(n724), .ZN(
        n6755) );
  MOAI22 U15685 ( .A1(n28407), .A2(n723), .B1(ram[2515]), .B2(n724), .ZN(
        n6756) );
  MOAI22 U15686 ( .A1(n28172), .A2(n723), .B1(ram[2516]), .B2(n724), .ZN(
        n6757) );
  MOAI22 U15687 ( .A1(n27937), .A2(n723), .B1(ram[2517]), .B2(n724), .ZN(
        n6758) );
  MOAI22 U15688 ( .A1(n27702), .A2(n723), .B1(ram[2518]), .B2(n724), .ZN(
        n6759) );
  MOAI22 U15689 ( .A1(n27467), .A2(n723), .B1(ram[2519]), .B2(n724), .ZN(
        n6760) );
  MOAI22 U15690 ( .A1(n29112), .A2(n725), .B1(ram[2520]), .B2(n726), .ZN(
        n6761) );
  MOAI22 U15691 ( .A1(n28877), .A2(n725), .B1(ram[2521]), .B2(n726), .ZN(
        n6762) );
  MOAI22 U15692 ( .A1(n28642), .A2(n725), .B1(ram[2522]), .B2(n726), .ZN(
        n6763) );
  MOAI22 U15693 ( .A1(n28407), .A2(n725), .B1(ram[2523]), .B2(n726), .ZN(
        n6764) );
  MOAI22 U15694 ( .A1(n28172), .A2(n725), .B1(ram[2524]), .B2(n726), .ZN(
        n6765) );
  MOAI22 U15695 ( .A1(n27937), .A2(n725), .B1(ram[2525]), .B2(n726), .ZN(
        n6766) );
  MOAI22 U15696 ( .A1(n27702), .A2(n725), .B1(ram[2526]), .B2(n726), .ZN(
        n6767) );
  MOAI22 U15697 ( .A1(n27467), .A2(n725), .B1(ram[2527]), .B2(n726), .ZN(
        n6768) );
  MOAI22 U15698 ( .A1(n29112), .A2(n727), .B1(ram[2528]), .B2(n728), .ZN(
        n6769) );
  MOAI22 U15699 ( .A1(n28877), .A2(n727), .B1(ram[2529]), .B2(n728), .ZN(
        n6770) );
  MOAI22 U15700 ( .A1(n28642), .A2(n727), .B1(ram[2530]), .B2(n728), .ZN(
        n6771) );
  MOAI22 U15701 ( .A1(n28407), .A2(n727), .B1(ram[2531]), .B2(n728), .ZN(
        n6772) );
  MOAI22 U15702 ( .A1(n28172), .A2(n727), .B1(ram[2532]), .B2(n728), .ZN(
        n6773) );
  MOAI22 U15703 ( .A1(n27937), .A2(n727), .B1(ram[2533]), .B2(n728), .ZN(
        n6774) );
  MOAI22 U15704 ( .A1(n27702), .A2(n727), .B1(ram[2534]), .B2(n728), .ZN(
        n6775) );
  MOAI22 U15705 ( .A1(n27467), .A2(n727), .B1(ram[2535]), .B2(n728), .ZN(
        n6776) );
  MOAI22 U15706 ( .A1(n29112), .A2(n729), .B1(ram[2536]), .B2(n730), .ZN(
        n6777) );
  MOAI22 U15707 ( .A1(n28877), .A2(n729), .B1(ram[2537]), .B2(n730), .ZN(
        n6778) );
  MOAI22 U15708 ( .A1(n28642), .A2(n729), .B1(ram[2538]), .B2(n730), .ZN(
        n6779) );
  MOAI22 U15709 ( .A1(n28407), .A2(n729), .B1(ram[2539]), .B2(n730), .ZN(
        n6780) );
  MOAI22 U15710 ( .A1(n28172), .A2(n729), .B1(ram[2540]), .B2(n730), .ZN(
        n6781) );
  MOAI22 U15711 ( .A1(n27937), .A2(n729), .B1(ram[2541]), .B2(n730), .ZN(
        n6782) );
  MOAI22 U15712 ( .A1(n27702), .A2(n729), .B1(ram[2542]), .B2(n730), .ZN(
        n6783) );
  MOAI22 U15713 ( .A1(n27467), .A2(n729), .B1(ram[2543]), .B2(n730), .ZN(
        n6784) );
  MOAI22 U15714 ( .A1(n29112), .A2(n731), .B1(ram[2544]), .B2(n732), .ZN(
        n6785) );
  MOAI22 U15715 ( .A1(n28877), .A2(n731), .B1(ram[2545]), .B2(n732), .ZN(
        n6786) );
  MOAI22 U15716 ( .A1(n28642), .A2(n731), .B1(ram[2546]), .B2(n732), .ZN(
        n6787) );
  MOAI22 U15717 ( .A1(n28407), .A2(n731), .B1(ram[2547]), .B2(n732), .ZN(
        n6788) );
  MOAI22 U15718 ( .A1(n28172), .A2(n731), .B1(ram[2548]), .B2(n732), .ZN(
        n6789) );
  MOAI22 U15719 ( .A1(n27937), .A2(n731), .B1(ram[2549]), .B2(n732), .ZN(
        n6790) );
  MOAI22 U15720 ( .A1(n27702), .A2(n731), .B1(ram[2550]), .B2(n732), .ZN(
        n6791) );
  MOAI22 U15721 ( .A1(n27467), .A2(n731), .B1(ram[2551]), .B2(n732), .ZN(
        n6792) );
  MOAI22 U15722 ( .A1(n29112), .A2(n733), .B1(ram[2552]), .B2(n734), .ZN(
        n6793) );
  MOAI22 U15723 ( .A1(n28877), .A2(n733), .B1(ram[2553]), .B2(n734), .ZN(
        n6794) );
  MOAI22 U15724 ( .A1(n28642), .A2(n733), .B1(ram[2554]), .B2(n734), .ZN(
        n6795) );
  MOAI22 U15725 ( .A1(n28407), .A2(n733), .B1(ram[2555]), .B2(n734), .ZN(
        n6796) );
  MOAI22 U15726 ( .A1(n28172), .A2(n733), .B1(ram[2556]), .B2(n734), .ZN(
        n6797) );
  MOAI22 U15727 ( .A1(n27937), .A2(n733), .B1(ram[2557]), .B2(n734), .ZN(
        n6798) );
  MOAI22 U15728 ( .A1(n27702), .A2(n733), .B1(ram[2558]), .B2(n734), .ZN(
        n6799) );
  MOAI22 U15729 ( .A1(n27467), .A2(n733), .B1(ram[2559]), .B2(n734), .ZN(
        n6800) );
  MOAI22 U15730 ( .A1(n29112), .A2(n736), .B1(ram[2560]), .B2(n737), .ZN(
        n6801) );
  MOAI22 U15731 ( .A1(n28877), .A2(n736), .B1(ram[2561]), .B2(n737), .ZN(
        n6802) );
  MOAI22 U15732 ( .A1(n28642), .A2(n736), .B1(ram[2562]), .B2(n737), .ZN(
        n6803) );
  MOAI22 U15733 ( .A1(n28407), .A2(n736), .B1(ram[2563]), .B2(n737), .ZN(
        n6804) );
  MOAI22 U15734 ( .A1(n28172), .A2(n736), .B1(ram[2564]), .B2(n737), .ZN(
        n6805) );
  MOAI22 U15735 ( .A1(n27937), .A2(n736), .B1(ram[2565]), .B2(n737), .ZN(
        n6806) );
  MOAI22 U15736 ( .A1(n27702), .A2(n736), .B1(ram[2566]), .B2(n737), .ZN(
        n6807) );
  MOAI22 U15737 ( .A1(n27467), .A2(n736), .B1(ram[2567]), .B2(n737), .ZN(
        n6808) );
  MOAI22 U15738 ( .A1(n29112), .A2(n739), .B1(ram[2568]), .B2(n740), .ZN(
        n6809) );
  MOAI22 U15739 ( .A1(n28877), .A2(n739), .B1(ram[2569]), .B2(n740), .ZN(
        n6810) );
  MOAI22 U15740 ( .A1(n28642), .A2(n739), .B1(ram[2570]), .B2(n740), .ZN(
        n6811) );
  MOAI22 U15741 ( .A1(n28407), .A2(n739), .B1(ram[2571]), .B2(n740), .ZN(
        n6812) );
  MOAI22 U15742 ( .A1(n28172), .A2(n739), .B1(ram[2572]), .B2(n740), .ZN(
        n6813) );
  MOAI22 U15743 ( .A1(n27937), .A2(n739), .B1(ram[2573]), .B2(n740), .ZN(
        n6814) );
  MOAI22 U15744 ( .A1(n27702), .A2(n739), .B1(ram[2574]), .B2(n740), .ZN(
        n6815) );
  MOAI22 U15745 ( .A1(n27467), .A2(n739), .B1(ram[2575]), .B2(n740), .ZN(
        n6816) );
  MOAI22 U15746 ( .A1(n29112), .A2(n741), .B1(ram[2576]), .B2(n742), .ZN(
        n6817) );
  MOAI22 U15747 ( .A1(n28877), .A2(n741), .B1(ram[2577]), .B2(n742), .ZN(
        n6818) );
  MOAI22 U15748 ( .A1(n28642), .A2(n741), .B1(ram[2578]), .B2(n742), .ZN(
        n6819) );
  MOAI22 U15749 ( .A1(n28407), .A2(n741), .B1(ram[2579]), .B2(n742), .ZN(
        n6820) );
  MOAI22 U15750 ( .A1(n28172), .A2(n741), .B1(ram[2580]), .B2(n742), .ZN(
        n6821) );
  MOAI22 U15751 ( .A1(n27937), .A2(n741), .B1(ram[2581]), .B2(n742), .ZN(
        n6822) );
  MOAI22 U15752 ( .A1(n27702), .A2(n741), .B1(ram[2582]), .B2(n742), .ZN(
        n6823) );
  MOAI22 U15753 ( .A1(n27467), .A2(n741), .B1(ram[2583]), .B2(n742), .ZN(
        n6824) );
  MOAI22 U15754 ( .A1(n29112), .A2(n743), .B1(ram[2584]), .B2(n744), .ZN(
        n6825) );
  MOAI22 U15755 ( .A1(n28877), .A2(n743), .B1(ram[2585]), .B2(n744), .ZN(
        n6826) );
  MOAI22 U15756 ( .A1(n28642), .A2(n743), .B1(ram[2586]), .B2(n744), .ZN(
        n6827) );
  MOAI22 U15757 ( .A1(n28407), .A2(n743), .B1(ram[2587]), .B2(n744), .ZN(
        n6828) );
  MOAI22 U15758 ( .A1(n28172), .A2(n743), .B1(ram[2588]), .B2(n744), .ZN(
        n6829) );
  MOAI22 U15759 ( .A1(n27937), .A2(n743), .B1(ram[2589]), .B2(n744), .ZN(
        n6830) );
  MOAI22 U15760 ( .A1(n27702), .A2(n743), .B1(ram[2590]), .B2(n744), .ZN(
        n6831) );
  MOAI22 U15761 ( .A1(n27467), .A2(n743), .B1(ram[2591]), .B2(n744), .ZN(
        n6832) );
  MOAI22 U15762 ( .A1(n29112), .A2(n745), .B1(ram[2592]), .B2(n746), .ZN(
        n6833) );
  MOAI22 U15763 ( .A1(n28877), .A2(n745), .B1(ram[2593]), .B2(n746), .ZN(
        n6834) );
  MOAI22 U15764 ( .A1(n28642), .A2(n745), .B1(ram[2594]), .B2(n746), .ZN(
        n6835) );
  MOAI22 U15765 ( .A1(n28407), .A2(n745), .B1(ram[2595]), .B2(n746), .ZN(
        n6836) );
  MOAI22 U15766 ( .A1(n28172), .A2(n745), .B1(ram[2596]), .B2(n746), .ZN(
        n6837) );
  MOAI22 U15767 ( .A1(n27937), .A2(n745), .B1(ram[2597]), .B2(n746), .ZN(
        n6838) );
  MOAI22 U15768 ( .A1(n27702), .A2(n745), .B1(ram[2598]), .B2(n746), .ZN(
        n6839) );
  MOAI22 U15769 ( .A1(n27467), .A2(n745), .B1(ram[2599]), .B2(n746), .ZN(
        n6840) );
  MOAI22 U15770 ( .A1(n29113), .A2(n747), .B1(ram[2600]), .B2(n748), .ZN(
        n6841) );
  MOAI22 U15771 ( .A1(n28878), .A2(n747), .B1(ram[2601]), .B2(n748), .ZN(
        n6842) );
  MOAI22 U15772 ( .A1(n28643), .A2(n747), .B1(ram[2602]), .B2(n748), .ZN(
        n6843) );
  MOAI22 U15773 ( .A1(n28408), .A2(n747), .B1(ram[2603]), .B2(n748), .ZN(
        n6844) );
  MOAI22 U15774 ( .A1(n28173), .A2(n747), .B1(ram[2604]), .B2(n748), .ZN(
        n6845) );
  MOAI22 U15775 ( .A1(n27938), .A2(n747), .B1(ram[2605]), .B2(n748), .ZN(
        n6846) );
  MOAI22 U15776 ( .A1(n27703), .A2(n747), .B1(ram[2606]), .B2(n748), .ZN(
        n6847) );
  MOAI22 U15777 ( .A1(n27468), .A2(n747), .B1(ram[2607]), .B2(n748), .ZN(
        n6848) );
  MOAI22 U15778 ( .A1(n29113), .A2(n749), .B1(ram[2608]), .B2(n750), .ZN(
        n6849) );
  MOAI22 U15779 ( .A1(n28878), .A2(n749), .B1(ram[2609]), .B2(n750), .ZN(
        n6850) );
  MOAI22 U15780 ( .A1(n28643), .A2(n749), .B1(ram[2610]), .B2(n750), .ZN(
        n6851) );
  MOAI22 U15781 ( .A1(n28408), .A2(n749), .B1(ram[2611]), .B2(n750), .ZN(
        n6852) );
  MOAI22 U15782 ( .A1(n28173), .A2(n749), .B1(ram[2612]), .B2(n750), .ZN(
        n6853) );
  MOAI22 U15783 ( .A1(n27938), .A2(n749), .B1(ram[2613]), .B2(n750), .ZN(
        n6854) );
  MOAI22 U15784 ( .A1(n27703), .A2(n749), .B1(ram[2614]), .B2(n750), .ZN(
        n6855) );
  MOAI22 U15785 ( .A1(n27468), .A2(n749), .B1(ram[2615]), .B2(n750), .ZN(
        n6856) );
  MOAI22 U15786 ( .A1(n29113), .A2(n751), .B1(ram[2616]), .B2(n752), .ZN(
        n6857) );
  MOAI22 U15787 ( .A1(n28878), .A2(n751), .B1(ram[2617]), .B2(n752), .ZN(
        n6858) );
  MOAI22 U15788 ( .A1(n28643), .A2(n751), .B1(ram[2618]), .B2(n752), .ZN(
        n6859) );
  MOAI22 U15789 ( .A1(n28408), .A2(n751), .B1(ram[2619]), .B2(n752), .ZN(
        n6860) );
  MOAI22 U15790 ( .A1(n28173), .A2(n751), .B1(ram[2620]), .B2(n752), .ZN(
        n6861) );
  MOAI22 U15791 ( .A1(n27938), .A2(n751), .B1(ram[2621]), .B2(n752), .ZN(
        n6862) );
  MOAI22 U15792 ( .A1(n27703), .A2(n751), .B1(ram[2622]), .B2(n752), .ZN(
        n6863) );
  MOAI22 U15793 ( .A1(n27468), .A2(n751), .B1(ram[2623]), .B2(n752), .ZN(
        n6864) );
  MOAI22 U15794 ( .A1(n29113), .A2(n753), .B1(ram[2624]), .B2(n754), .ZN(
        n6865) );
  MOAI22 U15795 ( .A1(n28878), .A2(n753), .B1(ram[2625]), .B2(n754), .ZN(
        n6866) );
  MOAI22 U15796 ( .A1(n28643), .A2(n753), .B1(ram[2626]), .B2(n754), .ZN(
        n6867) );
  MOAI22 U15797 ( .A1(n28408), .A2(n753), .B1(ram[2627]), .B2(n754), .ZN(
        n6868) );
  MOAI22 U15798 ( .A1(n28173), .A2(n753), .B1(ram[2628]), .B2(n754), .ZN(
        n6869) );
  MOAI22 U15799 ( .A1(n27938), .A2(n753), .B1(ram[2629]), .B2(n754), .ZN(
        n6870) );
  MOAI22 U15800 ( .A1(n27703), .A2(n753), .B1(ram[2630]), .B2(n754), .ZN(
        n6871) );
  MOAI22 U15801 ( .A1(n27468), .A2(n753), .B1(ram[2631]), .B2(n754), .ZN(
        n6872) );
  MOAI22 U15802 ( .A1(n29113), .A2(n755), .B1(ram[2632]), .B2(n756), .ZN(
        n6873) );
  MOAI22 U15803 ( .A1(n28878), .A2(n755), .B1(ram[2633]), .B2(n756), .ZN(
        n6874) );
  MOAI22 U15804 ( .A1(n28643), .A2(n755), .B1(ram[2634]), .B2(n756), .ZN(
        n6875) );
  MOAI22 U15805 ( .A1(n28408), .A2(n755), .B1(ram[2635]), .B2(n756), .ZN(
        n6876) );
  MOAI22 U15806 ( .A1(n28173), .A2(n755), .B1(ram[2636]), .B2(n756), .ZN(
        n6877) );
  MOAI22 U15807 ( .A1(n27938), .A2(n755), .B1(ram[2637]), .B2(n756), .ZN(
        n6878) );
  MOAI22 U15808 ( .A1(n27703), .A2(n755), .B1(ram[2638]), .B2(n756), .ZN(
        n6879) );
  MOAI22 U15809 ( .A1(n27468), .A2(n755), .B1(ram[2639]), .B2(n756), .ZN(
        n6880) );
  MOAI22 U15810 ( .A1(n29113), .A2(n757), .B1(ram[2640]), .B2(n758), .ZN(
        n6881) );
  MOAI22 U15811 ( .A1(n28878), .A2(n757), .B1(ram[2641]), .B2(n758), .ZN(
        n6882) );
  MOAI22 U15812 ( .A1(n28643), .A2(n757), .B1(ram[2642]), .B2(n758), .ZN(
        n6883) );
  MOAI22 U15813 ( .A1(n28408), .A2(n757), .B1(ram[2643]), .B2(n758), .ZN(
        n6884) );
  MOAI22 U15814 ( .A1(n28173), .A2(n757), .B1(ram[2644]), .B2(n758), .ZN(
        n6885) );
  MOAI22 U15815 ( .A1(n27938), .A2(n757), .B1(ram[2645]), .B2(n758), .ZN(
        n6886) );
  MOAI22 U15816 ( .A1(n27703), .A2(n757), .B1(ram[2646]), .B2(n758), .ZN(
        n6887) );
  MOAI22 U15817 ( .A1(n27468), .A2(n757), .B1(ram[2647]), .B2(n758), .ZN(
        n6888) );
  MOAI22 U15818 ( .A1(n29113), .A2(n759), .B1(ram[2648]), .B2(n760), .ZN(
        n6889) );
  MOAI22 U15819 ( .A1(n28878), .A2(n759), .B1(ram[2649]), .B2(n760), .ZN(
        n6890) );
  MOAI22 U15820 ( .A1(n28643), .A2(n759), .B1(ram[2650]), .B2(n760), .ZN(
        n6891) );
  MOAI22 U15821 ( .A1(n28408), .A2(n759), .B1(ram[2651]), .B2(n760), .ZN(
        n6892) );
  MOAI22 U15822 ( .A1(n28173), .A2(n759), .B1(ram[2652]), .B2(n760), .ZN(
        n6893) );
  MOAI22 U15823 ( .A1(n27938), .A2(n759), .B1(ram[2653]), .B2(n760), .ZN(
        n6894) );
  MOAI22 U15824 ( .A1(n27703), .A2(n759), .B1(ram[2654]), .B2(n760), .ZN(
        n6895) );
  MOAI22 U15825 ( .A1(n27468), .A2(n759), .B1(ram[2655]), .B2(n760), .ZN(
        n6896) );
  MOAI22 U15826 ( .A1(n29113), .A2(n761), .B1(ram[2656]), .B2(n762), .ZN(
        n6897) );
  MOAI22 U15827 ( .A1(n28878), .A2(n761), .B1(ram[2657]), .B2(n762), .ZN(
        n6898) );
  MOAI22 U15828 ( .A1(n28643), .A2(n761), .B1(ram[2658]), .B2(n762), .ZN(
        n6899) );
  MOAI22 U15829 ( .A1(n28408), .A2(n761), .B1(ram[2659]), .B2(n762), .ZN(
        n6900) );
  MOAI22 U15830 ( .A1(n28173), .A2(n761), .B1(ram[2660]), .B2(n762), .ZN(
        n6901) );
  MOAI22 U15831 ( .A1(n27938), .A2(n761), .B1(ram[2661]), .B2(n762), .ZN(
        n6902) );
  MOAI22 U15832 ( .A1(n27703), .A2(n761), .B1(ram[2662]), .B2(n762), .ZN(
        n6903) );
  MOAI22 U15833 ( .A1(n27468), .A2(n761), .B1(ram[2663]), .B2(n762), .ZN(
        n6904) );
  MOAI22 U15834 ( .A1(n29113), .A2(n763), .B1(ram[2664]), .B2(n764), .ZN(
        n6905) );
  MOAI22 U15835 ( .A1(n28878), .A2(n763), .B1(ram[2665]), .B2(n764), .ZN(
        n6906) );
  MOAI22 U15836 ( .A1(n28643), .A2(n763), .B1(ram[2666]), .B2(n764), .ZN(
        n6907) );
  MOAI22 U15837 ( .A1(n28408), .A2(n763), .B1(ram[2667]), .B2(n764), .ZN(
        n6908) );
  MOAI22 U15838 ( .A1(n28173), .A2(n763), .B1(ram[2668]), .B2(n764), .ZN(
        n6909) );
  MOAI22 U15839 ( .A1(n27938), .A2(n763), .B1(ram[2669]), .B2(n764), .ZN(
        n6910) );
  MOAI22 U15840 ( .A1(n27703), .A2(n763), .B1(ram[2670]), .B2(n764), .ZN(
        n6911) );
  MOAI22 U15841 ( .A1(n27468), .A2(n763), .B1(ram[2671]), .B2(n764), .ZN(
        n6912) );
  MOAI22 U15842 ( .A1(n29113), .A2(n765), .B1(ram[2672]), .B2(n766), .ZN(
        n6913) );
  MOAI22 U15843 ( .A1(n28878), .A2(n765), .B1(ram[2673]), .B2(n766), .ZN(
        n6914) );
  MOAI22 U15844 ( .A1(n28643), .A2(n765), .B1(ram[2674]), .B2(n766), .ZN(
        n6915) );
  MOAI22 U15845 ( .A1(n28408), .A2(n765), .B1(ram[2675]), .B2(n766), .ZN(
        n6916) );
  MOAI22 U15846 ( .A1(n28173), .A2(n765), .B1(ram[2676]), .B2(n766), .ZN(
        n6917) );
  MOAI22 U15847 ( .A1(n27938), .A2(n765), .B1(ram[2677]), .B2(n766), .ZN(
        n6918) );
  MOAI22 U15848 ( .A1(n27703), .A2(n765), .B1(ram[2678]), .B2(n766), .ZN(
        n6919) );
  MOAI22 U15849 ( .A1(n27468), .A2(n765), .B1(ram[2679]), .B2(n766), .ZN(
        n6920) );
  MOAI22 U15850 ( .A1(n29113), .A2(n767), .B1(ram[2680]), .B2(n768), .ZN(
        n6921) );
  MOAI22 U15851 ( .A1(n28878), .A2(n767), .B1(ram[2681]), .B2(n768), .ZN(
        n6922) );
  MOAI22 U15852 ( .A1(n28643), .A2(n767), .B1(ram[2682]), .B2(n768), .ZN(
        n6923) );
  MOAI22 U15853 ( .A1(n28408), .A2(n767), .B1(ram[2683]), .B2(n768), .ZN(
        n6924) );
  MOAI22 U15854 ( .A1(n28173), .A2(n767), .B1(ram[2684]), .B2(n768), .ZN(
        n6925) );
  MOAI22 U15855 ( .A1(n27938), .A2(n767), .B1(ram[2685]), .B2(n768), .ZN(
        n6926) );
  MOAI22 U15856 ( .A1(n27703), .A2(n767), .B1(ram[2686]), .B2(n768), .ZN(
        n6927) );
  MOAI22 U15857 ( .A1(n27468), .A2(n767), .B1(ram[2687]), .B2(n768), .ZN(
        n6928) );
  MOAI22 U15858 ( .A1(n29113), .A2(n769), .B1(ram[2688]), .B2(n770), .ZN(
        n6929) );
  MOAI22 U15859 ( .A1(n28878), .A2(n769), .B1(ram[2689]), .B2(n770), .ZN(
        n6930) );
  MOAI22 U15860 ( .A1(n28643), .A2(n769), .B1(ram[2690]), .B2(n770), .ZN(
        n6931) );
  MOAI22 U15861 ( .A1(n28408), .A2(n769), .B1(ram[2691]), .B2(n770), .ZN(
        n6932) );
  MOAI22 U15862 ( .A1(n28173), .A2(n769), .B1(ram[2692]), .B2(n770), .ZN(
        n6933) );
  MOAI22 U15863 ( .A1(n27938), .A2(n769), .B1(ram[2693]), .B2(n770), .ZN(
        n6934) );
  MOAI22 U15864 ( .A1(n27703), .A2(n769), .B1(ram[2694]), .B2(n770), .ZN(
        n6935) );
  MOAI22 U15865 ( .A1(n27468), .A2(n769), .B1(ram[2695]), .B2(n770), .ZN(
        n6936) );
  MOAI22 U15866 ( .A1(n29113), .A2(n771), .B1(ram[2696]), .B2(n772), .ZN(
        n6937) );
  MOAI22 U15867 ( .A1(n28878), .A2(n771), .B1(ram[2697]), .B2(n772), .ZN(
        n6938) );
  MOAI22 U15868 ( .A1(n28643), .A2(n771), .B1(ram[2698]), .B2(n772), .ZN(
        n6939) );
  MOAI22 U15869 ( .A1(n28408), .A2(n771), .B1(ram[2699]), .B2(n772), .ZN(
        n6940) );
  MOAI22 U15870 ( .A1(n28173), .A2(n771), .B1(ram[2700]), .B2(n772), .ZN(
        n6941) );
  MOAI22 U15871 ( .A1(n27938), .A2(n771), .B1(ram[2701]), .B2(n772), .ZN(
        n6942) );
  MOAI22 U15872 ( .A1(n27703), .A2(n771), .B1(ram[2702]), .B2(n772), .ZN(
        n6943) );
  MOAI22 U15873 ( .A1(n27468), .A2(n771), .B1(ram[2703]), .B2(n772), .ZN(
        n6944) );
  MOAI22 U15874 ( .A1(n29114), .A2(n773), .B1(ram[2704]), .B2(n774), .ZN(
        n6945) );
  MOAI22 U15875 ( .A1(n28879), .A2(n773), .B1(ram[2705]), .B2(n774), .ZN(
        n6946) );
  MOAI22 U15876 ( .A1(n28644), .A2(n773), .B1(ram[2706]), .B2(n774), .ZN(
        n6947) );
  MOAI22 U15877 ( .A1(n28409), .A2(n773), .B1(ram[2707]), .B2(n774), .ZN(
        n6948) );
  MOAI22 U15878 ( .A1(n28174), .A2(n773), .B1(ram[2708]), .B2(n774), .ZN(
        n6949) );
  MOAI22 U15879 ( .A1(n27939), .A2(n773), .B1(ram[2709]), .B2(n774), .ZN(
        n6950) );
  MOAI22 U15880 ( .A1(n27704), .A2(n773), .B1(ram[2710]), .B2(n774), .ZN(
        n6951) );
  MOAI22 U15881 ( .A1(n27469), .A2(n773), .B1(ram[2711]), .B2(n774), .ZN(
        n6952) );
  MOAI22 U15882 ( .A1(n29114), .A2(n775), .B1(ram[2712]), .B2(n776), .ZN(
        n6953) );
  MOAI22 U15883 ( .A1(n28879), .A2(n775), .B1(ram[2713]), .B2(n776), .ZN(
        n6954) );
  MOAI22 U15884 ( .A1(n28644), .A2(n775), .B1(ram[2714]), .B2(n776), .ZN(
        n6955) );
  MOAI22 U15885 ( .A1(n28409), .A2(n775), .B1(ram[2715]), .B2(n776), .ZN(
        n6956) );
  MOAI22 U15886 ( .A1(n28174), .A2(n775), .B1(ram[2716]), .B2(n776), .ZN(
        n6957) );
  MOAI22 U15887 ( .A1(n27939), .A2(n775), .B1(ram[2717]), .B2(n776), .ZN(
        n6958) );
  MOAI22 U15888 ( .A1(n27704), .A2(n775), .B1(ram[2718]), .B2(n776), .ZN(
        n6959) );
  MOAI22 U15889 ( .A1(n27469), .A2(n775), .B1(ram[2719]), .B2(n776), .ZN(
        n6960) );
  MOAI22 U15890 ( .A1(n29114), .A2(n777), .B1(ram[2720]), .B2(n778), .ZN(
        n6961) );
  MOAI22 U15891 ( .A1(n28879), .A2(n777), .B1(ram[2721]), .B2(n778), .ZN(
        n6962) );
  MOAI22 U15892 ( .A1(n28644), .A2(n777), .B1(ram[2722]), .B2(n778), .ZN(
        n6963) );
  MOAI22 U15893 ( .A1(n28409), .A2(n777), .B1(ram[2723]), .B2(n778), .ZN(
        n6964) );
  MOAI22 U15894 ( .A1(n28174), .A2(n777), .B1(ram[2724]), .B2(n778), .ZN(
        n6965) );
  MOAI22 U15895 ( .A1(n27939), .A2(n777), .B1(ram[2725]), .B2(n778), .ZN(
        n6966) );
  MOAI22 U15896 ( .A1(n27704), .A2(n777), .B1(ram[2726]), .B2(n778), .ZN(
        n6967) );
  MOAI22 U15897 ( .A1(n27469), .A2(n777), .B1(ram[2727]), .B2(n778), .ZN(
        n6968) );
  MOAI22 U15898 ( .A1(n29114), .A2(n779), .B1(ram[2728]), .B2(n780), .ZN(
        n6969) );
  MOAI22 U15899 ( .A1(n28879), .A2(n779), .B1(ram[2729]), .B2(n780), .ZN(
        n6970) );
  MOAI22 U15900 ( .A1(n28644), .A2(n779), .B1(ram[2730]), .B2(n780), .ZN(
        n6971) );
  MOAI22 U15901 ( .A1(n28409), .A2(n779), .B1(ram[2731]), .B2(n780), .ZN(
        n6972) );
  MOAI22 U15902 ( .A1(n28174), .A2(n779), .B1(ram[2732]), .B2(n780), .ZN(
        n6973) );
  MOAI22 U15903 ( .A1(n27939), .A2(n779), .B1(ram[2733]), .B2(n780), .ZN(
        n6974) );
  MOAI22 U15904 ( .A1(n27704), .A2(n779), .B1(ram[2734]), .B2(n780), .ZN(
        n6975) );
  MOAI22 U15905 ( .A1(n27469), .A2(n779), .B1(ram[2735]), .B2(n780), .ZN(
        n6976) );
  MOAI22 U15906 ( .A1(n29114), .A2(n781), .B1(ram[2736]), .B2(n782), .ZN(
        n6977) );
  MOAI22 U15907 ( .A1(n28879), .A2(n781), .B1(ram[2737]), .B2(n782), .ZN(
        n6978) );
  MOAI22 U15908 ( .A1(n28644), .A2(n781), .B1(ram[2738]), .B2(n782), .ZN(
        n6979) );
  MOAI22 U15909 ( .A1(n28409), .A2(n781), .B1(ram[2739]), .B2(n782), .ZN(
        n6980) );
  MOAI22 U15910 ( .A1(n28174), .A2(n781), .B1(ram[2740]), .B2(n782), .ZN(
        n6981) );
  MOAI22 U15911 ( .A1(n27939), .A2(n781), .B1(ram[2741]), .B2(n782), .ZN(
        n6982) );
  MOAI22 U15912 ( .A1(n27704), .A2(n781), .B1(ram[2742]), .B2(n782), .ZN(
        n6983) );
  MOAI22 U15913 ( .A1(n27469), .A2(n781), .B1(ram[2743]), .B2(n782), .ZN(
        n6984) );
  MOAI22 U15914 ( .A1(n29114), .A2(n783), .B1(ram[2744]), .B2(n784), .ZN(
        n6985) );
  MOAI22 U15915 ( .A1(n28879), .A2(n783), .B1(ram[2745]), .B2(n784), .ZN(
        n6986) );
  MOAI22 U15916 ( .A1(n28644), .A2(n783), .B1(ram[2746]), .B2(n784), .ZN(
        n6987) );
  MOAI22 U15917 ( .A1(n28409), .A2(n783), .B1(ram[2747]), .B2(n784), .ZN(
        n6988) );
  MOAI22 U15918 ( .A1(n28174), .A2(n783), .B1(ram[2748]), .B2(n784), .ZN(
        n6989) );
  MOAI22 U15919 ( .A1(n27939), .A2(n783), .B1(ram[2749]), .B2(n784), .ZN(
        n6990) );
  MOAI22 U15920 ( .A1(n27704), .A2(n783), .B1(ram[2750]), .B2(n784), .ZN(
        n6991) );
  MOAI22 U15921 ( .A1(n27469), .A2(n783), .B1(ram[2751]), .B2(n784), .ZN(
        n6992) );
  MOAI22 U15922 ( .A1(n29114), .A2(n785), .B1(ram[2752]), .B2(n786), .ZN(
        n6993) );
  MOAI22 U15923 ( .A1(n28879), .A2(n785), .B1(ram[2753]), .B2(n786), .ZN(
        n6994) );
  MOAI22 U15924 ( .A1(n28644), .A2(n785), .B1(ram[2754]), .B2(n786), .ZN(
        n6995) );
  MOAI22 U15925 ( .A1(n28409), .A2(n785), .B1(ram[2755]), .B2(n786), .ZN(
        n6996) );
  MOAI22 U15926 ( .A1(n28174), .A2(n785), .B1(ram[2756]), .B2(n786), .ZN(
        n6997) );
  MOAI22 U15927 ( .A1(n27939), .A2(n785), .B1(ram[2757]), .B2(n786), .ZN(
        n6998) );
  MOAI22 U15928 ( .A1(n27704), .A2(n785), .B1(ram[2758]), .B2(n786), .ZN(
        n6999) );
  MOAI22 U15929 ( .A1(n27469), .A2(n785), .B1(ram[2759]), .B2(n786), .ZN(
        n7000) );
  MOAI22 U15930 ( .A1(n29114), .A2(n787), .B1(ram[2760]), .B2(n788), .ZN(
        n7001) );
  MOAI22 U15931 ( .A1(n28879), .A2(n787), .B1(ram[2761]), .B2(n788), .ZN(
        n7002) );
  MOAI22 U15932 ( .A1(n28644), .A2(n787), .B1(ram[2762]), .B2(n788), .ZN(
        n7003) );
  MOAI22 U15933 ( .A1(n28409), .A2(n787), .B1(ram[2763]), .B2(n788), .ZN(
        n7004) );
  MOAI22 U15934 ( .A1(n28174), .A2(n787), .B1(ram[2764]), .B2(n788), .ZN(
        n7005) );
  MOAI22 U15935 ( .A1(n27939), .A2(n787), .B1(ram[2765]), .B2(n788), .ZN(
        n7006) );
  MOAI22 U15936 ( .A1(n27704), .A2(n787), .B1(ram[2766]), .B2(n788), .ZN(
        n7007) );
  MOAI22 U15937 ( .A1(n27469), .A2(n787), .B1(ram[2767]), .B2(n788), .ZN(
        n7008) );
  MOAI22 U15938 ( .A1(n29114), .A2(n789), .B1(ram[2768]), .B2(n790), .ZN(
        n7009) );
  MOAI22 U15939 ( .A1(n28879), .A2(n789), .B1(ram[2769]), .B2(n790), .ZN(
        n7010) );
  MOAI22 U15940 ( .A1(n28644), .A2(n789), .B1(ram[2770]), .B2(n790), .ZN(
        n7011) );
  MOAI22 U15941 ( .A1(n28409), .A2(n789), .B1(ram[2771]), .B2(n790), .ZN(
        n7012) );
  MOAI22 U15942 ( .A1(n28174), .A2(n789), .B1(ram[2772]), .B2(n790), .ZN(
        n7013) );
  MOAI22 U15943 ( .A1(n27939), .A2(n789), .B1(ram[2773]), .B2(n790), .ZN(
        n7014) );
  MOAI22 U15944 ( .A1(n27704), .A2(n789), .B1(ram[2774]), .B2(n790), .ZN(
        n7015) );
  MOAI22 U15945 ( .A1(n27469), .A2(n789), .B1(ram[2775]), .B2(n790), .ZN(
        n7016) );
  MOAI22 U15946 ( .A1(n29114), .A2(n791), .B1(ram[2776]), .B2(n792), .ZN(
        n7017) );
  MOAI22 U15947 ( .A1(n28879), .A2(n791), .B1(ram[2777]), .B2(n792), .ZN(
        n7018) );
  MOAI22 U15948 ( .A1(n28644), .A2(n791), .B1(ram[2778]), .B2(n792), .ZN(
        n7019) );
  MOAI22 U15949 ( .A1(n28409), .A2(n791), .B1(ram[2779]), .B2(n792), .ZN(
        n7020) );
  MOAI22 U15950 ( .A1(n28174), .A2(n791), .B1(ram[2780]), .B2(n792), .ZN(
        n7021) );
  MOAI22 U15951 ( .A1(n27939), .A2(n791), .B1(ram[2781]), .B2(n792), .ZN(
        n7022) );
  MOAI22 U15952 ( .A1(n27704), .A2(n791), .B1(ram[2782]), .B2(n792), .ZN(
        n7023) );
  MOAI22 U15953 ( .A1(n27469), .A2(n791), .B1(ram[2783]), .B2(n792), .ZN(
        n7024) );
  MOAI22 U15954 ( .A1(n29114), .A2(n793), .B1(ram[2784]), .B2(n794), .ZN(
        n7025) );
  MOAI22 U15955 ( .A1(n28879), .A2(n793), .B1(ram[2785]), .B2(n794), .ZN(
        n7026) );
  MOAI22 U15956 ( .A1(n28644), .A2(n793), .B1(ram[2786]), .B2(n794), .ZN(
        n7027) );
  MOAI22 U15957 ( .A1(n28409), .A2(n793), .B1(ram[2787]), .B2(n794), .ZN(
        n7028) );
  MOAI22 U15958 ( .A1(n28174), .A2(n793), .B1(ram[2788]), .B2(n794), .ZN(
        n7029) );
  MOAI22 U15959 ( .A1(n27939), .A2(n793), .B1(ram[2789]), .B2(n794), .ZN(
        n7030) );
  MOAI22 U15960 ( .A1(n27704), .A2(n793), .B1(ram[2790]), .B2(n794), .ZN(
        n7031) );
  MOAI22 U15961 ( .A1(n27469), .A2(n793), .B1(ram[2791]), .B2(n794), .ZN(
        n7032) );
  MOAI22 U15962 ( .A1(n29114), .A2(n795), .B1(ram[2792]), .B2(n796), .ZN(
        n7033) );
  MOAI22 U15963 ( .A1(n28879), .A2(n795), .B1(ram[2793]), .B2(n796), .ZN(
        n7034) );
  MOAI22 U15964 ( .A1(n28644), .A2(n795), .B1(ram[2794]), .B2(n796), .ZN(
        n7035) );
  MOAI22 U15965 ( .A1(n28409), .A2(n795), .B1(ram[2795]), .B2(n796), .ZN(
        n7036) );
  MOAI22 U15966 ( .A1(n28174), .A2(n795), .B1(ram[2796]), .B2(n796), .ZN(
        n7037) );
  MOAI22 U15967 ( .A1(n27939), .A2(n795), .B1(ram[2797]), .B2(n796), .ZN(
        n7038) );
  MOAI22 U15968 ( .A1(n27704), .A2(n795), .B1(ram[2798]), .B2(n796), .ZN(
        n7039) );
  MOAI22 U15969 ( .A1(n27469), .A2(n795), .B1(ram[2799]), .B2(n796), .ZN(
        n7040) );
  MOAI22 U15970 ( .A1(n29114), .A2(n797), .B1(ram[2800]), .B2(n798), .ZN(
        n7041) );
  MOAI22 U15971 ( .A1(n28879), .A2(n797), .B1(ram[2801]), .B2(n798), .ZN(
        n7042) );
  MOAI22 U15972 ( .A1(n28644), .A2(n797), .B1(ram[2802]), .B2(n798), .ZN(
        n7043) );
  MOAI22 U15973 ( .A1(n28409), .A2(n797), .B1(ram[2803]), .B2(n798), .ZN(
        n7044) );
  MOAI22 U15974 ( .A1(n28174), .A2(n797), .B1(ram[2804]), .B2(n798), .ZN(
        n7045) );
  MOAI22 U15975 ( .A1(n27939), .A2(n797), .B1(ram[2805]), .B2(n798), .ZN(
        n7046) );
  MOAI22 U15976 ( .A1(n27704), .A2(n797), .B1(ram[2806]), .B2(n798), .ZN(
        n7047) );
  MOAI22 U15977 ( .A1(n27469), .A2(n797), .B1(ram[2807]), .B2(n798), .ZN(
        n7048) );
  MOAI22 U15978 ( .A1(n29115), .A2(n799), .B1(ram[2808]), .B2(n800), .ZN(
        n7049) );
  MOAI22 U15979 ( .A1(n28880), .A2(n799), .B1(ram[2809]), .B2(n800), .ZN(
        n7050) );
  MOAI22 U15980 ( .A1(n28645), .A2(n799), .B1(ram[2810]), .B2(n800), .ZN(
        n7051) );
  MOAI22 U15981 ( .A1(n28410), .A2(n799), .B1(ram[2811]), .B2(n800), .ZN(
        n7052) );
  MOAI22 U15982 ( .A1(n28175), .A2(n799), .B1(ram[2812]), .B2(n800), .ZN(
        n7053) );
  MOAI22 U15983 ( .A1(n27940), .A2(n799), .B1(ram[2813]), .B2(n800), .ZN(
        n7054) );
  MOAI22 U15984 ( .A1(n27705), .A2(n799), .B1(ram[2814]), .B2(n800), .ZN(
        n7055) );
  MOAI22 U15985 ( .A1(n27470), .A2(n799), .B1(ram[2815]), .B2(n800), .ZN(
        n7056) );
  MOAI22 U15986 ( .A1(n29115), .A2(n801), .B1(ram[2816]), .B2(n802), .ZN(
        n7057) );
  MOAI22 U15987 ( .A1(n28880), .A2(n801), .B1(ram[2817]), .B2(n802), .ZN(
        n7058) );
  MOAI22 U15988 ( .A1(n28645), .A2(n801), .B1(ram[2818]), .B2(n802), .ZN(
        n7059) );
  MOAI22 U15989 ( .A1(n28410), .A2(n801), .B1(ram[2819]), .B2(n802), .ZN(
        n7060) );
  MOAI22 U15990 ( .A1(n28175), .A2(n801), .B1(ram[2820]), .B2(n802), .ZN(
        n7061) );
  MOAI22 U15991 ( .A1(n27940), .A2(n801), .B1(ram[2821]), .B2(n802), .ZN(
        n7062) );
  MOAI22 U15992 ( .A1(n27705), .A2(n801), .B1(ram[2822]), .B2(n802), .ZN(
        n7063) );
  MOAI22 U15993 ( .A1(n27470), .A2(n801), .B1(ram[2823]), .B2(n802), .ZN(
        n7064) );
  MOAI22 U15994 ( .A1(n29115), .A2(n803), .B1(ram[2824]), .B2(n804), .ZN(
        n7065) );
  MOAI22 U15995 ( .A1(n28880), .A2(n803), .B1(ram[2825]), .B2(n804), .ZN(
        n7066) );
  MOAI22 U15996 ( .A1(n28645), .A2(n803), .B1(ram[2826]), .B2(n804), .ZN(
        n7067) );
  MOAI22 U15997 ( .A1(n28410), .A2(n803), .B1(ram[2827]), .B2(n804), .ZN(
        n7068) );
  MOAI22 U15998 ( .A1(n28175), .A2(n803), .B1(ram[2828]), .B2(n804), .ZN(
        n7069) );
  MOAI22 U15999 ( .A1(n27940), .A2(n803), .B1(ram[2829]), .B2(n804), .ZN(
        n7070) );
  MOAI22 U16000 ( .A1(n27705), .A2(n803), .B1(ram[2830]), .B2(n804), .ZN(
        n7071) );
  MOAI22 U16001 ( .A1(n27470), .A2(n803), .B1(ram[2831]), .B2(n804), .ZN(
        n7072) );
  MOAI22 U16002 ( .A1(n29115), .A2(n805), .B1(ram[2832]), .B2(n806), .ZN(
        n7073) );
  MOAI22 U16003 ( .A1(n28880), .A2(n805), .B1(ram[2833]), .B2(n806), .ZN(
        n7074) );
  MOAI22 U16004 ( .A1(n28645), .A2(n805), .B1(ram[2834]), .B2(n806), .ZN(
        n7075) );
  MOAI22 U16005 ( .A1(n28410), .A2(n805), .B1(ram[2835]), .B2(n806), .ZN(
        n7076) );
  MOAI22 U16006 ( .A1(n28175), .A2(n805), .B1(ram[2836]), .B2(n806), .ZN(
        n7077) );
  MOAI22 U16007 ( .A1(n27940), .A2(n805), .B1(ram[2837]), .B2(n806), .ZN(
        n7078) );
  MOAI22 U16008 ( .A1(n27705), .A2(n805), .B1(ram[2838]), .B2(n806), .ZN(
        n7079) );
  MOAI22 U16009 ( .A1(n27470), .A2(n805), .B1(ram[2839]), .B2(n806), .ZN(
        n7080) );
  MOAI22 U16010 ( .A1(n29115), .A2(n807), .B1(ram[2840]), .B2(n808), .ZN(
        n7081) );
  MOAI22 U16011 ( .A1(n28880), .A2(n807), .B1(ram[2841]), .B2(n808), .ZN(
        n7082) );
  MOAI22 U16012 ( .A1(n28645), .A2(n807), .B1(ram[2842]), .B2(n808), .ZN(
        n7083) );
  MOAI22 U16013 ( .A1(n28410), .A2(n807), .B1(ram[2843]), .B2(n808), .ZN(
        n7084) );
  MOAI22 U16014 ( .A1(n28175), .A2(n807), .B1(ram[2844]), .B2(n808), .ZN(
        n7085) );
  MOAI22 U16015 ( .A1(n27940), .A2(n807), .B1(ram[2845]), .B2(n808), .ZN(
        n7086) );
  MOAI22 U16016 ( .A1(n27705), .A2(n807), .B1(ram[2846]), .B2(n808), .ZN(
        n7087) );
  MOAI22 U16017 ( .A1(n27470), .A2(n807), .B1(ram[2847]), .B2(n808), .ZN(
        n7088) );
  MOAI22 U16018 ( .A1(n29115), .A2(n809), .B1(ram[2848]), .B2(n810), .ZN(
        n7089) );
  MOAI22 U16019 ( .A1(n28880), .A2(n809), .B1(ram[2849]), .B2(n810), .ZN(
        n7090) );
  MOAI22 U16020 ( .A1(n28645), .A2(n809), .B1(ram[2850]), .B2(n810), .ZN(
        n7091) );
  MOAI22 U16021 ( .A1(n28410), .A2(n809), .B1(ram[2851]), .B2(n810), .ZN(
        n7092) );
  MOAI22 U16022 ( .A1(n28175), .A2(n809), .B1(ram[2852]), .B2(n810), .ZN(
        n7093) );
  MOAI22 U16023 ( .A1(n27940), .A2(n809), .B1(ram[2853]), .B2(n810), .ZN(
        n7094) );
  MOAI22 U16024 ( .A1(n27705), .A2(n809), .B1(ram[2854]), .B2(n810), .ZN(
        n7095) );
  MOAI22 U16025 ( .A1(n27470), .A2(n809), .B1(ram[2855]), .B2(n810), .ZN(
        n7096) );
  MOAI22 U16026 ( .A1(n29115), .A2(n811), .B1(ram[2856]), .B2(n812), .ZN(
        n7097) );
  MOAI22 U16027 ( .A1(n28880), .A2(n811), .B1(ram[2857]), .B2(n812), .ZN(
        n7098) );
  MOAI22 U16028 ( .A1(n28645), .A2(n811), .B1(ram[2858]), .B2(n812), .ZN(
        n7099) );
  MOAI22 U16029 ( .A1(n28410), .A2(n811), .B1(ram[2859]), .B2(n812), .ZN(
        n7100) );
  MOAI22 U16030 ( .A1(n28175), .A2(n811), .B1(ram[2860]), .B2(n812), .ZN(
        n7101) );
  MOAI22 U16031 ( .A1(n27940), .A2(n811), .B1(ram[2861]), .B2(n812), .ZN(
        n7102) );
  MOAI22 U16032 ( .A1(n27705), .A2(n811), .B1(ram[2862]), .B2(n812), .ZN(
        n7103) );
  MOAI22 U16033 ( .A1(n27470), .A2(n811), .B1(ram[2863]), .B2(n812), .ZN(
        n7104) );
  MOAI22 U16034 ( .A1(n29115), .A2(n813), .B1(ram[2864]), .B2(n814), .ZN(
        n7105) );
  MOAI22 U16035 ( .A1(n28880), .A2(n813), .B1(ram[2865]), .B2(n814), .ZN(
        n7106) );
  MOAI22 U16036 ( .A1(n28645), .A2(n813), .B1(ram[2866]), .B2(n814), .ZN(
        n7107) );
  MOAI22 U16037 ( .A1(n28410), .A2(n813), .B1(ram[2867]), .B2(n814), .ZN(
        n7108) );
  MOAI22 U16038 ( .A1(n28175), .A2(n813), .B1(ram[2868]), .B2(n814), .ZN(
        n7109) );
  MOAI22 U16039 ( .A1(n27940), .A2(n813), .B1(ram[2869]), .B2(n814), .ZN(
        n7110) );
  MOAI22 U16040 ( .A1(n27705), .A2(n813), .B1(ram[2870]), .B2(n814), .ZN(
        n7111) );
  MOAI22 U16041 ( .A1(n27470), .A2(n813), .B1(ram[2871]), .B2(n814), .ZN(
        n7112) );
  MOAI22 U16042 ( .A1(n29115), .A2(n815), .B1(ram[2872]), .B2(n816), .ZN(
        n7113) );
  MOAI22 U16043 ( .A1(n28880), .A2(n815), .B1(ram[2873]), .B2(n816), .ZN(
        n7114) );
  MOAI22 U16044 ( .A1(n28645), .A2(n815), .B1(ram[2874]), .B2(n816), .ZN(
        n7115) );
  MOAI22 U16045 ( .A1(n28410), .A2(n815), .B1(ram[2875]), .B2(n816), .ZN(
        n7116) );
  MOAI22 U16046 ( .A1(n28175), .A2(n815), .B1(ram[2876]), .B2(n816), .ZN(
        n7117) );
  MOAI22 U16047 ( .A1(n27940), .A2(n815), .B1(ram[2877]), .B2(n816), .ZN(
        n7118) );
  MOAI22 U16048 ( .A1(n27705), .A2(n815), .B1(ram[2878]), .B2(n816), .ZN(
        n7119) );
  MOAI22 U16049 ( .A1(n27470), .A2(n815), .B1(ram[2879]), .B2(n816), .ZN(
        n7120) );
  MOAI22 U16050 ( .A1(n29115), .A2(n817), .B1(ram[2880]), .B2(n818), .ZN(
        n7121) );
  MOAI22 U16051 ( .A1(n28880), .A2(n817), .B1(ram[2881]), .B2(n818), .ZN(
        n7122) );
  MOAI22 U16052 ( .A1(n28645), .A2(n817), .B1(ram[2882]), .B2(n818), .ZN(
        n7123) );
  MOAI22 U16053 ( .A1(n28410), .A2(n817), .B1(ram[2883]), .B2(n818), .ZN(
        n7124) );
  MOAI22 U16054 ( .A1(n28175), .A2(n817), .B1(ram[2884]), .B2(n818), .ZN(
        n7125) );
  MOAI22 U16055 ( .A1(n27940), .A2(n817), .B1(ram[2885]), .B2(n818), .ZN(
        n7126) );
  MOAI22 U16056 ( .A1(n27705), .A2(n817), .B1(ram[2886]), .B2(n818), .ZN(
        n7127) );
  MOAI22 U16057 ( .A1(n27470), .A2(n817), .B1(ram[2887]), .B2(n818), .ZN(
        n7128) );
  MOAI22 U16058 ( .A1(n29115), .A2(n819), .B1(ram[2888]), .B2(n820), .ZN(
        n7129) );
  MOAI22 U16059 ( .A1(n28880), .A2(n819), .B1(ram[2889]), .B2(n820), .ZN(
        n7130) );
  MOAI22 U16060 ( .A1(n28645), .A2(n819), .B1(ram[2890]), .B2(n820), .ZN(
        n7131) );
  MOAI22 U16061 ( .A1(n28410), .A2(n819), .B1(ram[2891]), .B2(n820), .ZN(
        n7132) );
  MOAI22 U16062 ( .A1(n28175), .A2(n819), .B1(ram[2892]), .B2(n820), .ZN(
        n7133) );
  MOAI22 U16063 ( .A1(n27940), .A2(n819), .B1(ram[2893]), .B2(n820), .ZN(
        n7134) );
  MOAI22 U16064 ( .A1(n27705), .A2(n819), .B1(ram[2894]), .B2(n820), .ZN(
        n7135) );
  MOAI22 U16065 ( .A1(n27470), .A2(n819), .B1(ram[2895]), .B2(n820), .ZN(
        n7136) );
  MOAI22 U16066 ( .A1(n29115), .A2(n821), .B1(ram[2896]), .B2(n822), .ZN(
        n7137) );
  MOAI22 U16067 ( .A1(n28880), .A2(n821), .B1(ram[2897]), .B2(n822), .ZN(
        n7138) );
  MOAI22 U16068 ( .A1(n28645), .A2(n821), .B1(ram[2898]), .B2(n822), .ZN(
        n7139) );
  MOAI22 U16069 ( .A1(n28410), .A2(n821), .B1(ram[2899]), .B2(n822), .ZN(
        n7140) );
  MOAI22 U16070 ( .A1(n28175), .A2(n821), .B1(ram[2900]), .B2(n822), .ZN(
        n7141) );
  MOAI22 U16071 ( .A1(n27940), .A2(n821), .B1(ram[2901]), .B2(n822), .ZN(
        n7142) );
  MOAI22 U16072 ( .A1(n27705), .A2(n821), .B1(ram[2902]), .B2(n822), .ZN(
        n7143) );
  MOAI22 U16073 ( .A1(n27470), .A2(n821), .B1(ram[2903]), .B2(n822), .ZN(
        n7144) );
  MOAI22 U16074 ( .A1(n29115), .A2(n823), .B1(ram[2904]), .B2(n824), .ZN(
        n7145) );
  MOAI22 U16075 ( .A1(n28880), .A2(n823), .B1(ram[2905]), .B2(n824), .ZN(
        n7146) );
  MOAI22 U16076 ( .A1(n28645), .A2(n823), .B1(ram[2906]), .B2(n824), .ZN(
        n7147) );
  MOAI22 U16077 ( .A1(n28410), .A2(n823), .B1(ram[2907]), .B2(n824), .ZN(
        n7148) );
  MOAI22 U16078 ( .A1(n28175), .A2(n823), .B1(ram[2908]), .B2(n824), .ZN(
        n7149) );
  MOAI22 U16079 ( .A1(n27940), .A2(n823), .B1(ram[2909]), .B2(n824), .ZN(
        n7150) );
  MOAI22 U16080 ( .A1(n27705), .A2(n823), .B1(ram[2910]), .B2(n824), .ZN(
        n7151) );
  MOAI22 U16081 ( .A1(n27470), .A2(n823), .B1(ram[2911]), .B2(n824), .ZN(
        n7152) );
  MOAI22 U16082 ( .A1(n29116), .A2(n825), .B1(ram[2912]), .B2(n826), .ZN(
        n7153) );
  MOAI22 U16083 ( .A1(n28881), .A2(n825), .B1(ram[2913]), .B2(n826), .ZN(
        n7154) );
  MOAI22 U16084 ( .A1(n28646), .A2(n825), .B1(ram[2914]), .B2(n826), .ZN(
        n7155) );
  MOAI22 U16085 ( .A1(n28411), .A2(n825), .B1(ram[2915]), .B2(n826), .ZN(
        n7156) );
  MOAI22 U16086 ( .A1(n28176), .A2(n825), .B1(ram[2916]), .B2(n826), .ZN(
        n7157) );
  MOAI22 U16087 ( .A1(n27941), .A2(n825), .B1(ram[2917]), .B2(n826), .ZN(
        n7158) );
  MOAI22 U16088 ( .A1(n27706), .A2(n825), .B1(ram[2918]), .B2(n826), .ZN(
        n7159) );
  MOAI22 U16089 ( .A1(n27471), .A2(n825), .B1(ram[2919]), .B2(n826), .ZN(
        n7160) );
  MOAI22 U16090 ( .A1(n29116), .A2(n827), .B1(ram[2920]), .B2(n828), .ZN(
        n7161) );
  MOAI22 U16091 ( .A1(n28881), .A2(n827), .B1(ram[2921]), .B2(n828), .ZN(
        n7162) );
  MOAI22 U16092 ( .A1(n28646), .A2(n827), .B1(ram[2922]), .B2(n828), .ZN(
        n7163) );
  MOAI22 U16093 ( .A1(n28411), .A2(n827), .B1(ram[2923]), .B2(n828), .ZN(
        n7164) );
  MOAI22 U16094 ( .A1(n28176), .A2(n827), .B1(ram[2924]), .B2(n828), .ZN(
        n7165) );
  MOAI22 U16095 ( .A1(n27941), .A2(n827), .B1(ram[2925]), .B2(n828), .ZN(
        n7166) );
  MOAI22 U16096 ( .A1(n27706), .A2(n827), .B1(ram[2926]), .B2(n828), .ZN(
        n7167) );
  MOAI22 U16097 ( .A1(n27471), .A2(n827), .B1(ram[2927]), .B2(n828), .ZN(
        n7168) );
  MOAI22 U16098 ( .A1(n29116), .A2(n829), .B1(ram[2928]), .B2(n830), .ZN(
        n7169) );
  MOAI22 U16099 ( .A1(n28881), .A2(n829), .B1(ram[2929]), .B2(n830), .ZN(
        n7170) );
  MOAI22 U16100 ( .A1(n28646), .A2(n829), .B1(ram[2930]), .B2(n830), .ZN(
        n7171) );
  MOAI22 U16101 ( .A1(n28411), .A2(n829), .B1(ram[2931]), .B2(n830), .ZN(
        n7172) );
  MOAI22 U16102 ( .A1(n28176), .A2(n829), .B1(ram[2932]), .B2(n830), .ZN(
        n7173) );
  MOAI22 U16103 ( .A1(n27941), .A2(n829), .B1(ram[2933]), .B2(n830), .ZN(
        n7174) );
  MOAI22 U16104 ( .A1(n27706), .A2(n829), .B1(ram[2934]), .B2(n830), .ZN(
        n7175) );
  MOAI22 U16105 ( .A1(n27471), .A2(n829), .B1(ram[2935]), .B2(n830), .ZN(
        n7176) );
  MOAI22 U16106 ( .A1(n29116), .A2(n831), .B1(ram[2936]), .B2(n832), .ZN(
        n7177) );
  MOAI22 U16107 ( .A1(n28881), .A2(n831), .B1(ram[2937]), .B2(n832), .ZN(
        n7178) );
  MOAI22 U16108 ( .A1(n28646), .A2(n831), .B1(ram[2938]), .B2(n832), .ZN(
        n7179) );
  MOAI22 U16109 ( .A1(n28411), .A2(n831), .B1(ram[2939]), .B2(n832), .ZN(
        n7180) );
  MOAI22 U16110 ( .A1(n28176), .A2(n831), .B1(ram[2940]), .B2(n832), .ZN(
        n7181) );
  MOAI22 U16111 ( .A1(n27941), .A2(n831), .B1(ram[2941]), .B2(n832), .ZN(
        n7182) );
  MOAI22 U16112 ( .A1(n27706), .A2(n831), .B1(ram[2942]), .B2(n832), .ZN(
        n7183) );
  MOAI22 U16113 ( .A1(n27471), .A2(n831), .B1(ram[2943]), .B2(n832), .ZN(
        n7184) );
  MOAI22 U16114 ( .A1(n29116), .A2(n833), .B1(ram[2944]), .B2(n834), .ZN(
        n7185) );
  MOAI22 U16115 ( .A1(n28881), .A2(n833), .B1(ram[2945]), .B2(n834), .ZN(
        n7186) );
  MOAI22 U16116 ( .A1(n28646), .A2(n833), .B1(ram[2946]), .B2(n834), .ZN(
        n7187) );
  MOAI22 U16117 ( .A1(n28411), .A2(n833), .B1(ram[2947]), .B2(n834), .ZN(
        n7188) );
  MOAI22 U16118 ( .A1(n28176), .A2(n833), .B1(ram[2948]), .B2(n834), .ZN(
        n7189) );
  MOAI22 U16119 ( .A1(n27941), .A2(n833), .B1(ram[2949]), .B2(n834), .ZN(
        n7190) );
  MOAI22 U16120 ( .A1(n27706), .A2(n833), .B1(ram[2950]), .B2(n834), .ZN(
        n7191) );
  MOAI22 U16121 ( .A1(n27471), .A2(n833), .B1(ram[2951]), .B2(n834), .ZN(
        n7192) );
  MOAI22 U16122 ( .A1(n29116), .A2(n835), .B1(ram[2952]), .B2(n836), .ZN(
        n7193) );
  MOAI22 U16123 ( .A1(n28881), .A2(n835), .B1(ram[2953]), .B2(n836), .ZN(
        n7194) );
  MOAI22 U16124 ( .A1(n28646), .A2(n835), .B1(ram[2954]), .B2(n836), .ZN(
        n7195) );
  MOAI22 U16125 ( .A1(n28411), .A2(n835), .B1(ram[2955]), .B2(n836), .ZN(
        n7196) );
  MOAI22 U16126 ( .A1(n28176), .A2(n835), .B1(ram[2956]), .B2(n836), .ZN(
        n7197) );
  MOAI22 U16127 ( .A1(n27941), .A2(n835), .B1(ram[2957]), .B2(n836), .ZN(
        n7198) );
  MOAI22 U16128 ( .A1(n27706), .A2(n835), .B1(ram[2958]), .B2(n836), .ZN(
        n7199) );
  MOAI22 U16129 ( .A1(n27471), .A2(n835), .B1(ram[2959]), .B2(n836), .ZN(
        n7200) );
  MOAI22 U16130 ( .A1(n29116), .A2(n837), .B1(ram[2960]), .B2(n838), .ZN(
        n7201) );
  MOAI22 U16131 ( .A1(n28881), .A2(n837), .B1(ram[2961]), .B2(n838), .ZN(
        n7202) );
  MOAI22 U16132 ( .A1(n28646), .A2(n837), .B1(ram[2962]), .B2(n838), .ZN(
        n7203) );
  MOAI22 U16133 ( .A1(n28411), .A2(n837), .B1(ram[2963]), .B2(n838), .ZN(
        n7204) );
  MOAI22 U16134 ( .A1(n28176), .A2(n837), .B1(ram[2964]), .B2(n838), .ZN(
        n7205) );
  MOAI22 U16135 ( .A1(n27941), .A2(n837), .B1(ram[2965]), .B2(n838), .ZN(
        n7206) );
  MOAI22 U16136 ( .A1(n27706), .A2(n837), .B1(ram[2966]), .B2(n838), .ZN(
        n7207) );
  MOAI22 U16137 ( .A1(n27471), .A2(n837), .B1(ram[2967]), .B2(n838), .ZN(
        n7208) );
  MOAI22 U16138 ( .A1(n29116), .A2(n839), .B1(ram[2968]), .B2(n840), .ZN(
        n7209) );
  MOAI22 U16139 ( .A1(n28881), .A2(n839), .B1(ram[2969]), .B2(n840), .ZN(
        n7210) );
  MOAI22 U16140 ( .A1(n28646), .A2(n839), .B1(ram[2970]), .B2(n840), .ZN(
        n7211) );
  MOAI22 U16141 ( .A1(n28411), .A2(n839), .B1(ram[2971]), .B2(n840), .ZN(
        n7212) );
  MOAI22 U16142 ( .A1(n28176), .A2(n839), .B1(ram[2972]), .B2(n840), .ZN(
        n7213) );
  MOAI22 U16143 ( .A1(n27941), .A2(n839), .B1(ram[2973]), .B2(n840), .ZN(
        n7214) );
  MOAI22 U16144 ( .A1(n27706), .A2(n839), .B1(ram[2974]), .B2(n840), .ZN(
        n7215) );
  MOAI22 U16145 ( .A1(n27471), .A2(n839), .B1(ram[2975]), .B2(n840), .ZN(
        n7216) );
  MOAI22 U16146 ( .A1(n29116), .A2(n841), .B1(ram[2976]), .B2(n842), .ZN(
        n7217) );
  MOAI22 U16147 ( .A1(n28881), .A2(n841), .B1(ram[2977]), .B2(n842), .ZN(
        n7218) );
  MOAI22 U16148 ( .A1(n28646), .A2(n841), .B1(ram[2978]), .B2(n842), .ZN(
        n7219) );
  MOAI22 U16149 ( .A1(n28411), .A2(n841), .B1(ram[2979]), .B2(n842), .ZN(
        n7220) );
  MOAI22 U16150 ( .A1(n28176), .A2(n841), .B1(ram[2980]), .B2(n842), .ZN(
        n7221) );
  MOAI22 U16151 ( .A1(n27941), .A2(n841), .B1(ram[2981]), .B2(n842), .ZN(
        n7222) );
  MOAI22 U16152 ( .A1(n27706), .A2(n841), .B1(ram[2982]), .B2(n842), .ZN(
        n7223) );
  MOAI22 U16153 ( .A1(n27471), .A2(n841), .B1(ram[2983]), .B2(n842), .ZN(
        n7224) );
  MOAI22 U16154 ( .A1(n29116), .A2(n843), .B1(ram[2984]), .B2(n844), .ZN(
        n7225) );
  MOAI22 U16155 ( .A1(n28881), .A2(n843), .B1(ram[2985]), .B2(n844), .ZN(
        n7226) );
  MOAI22 U16156 ( .A1(n28646), .A2(n843), .B1(ram[2986]), .B2(n844), .ZN(
        n7227) );
  MOAI22 U16157 ( .A1(n28411), .A2(n843), .B1(ram[2987]), .B2(n844), .ZN(
        n7228) );
  MOAI22 U16158 ( .A1(n28176), .A2(n843), .B1(ram[2988]), .B2(n844), .ZN(
        n7229) );
  MOAI22 U16159 ( .A1(n27941), .A2(n843), .B1(ram[2989]), .B2(n844), .ZN(
        n7230) );
  MOAI22 U16160 ( .A1(n27706), .A2(n843), .B1(ram[2990]), .B2(n844), .ZN(
        n7231) );
  MOAI22 U16161 ( .A1(n27471), .A2(n843), .B1(ram[2991]), .B2(n844), .ZN(
        n7232) );
  MOAI22 U16162 ( .A1(n29116), .A2(n845), .B1(ram[2992]), .B2(n846), .ZN(
        n7233) );
  MOAI22 U16163 ( .A1(n28881), .A2(n845), .B1(ram[2993]), .B2(n846), .ZN(
        n7234) );
  MOAI22 U16164 ( .A1(n28646), .A2(n845), .B1(ram[2994]), .B2(n846), .ZN(
        n7235) );
  MOAI22 U16165 ( .A1(n28411), .A2(n845), .B1(ram[2995]), .B2(n846), .ZN(
        n7236) );
  MOAI22 U16166 ( .A1(n28176), .A2(n845), .B1(ram[2996]), .B2(n846), .ZN(
        n7237) );
  MOAI22 U16167 ( .A1(n27941), .A2(n845), .B1(ram[2997]), .B2(n846), .ZN(
        n7238) );
  MOAI22 U16168 ( .A1(n27706), .A2(n845), .B1(ram[2998]), .B2(n846), .ZN(
        n7239) );
  MOAI22 U16169 ( .A1(n27471), .A2(n845), .B1(ram[2999]), .B2(n846), .ZN(
        n7240) );
  MOAI22 U16170 ( .A1(n29116), .A2(n847), .B1(ram[3000]), .B2(n848), .ZN(
        n7241) );
  MOAI22 U16171 ( .A1(n28881), .A2(n847), .B1(ram[3001]), .B2(n848), .ZN(
        n7242) );
  MOAI22 U16172 ( .A1(n28646), .A2(n847), .B1(ram[3002]), .B2(n848), .ZN(
        n7243) );
  MOAI22 U16173 ( .A1(n28411), .A2(n847), .B1(ram[3003]), .B2(n848), .ZN(
        n7244) );
  MOAI22 U16174 ( .A1(n28176), .A2(n847), .B1(ram[3004]), .B2(n848), .ZN(
        n7245) );
  MOAI22 U16175 ( .A1(n27941), .A2(n847), .B1(ram[3005]), .B2(n848), .ZN(
        n7246) );
  MOAI22 U16176 ( .A1(n27706), .A2(n847), .B1(ram[3006]), .B2(n848), .ZN(
        n7247) );
  MOAI22 U16177 ( .A1(n27471), .A2(n847), .B1(ram[3007]), .B2(n848), .ZN(
        n7248) );
  MOAI22 U16178 ( .A1(n29116), .A2(n849), .B1(ram[3008]), .B2(n850), .ZN(
        n7249) );
  MOAI22 U16179 ( .A1(n28881), .A2(n849), .B1(ram[3009]), .B2(n850), .ZN(
        n7250) );
  MOAI22 U16180 ( .A1(n28646), .A2(n849), .B1(ram[3010]), .B2(n850), .ZN(
        n7251) );
  MOAI22 U16181 ( .A1(n28411), .A2(n849), .B1(ram[3011]), .B2(n850), .ZN(
        n7252) );
  MOAI22 U16182 ( .A1(n28176), .A2(n849), .B1(ram[3012]), .B2(n850), .ZN(
        n7253) );
  MOAI22 U16183 ( .A1(n27941), .A2(n849), .B1(ram[3013]), .B2(n850), .ZN(
        n7254) );
  MOAI22 U16184 ( .A1(n27706), .A2(n849), .B1(ram[3014]), .B2(n850), .ZN(
        n7255) );
  MOAI22 U16185 ( .A1(n27471), .A2(n849), .B1(ram[3015]), .B2(n850), .ZN(
        n7256) );
  MOAI22 U16186 ( .A1(n29117), .A2(n851), .B1(ram[3016]), .B2(n852), .ZN(
        n7257) );
  MOAI22 U16187 ( .A1(n28882), .A2(n851), .B1(ram[3017]), .B2(n852), .ZN(
        n7258) );
  MOAI22 U16188 ( .A1(n28647), .A2(n851), .B1(ram[3018]), .B2(n852), .ZN(
        n7259) );
  MOAI22 U16189 ( .A1(n28412), .A2(n851), .B1(ram[3019]), .B2(n852), .ZN(
        n7260) );
  MOAI22 U16190 ( .A1(n28177), .A2(n851), .B1(ram[3020]), .B2(n852), .ZN(
        n7261) );
  MOAI22 U16191 ( .A1(n27942), .A2(n851), .B1(ram[3021]), .B2(n852), .ZN(
        n7262) );
  MOAI22 U16192 ( .A1(n27707), .A2(n851), .B1(ram[3022]), .B2(n852), .ZN(
        n7263) );
  MOAI22 U16193 ( .A1(n27472), .A2(n851), .B1(ram[3023]), .B2(n852), .ZN(
        n7264) );
  MOAI22 U16194 ( .A1(n29117), .A2(n853), .B1(ram[3024]), .B2(n854), .ZN(
        n7265) );
  MOAI22 U16195 ( .A1(n28882), .A2(n853), .B1(ram[3025]), .B2(n854), .ZN(
        n7266) );
  MOAI22 U16196 ( .A1(n28647), .A2(n853), .B1(ram[3026]), .B2(n854), .ZN(
        n7267) );
  MOAI22 U16197 ( .A1(n28412), .A2(n853), .B1(ram[3027]), .B2(n854), .ZN(
        n7268) );
  MOAI22 U16198 ( .A1(n28177), .A2(n853), .B1(ram[3028]), .B2(n854), .ZN(
        n7269) );
  MOAI22 U16199 ( .A1(n27942), .A2(n853), .B1(ram[3029]), .B2(n854), .ZN(
        n7270) );
  MOAI22 U16200 ( .A1(n27707), .A2(n853), .B1(ram[3030]), .B2(n854), .ZN(
        n7271) );
  MOAI22 U16201 ( .A1(n27472), .A2(n853), .B1(ram[3031]), .B2(n854), .ZN(
        n7272) );
  MOAI22 U16202 ( .A1(n29117), .A2(n855), .B1(ram[3032]), .B2(n856), .ZN(
        n7273) );
  MOAI22 U16203 ( .A1(n28882), .A2(n855), .B1(ram[3033]), .B2(n856), .ZN(
        n7274) );
  MOAI22 U16204 ( .A1(n28647), .A2(n855), .B1(ram[3034]), .B2(n856), .ZN(
        n7275) );
  MOAI22 U16205 ( .A1(n28412), .A2(n855), .B1(ram[3035]), .B2(n856), .ZN(
        n7276) );
  MOAI22 U16206 ( .A1(n28177), .A2(n855), .B1(ram[3036]), .B2(n856), .ZN(
        n7277) );
  MOAI22 U16207 ( .A1(n27942), .A2(n855), .B1(ram[3037]), .B2(n856), .ZN(
        n7278) );
  MOAI22 U16208 ( .A1(n27707), .A2(n855), .B1(ram[3038]), .B2(n856), .ZN(
        n7279) );
  MOAI22 U16209 ( .A1(n27472), .A2(n855), .B1(ram[3039]), .B2(n856), .ZN(
        n7280) );
  MOAI22 U16210 ( .A1(n29117), .A2(n857), .B1(ram[3040]), .B2(n858), .ZN(
        n7281) );
  MOAI22 U16211 ( .A1(n28882), .A2(n857), .B1(ram[3041]), .B2(n858), .ZN(
        n7282) );
  MOAI22 U16212 ( .A1(n28647), .A2(n857), .B1(ram[3042]), .B2(n858), .ZN(
        n7283) );
  MOAI22 U16213 ( .A1(n28412), .A2(n857), .B1(ram[3043]), .B2(n858), .ZN(
        n7284) );
  MOAI22 U16214 ( .A1(n28177), .A2(n857), .B1(ram[3044]), .B2(n858), .ZN(
        n7285) );
  MOAI22 U16215 ( .A1(n27942), .A2(n857), .B1(ram[3045]), .B2(n858), .ZN(
        n7286) );
  MOAI22 U16216 ( .A1(n27707), .A2(n857), .B1(ram[3046]), .B2(n858), .ZN(
        n7287) );
  MOAI22 U16217 ( .A1(n27472), .A2(n857), .B1(ram[3047]), .B2(n858), .ZN(
        n7288) );
  MOAI22 U16218 ( .A1(n29117), .A2(n859), .B1(ram[3048]), .B2(n860), .ZN(
        n7289) );
  MOAI22 U16219 ( .A1(n28882), .A2(n859), .B1(ram[3049]), .B2(n860), .ZN(
        n7290) );
  MOAI22 U16220 ( .A1(n28647), .A2(n859), .B1(ram[3050]), .B2(n860), .ZN(
        n7291) );
  MOAI22 U16221 ( .A1(n28412), .A2(n859), .B1(ram[3051]), .B2(n860), .ZN(
        n7292) );
  MOAI22 U16222 ( .A1(n28177), .A2(n859), .B1(ram[3052]), .B2(n860), .ZN(
        n7293) );
  MOAI22 U16223 ( .A1(n27942), .A2(n859), .B1(ram[3053]), .B2(n860), .ZN(
        n7294) );
  MOAI22 U16224 ( .A1(n27707), .A2(n859), .B1(ram[3054]), .B2(n860), .ZN(
        n7295) );
  MOAI22 U16225 ( .A1(n27472), .A2(n859), .B1(ram[3055]), .B2(n860), .ZN(
        n7296) );
  MOAI22 U16226 ( .A1(n29117), .A2(n861), .B1(ram[3056]), .B2(n862), .ZN(
        n7297) );
  MOAI22 U16227 ( .A1(n28882), .A2(n861), .B1(ram[3057]), .B2(n862), .ZN(
        n7298) );
  MOAI22 U16228 ( .A1(n28647), .A2(n861), .B1(ram[3058]), .B2(n862), .ZN(
        n7299) );
  MOAI22 U16229 ( .A1(n28412), .A2(n861), .B1(ram[3059]), .B2(n862), .ZN(
        n7300) );
  MOAI22 U16230 ( .A1(n28177), .A2(n861), .B1(ram[3060]), .B2(n862), .ZN(
        n7301) );
  MOAI22 U16231 ( .A1(n27942), .A2(n861), .B1(ram[3061]), .B2(n862), .ZN(
        n7302) );
  MOAI22 U16232 ( .A1(n27707), .A2(n861), .B1(ram[3062]), .B2(n862), .ZN(
        n7303) );
  MOAI22 U16233 ( .A1(n27472), .A2(n861), .B1(ram[3063]), .B2(n862), .ZN(
        n7304) );
  MOAI22 U16234 ( .A1(n29117), .A2(n863), .B1(ram[3064]), .B2(n864), .ZN(
        n7305) );
  MOAI22 U16235 ( .A1(n28882), .A2(n863), .B1(ram[3065]), .B2(n864), .ZN(
        n7306) );
  MOAI22 U16236 ( .A1(n28647), .A2(n863), .B1(ram[3066]), .B2(n864), .ZN(
        n7307) );
  MOAI22 U16237 ( .A1(n28412), .A2(n863), .B1(ram[3067]), .B2(n864), .ZN(
        n7308) );
  MOAI22 U16238 ( .A1(n28177), .A2(n863), .B1(ram[3068]), .B2(n864), .ZN(
        n7309) );
  MOAI22 U16239 ( .A1(n27942), .A2(n863), .B1(ram[3069]), .B2(n864), .ZN(
        n7310) );
  MOAI22 U16240 ( .A1(n27707), .A2(n863), .B1(ram[3070]), .B2(n864), .ZN(
        n7311) );
  MOAI22 U16241 ( .A1(n27472), .A2(n863), .B1(ram[3071]), .B2(n864), .ZN(
        n7312) );
  MOAI22 U16242 ( .A1(n29117), .A2(n866), .B1(ram[3072]), .B2(n867), .ZN(
        n7313) );
  MOAI22 U16243 ( .A1(n28882), .A2(n866), .B1(ram[3073]), .B2(n867), .ZN(
        n7314) );
  MOAI22 U16244 ( .A1(n28647), .A2(n866), .B1(ram[3074]), .B2(n867), .ZN(
        n7315) );
  MOAI22 U16245 ( .A1(n28412), .A2(n866), .B1(ram[3075]), .B2(n867), .ZN(
        n7316) );
  MOAI22 U16246 ( .A1(n28177), .A2(n866), .B1(ram[3076]), .B2(n867), .ZN(
        n7317) );
  MOAI22 U16247 ( .A1(n27942), .A2(n866), .B1(ram[3077]), .B2(n867), .ZN(
        n7318) );
  MOAI22 U16248 ( .A1(n27707), .A2(n866), .B1(ram[3078]), .B2(n867), .ZN(
        n7319) );
  MOAI22 U16249 ( .A1(n27472), .A2(n866), .B1(ram[3079]), .B2(n867), .ZN(
        n7320) );
  MOAI22 U16250 ( .A1(n29117), .A2(n869), .B1(ram[3080]), .B2(n870), .ZN(
        n7321) );
  MOAI22 U16251 ( .A1(n28882), .A2(n869), .B1(ram[3081]), .B2(n870), .ZN(
        n7322) );
  MOAI22 U16252 ( .A1(n28647), .A2(n869), .B1(ram[3082]), .B2(n870), .ZN(
        n7323) );
  MOAI22 U16253 ( .A1(n28412), .A2(n869), .B1(ram[3083]), .B2(n870), .ZN(
        n7324) );
  MOAI22 U16254 ( .A1(n28177), .A2(n869), .B1(ram[3084]), .B2(n870), .ZN(
        n7325) );
  MOAI22 U16255 ( .A1(n27942), .A2(n869), .B1(ram[3085]), .B2(n870), .ZN(
        n7326) );
  MOAI22 U16256 ( .A1(n27707), .A2(n869), .B1(ram[3086]), .B2(n870), .ZN(
        n7327) );
  MOAI22 U16257 ( .A1(n27472), .A2(n869), .B1(ram[3087]), .B2(n870), .ZN(
        n7328) );
  MOAI22 U16258 ( .A1(n29117), .A2(n871), .B1(ram[3088]), .B2(n872), .ZN(
        n7329) );
  MOAI22 U16259 ( .A1(n28882), .A2(n871), .B1(ram[3089]), .B2(n872), .ZN(
        n7330) );
  MOAI22 U16260 ( .A1(n28647), .A2(n871), .B1(ram[3090]), .B2(n872), .ZN(
        n7331) );
  MOAI22 U16261 ( .A1(n28412), .A2(n871), .B1(ram[3091]), .B2(n872), .ZN(
        n7332) );
  MOAI22 U16262 ( .A1(n28177), .A2(n871), .B1(ram[3092]), .B2(n872), .ZN(
        n7333) );
  MOAI22 U16263 ( .A1(n27942), .A2(n871), .B1(ram[3093]), .B2(n872), .ZN(
        n7334) );
  MOAI22 U16264 ( .A1(n27707), .A2(n871), .B1(ram[3094]), .B2(n872), .ZN(
        n7335) );
  MOAI22 U16265 ( .A1(n27472), .A2(n871), .B1(ram[3095]), .B2(n872), .ZN(
        n7336) );
  MOAI22 U16266 ( .A1(n29117), .A2(n873), .B1(ram[3096]), .B2(n874), .ZN(
        n7337) );
  MOAI22 U16267 ( .A1(n28882), .A2(n873), .B1(ram[3097]), .B2(n874), .ZN(
        n7338) );
  MOAI22 U16268 ( .A1(n28647), .A2(n873), .B1(ram[3098]), .B2(n874), .ZN(
        n7339) );
  MOAI22 U16269 ( .A1(n28412), .A2(n873), .B1(ram[3099]), .B2(n874), .ZN(
        n7340) );
  MOAI22 U16270 ( .A1(n28177), .A2(n873), .B1(ram[3100]), .B2(n874), .ZN(
        n7341) );
  MOAI22 U16271 ( .A1(n27942), .A2(n873), .B1(ram[3101]), .B2(n874), .ZN(
        n7342) );
  MOAI22 U16272 ( .A1(n27707), .A2(n873), .B1(ram[3102]), .B2(n874), .ZN(
        n7343) );
  MOAI22 U16273 ( .A1(n27472), .A2(n873), .B1(ram[3103]), .B2(n874), .ZN(
        n7344) );
  MOAI22 U16274 ( .A1(n29117), .A2(n875), .B1(ram[3104]), .B2(n876), .ZN(
        n7345) );
  MOAI22 U16275 ( .A1(n28882), .A2(n875), .B1(ram[3105]), .B2(n876), .ZN(
        n7346) );
  MOAI22 U16276 ( .A1(n28647), .A2(n875), .B1(ram[3106]), .B2(n876), .ZN(
        n7347) );
  MOAI22 U16277 ( .A1(n28412), .A2(n875), .B1(ram[3107]), .B2(n876), .ZN(
        n7348) );
  MOAI22 U16278 ( .A1(n28177), .A2(n875), .B1(ram[3108]), .B2(n876), .ZN(
        n7349) );
  MOAI22 U16279 ( .A1(n27942), .A2(n875), .B1(ram[3109]), .B2(n876), .ZN(
        n7350) );
  MOAI22 U16280 ( .A1(n27707), .A2(n875), .B1(ram[3110]), .B2(n876), .ZN(
        n7351) );
  MOAI22 U16281 ( .A1(n27472), .A2(n875), .B1(ram[3111]), .B2(n876), .ZN(
        n7352) );
  MOAI22 U16282 ( .A1(n29117), .A2(n877), .B1(ram[3112]), .B2(n878), .ZN(
        n7353) );
  MOAI22 U16283 ( .A1(n28882), .A2(n877), .B1(ram[3113]), .B2(n878), .ZN(
        n7354) );
  MOAI22 U16284 ( .A1(n28647), .A2(n877), .B1(ram[3114]), .B2(n878), .ZN(
        n7355) );
  MOAI22 U16285 ( .A1(n28412), .A2(n877), .B1(ram[3115]), .B2(n878), .ZN(
        n7356) );
  MOAI22 U16286 ( .A1(n28177), .A2(n877), .B1(ram[3116]), .B2(n878), .ZN(
        n7357) );
  MOAI22 U16287 ( .A1(n27942), .A2(n877), .B1(ram[3117]), .B2(n878), .ZN(
        n7358) );
  MOAI22 U16288 ( .A1(n27707), .A2(n877), .B1(ram[3118]), .B2(n878), .ZN(
        n7359) );
  MOAI22 U16289 ( .A1(n27472), .A2(n877), .B1(ram[3119]), .B2(n878), .ZN(
        n7360) );
  MOAI22 U16290 ( .A1(n29118), .A2(n879), .B1(ram[3120]), .B2(n880), .ZN(
        n7361) );
  MOAI22 U16291 ( .A1(n28883), .A2(n879), .B1(ram[3121]), .B2(n880), .ZN(
        n7362) );
  MOAI22 U16292 ( .A1(n28648), .A2(n879), .B1(ram[3122]), .B2(n880), .ZN(
        n7363) );
  MOAI22 U16293 ( .A1(n28413), .A2(n879), .B1(ram[3123]), .B2(n880), .ZN(
        n7364) );
  MOAI22 U16294 ( .A1(n28178), .A2(n879), .B1(ram[3124]), .B2(n880), .ZN(
        n7365) );
  MOAI22 U16295 ( .A1(n27943), .A2(n879), .B1(ram[3125]), .B2(n880), .ZN(
        n7366) );
  MOAI22 U16296 ( .A1(n27708), .A2(n879), .B1(ram[3126]), .B2(n880), .ZN(
        n7367) );
  MOAI22 U16297 ( .A1(n27473), .A2(n879), .B1(ram[3127]), .B2(n880), .ZN(
        n7368) );
  MOAI22 U16298 ( .A1(n29118), .A2(n881), .B1(ram[3128]), .B2(n882), .ZN(
        n7369) );
  MOAI22 U16299 ( .A1(n28883), .A2(n881), .B1(ram[3129]), .B2(n882), .ZN(
        n7370) );
  MOAI22 U16300 ( .A1(n28648), .A2(n881), .B1(ram[3130]), .B2(n882), .ZN(
        n7371) );
  MOAI22 U16301 ( .A1(n28413), .A2(n881), .B1(ram[3131]), .B2(n882), .ZN(
        n7372) );
  MOAI22 U16302 ( .A1(n28178), .A2(n881), .B1(ram[3132]), .B2(n882), .ZN(
        n7373) );
  MOAI22 U16303 ( .A1(n27943), .A2(n881), .B1(ram[3133]), .B2(n882), .ZN(
        n7374) );
  MOAI22 U16304 ( .A1(n27708), .A2(n881), .B1(ram[3134]), .B2(n882), .ZN(
        n7375) );
  MOAI22 U16305 ( .A1(n27473), .A2(n881), .B1(ram[3135]), .B2(n882), .ZN(
        n7376) );
  MOAI22 U16306 ( .A1(n29118), .A2(n883), .B1(ram[3136]), .B2(n884), .ZN(
        n7377) );
  MOAI22 U16307 ( .A1(n28883), .A2(n883), .B1(ram[3137]), .B2(n884), .ZN(
        n7378) );
  MOAI22 U16308 ( .A1(n28648), .A2(n883), .B1(ram[3138]), .B2(n884), .ZN(
        n7379) );
  MOAI22 U16309 ( .A1(n28413), .A2(n883), .B1(ram[3139]), .B2(n884), .ZN(
        n7380) );
  MOAI22 U16310 ( .A1(n28178), .A2(n883), .B1(ram[3140]), .B2(n884), .ZN(
        n7381) );
  MOAI22 U16311 ( .A1(n27943), .A2(n883), .B1(ram[3141]), .B2(n884), .ZN(
        n7382) );
  MOAI22 U16312 ( .A1(n27708), .A2(n883), .B1(ram[3142]), .B2(n884), .ZN(
        n7383) );
  MOAI22 U16313 ( .A1(n27473), .A2(n883), .B1(ram[3143]), .B2(n884), .ZN(
        n7384) );
  MOAI22 U16314 ( .A1(n29118), .A2(n885), .B1(ram[3144]), .B2(n886), .ZN(
        n7385) );
  MOAI22 U16315 ( .A1(n28883), .A2(n885), .B1(ram[3145]), .B2(n886), .ZN(
        n7386) );
  MOAI22 U16316 ( .A1(n28648), .A2(n885), .B1(ram[3146]), .B2(n886), .ZN(
        n7387) );
  MOAI22 U16317 ( .A1(n28413), .A2(n885), .B1(ram[3147]), .B2(n886), .ZN(
        n7388) );
  MOAI22 U16318 ( .A1(n28178), .A2(n885), .B1(ram[3148]), .B2(n886), .ZN(
        n7389) );
  MOAI22 U16319 ( .A1(n27943), .A2(n885), .B1(ram[3149]), .B2(n886), .ZN(
        n7390) );
  MOAI22 U16320 ( .A1(n27708), .A2(n885), .B1(ram[3150]), .B2(n886), .ZN(
        n7391) );
  MOAI22 U16321 ( .A1(n27473), .A2(n885), .B1(ram[3151]), .B2(n886), .ZN(
        n7392) );
  MOAI22 U16322 ( .A1(n29118), .A2(n887), .B1(ram[3152]), .B2(n888), .ZN(
        n7393) );
  MOAI22 U16323 ( .A1(n28883), .A2(n887), .B1(ram[3153]), .B2(n888), .ZN(
        n7394) );
  MOAI22 U16324 ( .A1(n28648), .A2(n887), .B1(ram[3154]), .B2(n888), .ZN(
        n7395) );
  MOAI22 U16325 ( .A1(n28413), .A2(n887), .B1(ram[3155]), .B2(n888), .ZN(
        n7396) );
  MOAI22 U16326 ( .A1(n28178), .A2(n887), .B1(ram[3156]), .B2(n888), .ZN(
        n7397) );
  MOAI22 U16327 ( .A1(n27943), .A2(n887), .B1(ram[3157]), .B2(n888), .ZN(
        n7398) );
  MOAI22 U16328 ( .A1(n27708), .A2(n887), .B1(ram[3158]), .B2(n888), .ZN(
        n7399) );
  MOAI22 U16329 ( .A1(n27473), .A2(n887), .B1(ram[3159]), .B2(n888), .ZN(
        n7400) );
  MOAI22 U16330 ( .A1(n29118), .A2(n889), .B1(ram[3160]), .B2(n890), .ZN(
        n7401) );
  MOAI22 U16331 ( .A1(n28883), .A2(n889), .B1(ram[3161]), .B2(n890), .ZN(
        n7402) );
  MOAI22 U16332 ( .A1(n28648), .A2(n889), .B1(ram[3162]), .B2(n890), .ZN(
        n7403) );
  MOAI22 U16333 ( .A1(n28413), .A2(n889), .B1(ram[3163]), .B2(n890), .ZN(
        n7404) );
  MOAI22 U16334 ( .A1(n28178), .A2(n889), .B1(ram[3164]), .B2(n890), .ZN(
        n7405) );
  MOAI22 U16335 ( .A1(n27943), .A2(n889), .B1(ram[3165]), .B2(n890), .ZN(
        n7406) );
  MOAI22 U16336 ( .A1(n27708), .A2(n889), .B1(ram[3166]), .B2(n890), .ZN(
        n7407) );
  MOAI22 U16337 ( .A1(n27473), .A2(n889), .B1(ram[3167]), .B2(n890), .ZN(
        n7408) );
  MOAI22 U16338 ( .A1(n29118), .A2(n891), .B1(ram[3168]), .B2(n892), .ZN(
        n7409) );
  MOAI22 U16339 ( .A1(n28883), .A2(n891), .B1(ram[3169]), .B2(n892), .ZN(
        n7410) );
  MOAI22 U16340 ( .A1(n28648), .A2(n891), .B1(ram[3170]), .B2(n892), .ZN(
        n7411) );
  MOAI22 U16341 ( .A1(n28413), .A2(n891), .B1(ram[3171]), .B2(n892), .ZN(
        n7412) );
  MOAI22 U16342 ( .A1(n28178), .A2(n891), .B1(ram[3172]), .B2(n892), .ZN(
        n7413) );
  MOAI22 U16343 ( .A1(n27943), .A2(n891), .B1(ram[3173]), .B2(n892), .ZN(
        n7414) );
  MOAI22 U16344 ( .A1(n27708), .A2(n891), .B1(ram[3174]), .B2(n892), .ZN(
        n7415) );
  MOAI22 U16345 ( .A1(n27473), .A2(n891), .B1(ram[3175]), .B2(n892), .ZN(
        n7416) );
  MOAI22 U16346 ( .A1(n29118), .A2(n893), .B1(ram[3176]), .B2(n894), .ZN(
        n7417) );
  MOAI22 U16347 ( .A1(n28883), .A2(n893), .B1(ram[3177]), .B2(n894), .ZN(
        n7418) );
  MOAI22 U16348 ( .A1(n28648), .A2(n893), .B1(ram[3178]), .B2(n894), .ZN(
        n7419) );
  MOAI22 U16349 ( .A1(n28413), .A2(n893), .B1(ram[3179]), .B2(n894), .ZN(
        n7420) );
  MOAI22 U16350 ( .A1(n28178), .A2(n893), .B1(ram[3180]), .B2(n894), .ZN(
        n7421) );
  MOAI22 U16351 ( .A1(n27943), .A2(n893), .B1(ram[3181]), .B2(n894), .ZN(
        n7422) );
  MOAI22 U16352 ( .A1(n27708), .A2(n893), .B1(ram[3182]), .B2(n894), .ZN(
        n7423) );
  MOAI22 U16353 ( .A1(n27473), .A2(n893), .B1(ram[3183]), .B2(n894), .ZN(
        n7424) );
  MOAI22 U16354 ( .A1(n29118), .A2(n895), .B1(ram[3184]), .B2(n896), .ZN(
        n7425) );
  MOAI22 U16355 ( .A1(n28883), .A2(n895), .B1(ram[3185]), .B2(n896), .ZN(
        n7426) );
  MOAI22 U16356 ( .A1(n28648), .A2(n895), .B1(ram[3186]), .B2(n896), .ZN(
        n7427) );
  MOAI22 U16357 ( .A1(n28413), .A2(n895), .B1(ram[3187]), .B2(n896), .ZN(
        n7428) );
  MOAI22 U16358 ( .A1(n28178), .A2(n895), .B1(ram[3188]), .B2(n896), .ZN(
        n7429) );
  MOAI22 U16359 ( .A1(n27943), .A2(n895), .B1(ram[3189]), .B2(n896), .ZN(
        n7430) );
  MOAI22 U16360 ( .A1(n27708), .A2(n895), .B1(ram[3190]), .B2(n896), .ZN(
        n7431) );
  MOAI22 U16361 ( .A1(n27473), .A2(n895), .B1(ram[3191]), .B2(n896), .ZN(
        n7432) );
  MOAI22 U16362 ( .A1(n29118), .A2(n897), .B1(ram[3192]), .B2(n898), .ZN(
        n7433) );
  MOAI22 U16363 ( .A1(n28883), .A2(n897), .B1(ram[3193]), .B2(n898), .ZN(
        n7434) );
  MOAI22 U16364 ( .A1(n28648), .A2(n897), .B1(ram[3194]), .B2(n898), .ZN(
        n7435) );
  MOAI22 U16365 ( .A1(n28413), .A2(n897), .B1(ram[3195]), .B2(n898), .ZN(
        n7436) );
  MOAI22 U16366 ( .A1(n28178), .A2(n897), .B1(ram[3196]), .B2(n898), .ZN(
        n7437) );
  MOAI22 U16367 ( .A1(n27943), .A2(n897), .B1(ram[3197]), .B2(n898), .ZN(
        n7438) );
  MOAI22 U16368 ( .A1(n27708), .A2(n897), .B1(ram[3198]), .B2(n898), .ZN(
        n7439) );
  MOAI22 U16369 ( .A1(n27473), .A2(n897), .B1(ram[3199]), .B2(n898), .ZN(
        n7440) );
  MOAI22 U16370 ( .A1(n29118), .A2(n899), .B1(ram[3200]), .B2(n900), .ZN(
        n7441) );
  MOAI22 U16371 ( .A1(n28883), .A2(n899), .B1(ram[3201]), .B2(n900), .ZN(
        n7442) );
  MOAI22 U16372 ( .A1(n28648), .A2(n899), .B1(ram[3202]), .B2(n900), .ZN(
        n7443) );
  MOAI22 U16373 ( .A1(n28413), .A2(n899), .B1(ram[3203]), .B2(n900), .ZN(
        n7444) );
  MOAI22 U16374 ( .A1(n28178), .A2(n899), .B1(ram[3204]), .B2(n900), .ZN(
        n7445) );
  MOAI22 U16375 ( .A1(n27943), .A2(n899), .B1(ram[3205]), .B2(n900), .ZN(
        n7446) );
  MOAI22 U16376 ( .A1(n27708), .A2(n899), .B1(ram[3206]), .B2(n900), .ZN(
        n7447) );
  MOAI22 U16377 ( .A1(n27473), .A2(n899), .B1(ram[3207]), .B2(n900), .ZN(
        n7448) );
  MOAI22 U16378 ( .A1(n29118), .A2(n901), .B1(ram[3208]), .B2(n902), .ZN(
        n7449) );
  MOAI22 U16379 ( .A1(n28883), .A2(n901), .B1(ram[3209]), .B2(n902), .ZN(
        n7450) );
  MOAI22 U16380 ( .A1(n28648), .A2(n901), .B1(ram[3210]), .B2(n902), .ZN(
        n7451) );
  MOAI22 U16381 ( .A1(n28413), .A2(n901), .B1(ram[3211]), .B2(n902), .ZN(
        n7452) );
  MOAI22 U16382 ( .A1(n28178), .A2(n901), .B1(ram[3212]), .B2(n902), .ZN(
        n7453) );
  MOAI22 U16383 ( .A1(n27943), .A2(n901), .B1(ram[3213]), .B2(n902), .ZN(
        n7454) );
  MOAI22 U16384 ( .A1(n27708), .A2(n901), .B1(ram[3214]), .B2(n902), .ZN(
        n7455) );
  MOAI22 U16385 ( .A1(n27473), .A2(n901), .B1(ram[3215]), .B2(n902), .ZN(
        n7456) );
  MOAI22 U16386 ( .A1(n29118), .A2(n903), .B1(ram[3216]), .B2(n904), .ZN(
        n7457) );
  MOAI22 U16387 ( .A1(n28883), .A2(n903), .B1(ram[3217]), .B2(n904), .ZN(
        n7458) );
  MOAI22 U16388 ( .A1(n28648), .A2(n903), .B1(ram[3218]), .B2(n904), .ZN(
        n7459) );
  MOAI22 U16389 ( .A1(n28413), .A2(n903), .B1(ram[3219]), .B2(n904), .ZN(
        n7460) );
  MOAI22 U16390 ( .A1(n28178), .A2(n903), .B1(ram[3220]), .B2(n904), .ZN(
        n7461) );
  MOAI22 U16391 ( .A1(n27943), .A2(n903), .B1(ram[3221]), .B2(n904), .ZN(
        n7462) );
  MOAI22 U16392 ( .A1(n27708), .A2(n903), .B1(ram[3222]), .B2(n904), .ZN(
        n7463) );
  MOAI22 U16393 ( .A1(n27473), .A2(n903), .B1(ram[3223]), .B2(n904), .ZN(
        n7464) );
  MOAI22 U16394 ( .A1(n29119), .A2(n905), .B1(ram[3224]), .B2(n906), .ZN(
        n7465) );
  MOAI22 U16395 ( .A1(n28884), .A2(n905), .B1(ram[3225]), .B2(n906), .ZN(
        n7466) );
  MOAI22 U16396 ( .A1(n28649), .A2(n905), .B1(ram[3226]), .B2(n906), .ZN(
        n7467) );
  MOAI22 U16397 ( .A1(n28414), .A2(n905), .B1(ram[3227]), .B2(n906), .ZN(
        n7468) );
  MOAI22 U16398 ( .A1(n28179), .A2(n905), .B1(ram[3228]), .B2(n906), .ZN(
        n7469) );
  MOAI22 U16399 ( .A1(n27944), .A2(n905), .B1(ram[3229]), .B2(n906), .ZN(
        n7470) );
  MOAI22 U16400 ( .A1(n27709), .A2(n905), .B1(ram[3230]), .B2(n906), .ZN(
        n7471) );
  MOAI22 U16401 ( .A1(n27474), .A2(n905), .B1(ram[3231]), .B2(n906), .ZN(
        n7472) );
  MOAI22 U16402 ( .A1(n29119), .A2(n907), .B1(ram[3232]), .B2(n908), .ZN(
        n7473) );
  MOAI22 U16403 ( .A1(n28884), .A2(n907), .B1(ram[3233]), .B2(n908), .ZN(
        n7474) );
  MOAI22 U16404 ( .A1(n28649), .A2(n907), .B1(ram[3234]), .B2(n908), .ZN(
        n7475) );
  MOAI22 U16405 ( .A1(n28414), .A2(n907), .B1(ram[3235]), .B2(n908), .ZN(
        n7476) );
  MOAI22 U16406 ( .A1(n28179), .A2(n907), .B1(ram[3236]), .B2(n908), .ZN(
        n7477) );
  MOAI22 U16407 ( .A1(n27944), .A2(n907), .B1(ram[3237]), .B2(n908), .ZN(
        n7478) );
  MOAI22 U16408 ( .A1(n27709), .A2(n907), .B1(ram[3238]), .B2(n908), .ZN(
        n7479) );
  MOAI22 U16409 ( .A1(n27474), .A2(n907), .B1(ram[3239]), .B2(n908), .ZN(
        n7480) );
  MOAI22 U16410 ( .A1(n29119), .A2(n909), .B1(ram[3240]), .B2(n910), .ZN(
        n7481) );
  MOAI22 U16411 ( .A1(n28884), .A2(n909), .B1(ram[3241]), .B2(n910), .ZN(
        n7482) );
  MOAI22 U16412 ( .A1(n28649), .A2(n909), .B1(ram[3242]), .B2(n910), .ZN(
        n7483) );
  MOAI22 U16413 ( .A1(n28414), .A2(n909), .B1(ram[3243]), .B2(n910), .ZN(
        n7484) );
  MOAI22 U16414 ( .A1(n28179), .A2(n909), .B1(ram[3244]), .B2(n910), .ZN(
        n7485) );
  MOAI22 U16415 ( .A1(n27944), .A2(n909), .B1(ram[3245]), .B2(n910), .ZN(
        n7486) );
  MOAI22 U16416 ( .A1(n27709), .A2(n909), .B1(ram[3246]), .B2(n910), .ZN(
        n7487) );
  MOAI22 U16417 ( .A1(n27474), .A2(n909), .B1(ram[3247]), .B2(n910), .ZN(
        n7488) );
  MOAI22 U16418 ( .A1(n29119), .A2(n911), .B1(ram[3248]), .B2(n912), .ZN(
        n7489) );
  MOAI22 U16419 ( .A1(n28884), .A2(n911), .B1(ram[3249]), .B2(n912), .ZN(
        n7490) );
  MOAI22 U16420 ( .A1(n28649), .A2(n911), .B1(ram[3250]), .B2(n912), .ZN(
        n7491) );
  MOAI22 U16421 ( .A1(n28414), .A2(n911), .B1(ram[3251]), .B2(n912), .ZN(
        n7492) );
  MOAI22 U16422 ( .A1(n28179), .A2(n911), .B1(ram[3252]), .B2(n912), .ZN(
        n7493) );
  MOAI22 U16423 ( .A1(n27944), .A2(n911), .B1(ram[3253]), .B2(n912), .ZN(
        n7494) );
  MOAI22 U16424 ( .A1(n27709), .A2(n911), .B1(ram[3254]), .B2(n912), .ZN(
        n7495) );
  MOAI22 U16425 ( .A1(n27474), .A2(n911), .B1(ram[3255]), .B2(n912), .ZN(
        n7496) );
  MOAI22 U16426 ( .A1(n29119), .A2(n913), .B1(ram[3256]), .B2(n914), .ZN(
        n7497) );
  MOAI22 U16427 ( .A1(n28884), .A2(n913), .B1(ram[3257]), .B2(n914), .ZN(
        n7498) );
  MOAI22 U16428 ( .A1(n28649), .A2(n913), .B1(ram[3258]), .B2(n914), .ZN(
        n7499) );
  MOAI22 U16429 ( .A1(n28414), .A2(n913), .B1(ram[3259]), .B2(n914), .ZN(
        n7500) );
  MOAI22 U16430 ( .A1(n28179), .A2(n913), .B1(ram[3260]), .B2(n914), .ZN(
        n7501) );
  MOAI22 U16431 ( .A1(n27944), .A2(n913), .B1(ram[3261]), .B2(n914), .ZN(
        n7502) );
  MOAI22 U16432 ( .A1(n27709), .A2(n913), .B1(ram[3262]), .B2(n914), .ZN(
        n7503) );
  MOAI22 U16433 ( .A1(n27474), .A2(n913), .B1(ram[3263]), .B2(n914), .ZN(
        n7504) );
  MOAI22 U16434 ( .A1(n29119), .A2(n915), .B1(ram[3264]), .B2(n916), .ZN(
        n7505) );
  MOAI22 U16435 ( .A1(n28884), .A2(n915), .B1(ram[3265]), .B2(n916), .ZN(
        n7506) );
  MOAI22 U16436 ( .A1(n28649), .A2(n915), .B1(ram[3266]), .B2(n916), .ZN(
        n7507) );
  MOAI22 U16437 ( .A1(n28414), .A2(n915), .B1(ram[3267]), .B2(n916), .ZN(
        n7508) );
  MOAI22 U16438 ( .A1(n28179), .A2(n915), .B1(ram[3268]), .B2(n916), .ZN(
        n7509) );
  MOAI22 U16439 ( .A1(n27944), .A2(n915), .B1(ram[3269]), .B2(n916), .ZN(
        n7510) );
  MOAI22 U16440 ( .A1(n27709), .A2(n915), .B1(ram[3270]), .B2(n916), .ZN(
        n7511) );
  MOAI22 U16441 ( .A1(n27474), .A2(n915), .B1(ram[3271]), .B2(n916), .ZN(
        n7512) );
  MOAI22 U16442 ( .A1(n29119), .A2(n917), .B1(ram[3272]), .B2(n918), .ZN(
        n7513) );
  MOAI22 U16443 ( .A1(n28884), .A2(n917), .B1(ram[3273]), .B2(n918), .ZN(
        n7514) );
  MOAI22 U16444 ( .A1(n28649), .A2(n917), .B1(ram[3274]), .B2(n918), .ZN(
        n7515) );
  MOAI22 U16445 ( .A1(n28414), .A2(n917), .B1(ram[3275]), .B2(n918), .ZN(
        n7516) );
  MOAI22 U16446 ( .A1(n28179), .A2(n917), .B1(ram[3276]), .B2(n918), .ZN(
        n7517) );
  MOAI22 U16447 ( .A1(n27944), .A2(n917), .B1(ram[3277]), .B2(n918), .ZN(
        n7518) );
  MOAI22 U16448 ( .A1(n27709), .A2(n917), .B1(ram[3278]), .B2(n918), .ZN(
        n7519) );
  MOAI22 U16449 ( .A1(n27474), .A2(n917), .B1(ram[3279]), .B2(n918), .ZN(
        n7520) );
  MOAI22 U16450 ( .A1(n29119), .A2(n919), .B1(ram[3280]), .B2(n920), .ZN(
        n7521) );
  MOAI22 U16451 ( .A1(n28884), .A2(n919), .B1(ram[3281]), .B2(n920), .ZN(
        n7522) );
  MOAI22 U16452 ( .A1(n28649), .A2(n919), .B1(ram[3282]), .B2(n920), .ZN(
        n7523) );
  MOAI22 U16453 ( .A1(n28414), .A2(n919), .B1(ram[3283]), .B2(n920), .ZN(
        n7524) );
  MOAI22 U16454 ( .A1(n28179), .A2(n919), .B1(ram[3284]), .B2(n920), .ZN(
        n7525) );
  MOAI22 U16455 ( .A1(n27944), .A2(n919), .B1(ram[3285]), .B2(n920), .ZN(
        n7526) );
  MOAI22 U16456 ( .A1(n27709), .A2(n919), .B1(ram[3286]), .B2(n920), .ZN(
        n7527) );
  MOAI22 U16457 ( .A1(n27474), .A2(n919), .B1(ram[3287]), .B2(n920), .ZN(
        n7528) );
  MOAI22 U16458 ( .A1(n29119), .A2(n921), .B1(ram[3288]), .B2(n922), .ZN(
        n7529) );
  MOAI22 U16459 ( .A1(n28884), .A2(n921), .B1(ram[3289]), .B2(n922), .ZN(
        n7530) );
  MOAI22 U16460 ( .A1(n28649), .A2(n921), .B1(ram[3290]), .B2(n922), .ZN(
        n7531) );
  MOAI22 U16461 ( .A1(n28414), .A2(n921), .B1(ram[3291]), .B2(n922), .ZN(
        n7532) );
  MOAI22 U16462 ( .A1(n28179), .A2(n921), .B1(ram[3292]), .B2(n922), .ZN(
        n7533) );
  MOAI22 U16463 ( .A1(n27944), .A2(n921), .B1(ram[3293]), .B2(n922), .ZN(
        n7534) );
  MOAI22 U16464 ( .A1(n27709), .A2(n921), .B1(ram[3294]), .B2(n922), .ZN(
        n7535) );
  MOAI22 U16465 ( .A1(n27474), .A2(n921), .B1(ram[3295]), .B2(n922), .ZN(
        n7536) );
  MOAI22 U16466 ( .A1(n29119), .A2(n923), .B1(ram[3296]), .B2(n924), .ZN(
        n7537) );
  MOAI22 U16467 ( .A1(n28884), .A2(n923), .B1(ram[3297]), .B2(n924), .ZN(
        n7538) );
  MOAI22 U16468 ( .A1(n28649), .A2(n923), .B1(ram[3298]), .B2(n924), .ZN(
        n7539) );
  MOAI22 U16469 ( .A1(n28414), .A2(n923), .B1(ram[3299]), .B2(n924), .ZN(
        n7540) );
  MOAI22 U16470 ( .A1(n28179), .A2(n923), .B1(ram[3300]), .B2(n924), .ZN(
        n7541) );
  MOAI22 U16471 ( .A1(n27944), .A2(n923), .B1(ram[3301]), .B2(n924), .ZN(
        n7542) );
  MOAI22 U16472 ( .A1(n27709), .A2(n923), .B1(ram[3302]), .B2(n924), .ZN(
        n7543) );
  MOAI22 U16473 ( .A1(n27474), .A2(n923), .B1(ram[3303]), .B2(n924), .ZN(
        n7544) );
  MOAI22 U16474 ( .A1(n29119), .A2(n925), .B1(ram[3304]), .B2(n926), .ZN(
        n7545) );
  MOAI22 U16475 ( .A1(n28884), .A2(n925), .B1(ram[3305]), .B2(n926), .ZN(
        n7546) );
  MOAI22 U16476 ( .A1(n28649), .A2(n925), .B1(ram[3306]), .B2(n926), .ZN(
        n7547) );
  MOAI22 U16477 ( .A1(n28414), .A2(n925), .B1(ram[3307]), .B2(n926), .ZN(
        n7548) );
  MOAI22 U16478 ( .A1(n28179), .A2(n925), .B1(ram[3308]), .B2(n926), .ZN(
        n7549) );
  MOAI22 U16479 ( .A1(n27944), .A2(n925), .B1(ram[3309]), .B2(n926), .ZN(
        n7550) );
  MOAI22 U16480 ( .A1(n27709), .A2(n925), .B1(ram[3310]), .B2(n926), .ZN(
        n7551) );
  MOAI22 U16481 ( .A1(n27474), .A2(n925), .B1(ram[3311]), .B2(n926), .ZN(
        n7552) );
  MOAI22 U16482 ( .A1(n29119), .A2(n927), .B1(ram[3312]), .B2(n928), .ZN(
        n7553) );
  MOAI22 U16483 ( .A1(n28884), .A2(n927), .B1(ram[3313]), .B2(n928), .ZN(
        n7554) );
  MOAI22 U16484 ( .A1(n28649), .A2(n927), .B1(ram[3314]), .B2(n928), .ZN(
        n7555) );
  MOAI22 U16485 ( .A1(n28414), .A2(n927), .B1(ram[3315]), .B2(n928), .ZN(
        n7556) );
  MOAI22 U16486 ( .A1(n28179), .A2(n927), .B1(ram[3316]), .B2(n928), .ZN(
        n7557) );
  MOAI22 U16487 ( .A1(n27944), .A2(n927), .B1(ram[3317]), .B2(n928), .ZN(
        n7558) );
  MOAI22 U16488 ( .A1(n27709), .A2(n927), .B1(ram[3318]), .B2(n928), .ZN(
        n7559) );
  MOAI22 U16489 ( .A1(n27474), .A2(n927), .B1(ram[3319]), .B2(n928), .ZN(
        n7560) );
  MOAI22 U16490 ( .A1(n29119), .A2(n929), .B1(ram[3320]), .B2(n930), .ZN(
        n7561) );
  MOAI22 U16491 ( .A1(n28884), .A2(n929), .B1(ram[3321]), .B2(n930), .ZN(
        n7562) );
  MOAI22 U16492 ( .A1(n28649), .A2(n929), .B1(ram[3322]), .B2(n930), .ZN(
        n7563) );
  MOAI22 U16493 ( .A1(n28414), .A2(n929), .B1(ram[3323]), .B2(n930), .ZN(
        n7564) );
  MOAI22 U16494 ( .A1(n28179), .A2(n929), .B1(ram[3324]), .B2(n930), .ZN(
        n7565) );
  MOAI22 U16495 ( .A1(n27944), .A2(n929), .B1(ram[3325]), .B2(n930), .ZN(
        n7566) );
  MOAI22 U16496 ( .A1(n27709), .A2(n929), .B1(ram[3326]), .B2(n930), .ZN(
        n7567) );
  MOAI22 U16497 ( .A1(n27474), .A2(n929), .B1(ram[3327]), .B2(n930), .ZN(
        n7568) );
  MOAI22 U16498 ( .A1(n29120), .A2(n931), .B1(ram[3328]), .B2(n932), .ZN(
        n7569) );
  MOAI22 U16499 ( .A1(n28885), .A2(n931), .B1(ram[3329]), .B2(n932), .ZN(
        n7570) );
  MOAI22 U16500 ( .A1(n28650), .A2(n931), .B1(ram[3330]), .B2(n932), .ZN(
        n7571) );
  MOAI22 U16501 ( .A1(n28415), .A2(n931), .B1(ram[3331]), .B2(n932), .ZN(
        n7572) );
  MOAI22 U16502 ( .A1(n28180), .A2(n931), .B1(ram[3332]), .B2(n932), .ZN(
        n7573) );
  MOAI22 U16503 ( .A1(n27945), .A2(n931), .B1(ram[3333]), .B2(n932), .ZN(
        n7574) );
  MOAI22 U16504 ( .A1(n27710), .A2(n931), .B1(ram[3334]), .B2(n932), .ZN(
        n7575) );
  MOAI22 U16505 ( .A1(n27475), .A2(n931), .B1(ram[3335]), .B2(n932), .ZN(
        n7576) );
  MOAI22 U16506 ( .A1(n29120), .A2(n933), .B1(ram[3336]), .B2(n934), .ZN(
        n7577) );
  MOAI22 U16507 ( .A1(n28885), .A2(n933), .B1(ram[3337]), .B2(n934), .ZN(
        n7578) );
  MOAI22 U16508 ( .A1(n28650), .A2(n933), .B1(ram[3338]), .B2(n934), .ZN(
        n7579) );
  MOAI22 U16509 ( .A1(n28415), .A2(n933), .B1(ram[3339]), .B2(n934), .ZN(
        n7580) );
  MOAI22 U16510 ( .A1(n28180), .A2(n933), .B1(ram[3340]), .B2(n934), .ZN(
        n7581) );
  MOAI22 U16511 ( .A1(n27945), .A2(n933), .B1(ram[3341]), .B2(n934), .ZN(
        n7582) );
  MOAI22 U16512 ( .A1(n27710), .A2(n933), .B1(ram[3342]), .B2(n934), .ZN(
        n7583) );
  MOAI22 U16513 ( .A1(n27475), .A2(n933), .B1(ram[3343]), .B2(n934), .ZN(
        n7584) );
  MOAI22 U16514 ( .A1(n29120), .A2(n935), .B1(ram[3344]), .B2(n936), .ZN(
        n7585) );
  MOAI22 U16515 ( .A1(n28885), .A2(n935), .B1(ram[3345]), .B2(n936), .ZN(
        n7586) );
  MOAI22 U16516 ( .A1(n28650), .A2(n935), .B1(ram[3346]), .B2(n936), .ZN(
        n7587) );
  MOAI22 U16517 ( .A1(n28415), .A2(n935), .B1(ram[3347]), .B2(n936), .ZN(
        n7588) );
  MOAI22 U16518 ( .A1(n28180), .A2(n935), .B1(ram[3348]), .B2(n936), .ZN(
        n7589) );
  MOAI22 U16519 ( .A1(n27945), .A2(n935), .B1(ram[3349]), .B2(n936), .ZN(
        n7590) );
  MOAI22 U16520 ( .A1(n27710), .A2(n935), .B1(ram[3350]), .B2(n936), .ZN(
        n7591) );
  MOAI22 U16521 ( .A1(n27475), .A2(n935), .B1(ram[3351]), .B2(n936), .ZN(
        n7592) );
  MOAI22 U16522 ( .A1(n29120), .A2(n937), .B1(ram[3352]), .B2(n938), .ZN(
        n7593) );
  MOAI22 U16523 ( .A1(n28885), .A2(n937), .B1(ram[3353]), .B2(n938), .ZN(
        n7594) );
  MOAI22 U16524 ( .A1(n28650), .A2(n937), .B1(ram[3354]), .B2(n938), .ZN(
        n7595) );
  MOAI22 U16525 ( .A1(n28415), .A2(n937), .B1(ram[3355]), .B2(n938), .ZN(
        n7596) );
  MOAI22 U16526 ( .A1(n28180), .A2(n937), .B1(ram[3356]), .B2(n938), .ZN(
        n7597) );
  MOAI22 U16527 ( .A1(n27945), .A2(n937), .B1(ram[3357]), .B2(n938), .ZN(
        n7598) );
  MOAI22 U16528 ( .A1(n27710), .A2(n937), .B1(ram[3358]), .B2(n938), .ZN(
        n7599) );
  MOAI22 U16529 ( .A1(n27475), .A2(n937), .B1(ram[3359]), .B2(n938), .ZN(
        n7600) );
  MOAI22 U16530 ( .A1(n29120), .A2(n939), .B1(ram[3360]), .B2(n940), .ZN(
        n7601) );
  MOAI22 U16531 ( .A1(n28885), .A2(n939), .B1(ram[3361]), .B2(n940), .ZN(
        n7602) );
  MOAI22 U16532 ( .A1(n28650), .A2(n939), .B1(ram[3362]), .B2(n940), .ZN(
        n7603) );
  MOAI22 U16533 ( .A1(n28415), .A2(n939), .B1(ram[3363]), .B2(n940), .ZN(
        n7604) );
  MOAI22 U16534 ( .A1(n28180), .A2(n939), .B1(ram[3364]), .B2(n940), .ZN(
        n7605) );
  MOAI22 U16535 ( .A1(n27945), .A2(n939), .B1(ram[3365]), .B2(n940), .ZN(
        n7606) );
  MOAI22 U16536 ( .A1(n27710), .A2(n939), .B1(ram[3366]), .B2(n940), .ZN(
        n7607) );
  MOAI22 U16537 ( .A1(n27475), .A2(n939), .B1(ram[3367]), .B2(n940), .ZN(
        n7608) );
  MOAI22 U16538 ( .A1(n29120), .A2(n941), .B1(ram[3368]), .B2(n942), .ZN(
        n7609) );
  MOAI22 U16539 ( .A1(n28885), .A2(n941), .B1(ram[3369]), .B2(n942), .ZN(
        n7610) );
  MOAI22 U16540 ( .A1(n28650), .A2(n941), .B1(ram[3370]), .B2(n942), .ZN(
        n7611) );
  MOAI22 U16541 ( .A1(n28415), .A2(n941), .B1(ram[3371]), .B2(n942), .ZN(
        n7612) );
  MOAI22 U16542 ( .A1(n28180), .A2(n941), .B1(ram[3372]), .B2(n942), .ZN(
        n7613) );
  MOAI22 U16543 ( .A1(n27945), .A2(n941), .B1(ram[3373]), .B2(n942), .ZN(
        n7614) );
  MOAI22 U16544 ( .A1(n27710), .A2(n941), .B1(ram[3374]), .B2(n942), .ZN(
        n7615) );
  MOAI22 U16545 ( .A1(n27475), .A2(n941), .B1(ram[3375]), .B2(n942), .ZN(
        n7616) );
  MOAI22 U16546 ( .A1(n29120), .A2(n943), .B1(ram[3376]), .B2(n944), .ZN(
        n7617) );
  MOAI22 U16547 ( .A1(n28885), .A2(n943), .B1(ram[3377]), .B2(n944), .ZN(
        n7618) );
  MOAI22 U16548 ( .A1(n28650), .A2(n943), .B1(ram[3378]), .B2(n944), .ZN(
        n7619) );
  MOAI22 U16549 ( .A1(n28415), .A2(n943), .B1(ram[3379]), .B2(n944), .ZN(
        n7620) );
  MOAI22 U16550 ( .A1(n28180), .A2(n943), .B1(ram[3380]), .B2(n944), .ZN(
        n7621) );
  MOAI22 U16551 ( .A1(n27945), .A2(n943), .B1(ram[3381]), .B2(n944), .ZN(
        n7622) );
  MOAI22 U16552 ( .A1(n27710), .A2(n943), .B1(ram[3382]), .B2(n944), .ZN(
        n7623) );
  MOAI22 U16553 ( .A1(n27475), .A2(n943), .B1(ram[3383]), .B2(n944), .ZN(
        n7624) );
  MOAI22 U16554 ( .A1(n29120), .A2(n945), .B1(ram[3384]), .B2(n946), .ZN(
        n7625) );
  MOAI22 U16555 ( .A1(n28885), .A2(n945), .B1(ram[3385]), .B2(n946), .ZN(
        n7626) );
  MOAI22 U16556 ( .A1(n28650), .A2(n945), .B1(ram[3386]), .B2(n946), .ZN(
        n7627) );
  MOAI22 U16557 ( .A1(n28415), .A2(n945), .B1(ram[3387]), .B2(n946), .ZN(
        n7628) );
  MOAI22 U16558 ( .A1(n28180), .A2(n945), .B1(ram[3388]), .B2(n946), .ZN(
        n7629) );
  MOAI22 U16559 ( .A1(n27945), .A2(n945), .B1(ram[3389]), .B2(n946), .ZN(
        n7630) );
  MOAI22 U16560 ( .A1(n27710), .A2(n945), .B1(ram[3390]), .B2(n946), .ZN(
        n7631) );
  MOAI22 U16561 ( .A1(n27475), .A2(n945), .B1(ram[3391]), .B2(n946), .ZN(
        n7632) );
  MOAI22 U16562 ( .A1(n29120), .A2(n947), .B1(ram[3392]), .B2(n948), .ZN(
        n7633) );
  MOAI22 U16563 ( .A1(n28885), .A2(n947), .B1(ram[3393]), .B2(n948), .ZN(
        n7634) );
  MOAI22 U16564 ( .A1(n28650), .A2(n947), .B1(ram[3394]), .B2(n948), .ZN(
        n7635) );
  MOAI22 U16565 ( .A1(n28415), .A2(n947), .B1(ram[3395]), .B2(n948), .ZN(
        n7636) );
  MOAI22 U16566 ( .A1(n28180), .A2(n947), .B1(ram[3396]), .B2(n948), .ZN(
        n7637) );
  MOAI22 U16567 ( .A1(n27945), .A2(n947), .B1(ram[3397]), .B2(n948), .ZN(
        n7638) );
  MOAI22 U16568 ( .A1(n27710), .A2(n947), .B1(ram[3398]), .B2(n948), .ZN(
        n7639) );
  MOAI22 U16569 ( .A1(n27475), .A2(n947), .B1(ram[3399]), .B2(n948), .ZN(
        n7640) );
  MOAI22 U16570 ( .A1(n29120), .A2(n949), .B1(ram[3400]), .B2(n950), .ZN(
        n7641) );
  MOAI22 U16571 ( .A1(n28885), .A2(n949), .B1(ram[3401]), .B2(n950), .ZN(
        n7642) );
  MOAI22 U16572 ( .A1(n28650), .A2(n949), .B1(ram[3402]), .B2(n950), .ZN(
        n7643) );
  MOAI22 U16573 ( .A1(n28415), .A2(n949), .B1(ram[3403]), .B2(n950), .ZN(
        n7644) );
  MOAI22 U16574 ( .A1(n28180), .A2(n949), .B1(ram[3404]), .B2(n950), .ZN(
        n7645) );
  MOAI22 U16575 ( .A1(n27945), .A2(n949), .B1(ram[3405]), .B2(n950), .ZN(
        n7646) );
  MOAI22 U16576 ( .A1(n27710), .A2(n949), .B1(ram[3406]), .B2(n950), .ZN(
        n7647) );
  MOAI22 U16577 ( .A1(n27475), .A2(n949), .B1(ram[3407]), .B2(n950), .ZN(
        n7648) );
  MOAI22 U16578 ( .A1(n29120), .A2(n951), .B1(ram[3408]), .B2(n952), .ZN(
        n7649) );
  MOAI22 U16579 ( .A1(n28885), .A2(n951), .B1(ram[3409]), .B2(n952), .ZN(
        n7650) );
  MOAI22 U16580 ( .A1(n28650), .A2(n951), .B1(ram[3410]), .B2(n952), .ZN(
        n7651) );
  MOAI22 U16581 ( .A1(n28415), .A2(n951), .B1(ram[3411]), .B2(n952), .ZN(
        n7652) );
  MOAI22 U16582 ( .A1(n28180), .A2(n951), .B1(ram[3412]), .B2(n952), .ZN(
        n7653) );
  MOAI22 U16583 ( .A1(n27945), .A2(n951), .B1(ram[3413]), .B2(n952), .ZN(
        n7654) );
  MOAI22 U16584 ( .A1(n27710), .A2(n951), .B1(ram[3414]), .B2(n952), .ZN(
        n7655) );
  MOAI22 U16585 ( .A1(n27475), .A2(n951), .B1(ram[3415]), .B2(n952), .ZN(
        n7656) );
  MOAI22 U16586 ( .A1(n29120), .A2(n953), .B1(ram[3416]), .B2(n954), .ZN(
        n7657) );
  MOAI22 U16587 ( .A1(n28885), .A2(n953), .B1(ram[3417]), .B2(n954), .ZN(
        n7658) );
  MOAI22 U16588 ( .A1(n28650), .A2(n953), .B1(ram[3418]), .B2(n954), .ZN(
        n7659) );
  MOAI22 U16589 ( .A1(n28415), .A2(n953), .B1(ram[3419]), .B2(n954), .ZN(
        n7660) );
  MOAI22 U16590 ( .A1(n28180), .A2(n953), .B1(ram[3420]), .B2(n954), .ZN(
        n7661) );
  MOAI22 U16591 ( .A1(n27945), .A2(n953), .B1(ram[3421]), .B2(n954), .ZN(
        n7662) );
  MOAI22 U16592 ( .A1(n27710), .A2(n953), .B1(ram[3422]), .B2(n954), .ZN(
        n7663) );
  MOAI22 U16593 ( .A1(n27475), .A2(n953), .B1(ram[3423]), .B2(n954), .ZN(
        n7664) );
  MOAI22 U16594 ( .A1(n29120), .A2(n955), .B1(ram[3424]), .B2(n956), .ZN(
        n7665) );
  MOAI22 U16595 ( .A1(n28885), .A2(n955), .B1(ram[3425]), .B2(n956), .ZN(
        n7666) );
  MOAI22 U16596 ( .A1(n28650), .A2(n955), .B1(ram[3426]), .B2(n956), .ZN(
        n7667) );
  MOAI22 U16597 ( .A1(n28415), .A2(n955), .B1(ram[3427]), .B2(n956), .ZN(
        n7668) );
  MOAI22 U16598 ( .A1(n28180), .A2(n955), .B1(ram[3428]), .B2(n956), .ZN(
        n7669) );
  MOAI22 U16599 ( .A1(n27945), .A2(n955), .B1(ram[3429]), .B2(n956), .ZN(
        n7670) );
  MOAI22 U16600 ( .A1(n27710), .A2(n955), .B1(ram[3430]), .B2(n956), .ZN(
        n7671) );
  MOAI22 U16601 ( .A1(n27475), .A2(n955), .B1(ram[3431]), .B2(n956), .ZN(
        n7672) );
  MOAI22 U16602 ( .A1(n29121), .A2(n957), .B1(ram[3432]), .B2(n958), .ZN(
        n7673) );
  MOAI22 U16603 ( .A1(n28886), .A2(n957), .B1(ram[3433]), .B2(n958), .ZN(
        n7674) );
  MOAI22 U16604 ( .A1(n28651), .A2(n957), .B1(ram[3434]), .B2(n958), .ZN(
        n7675) );
  MOAI22 U16605 ( .A1(n28416), .A2(n957), .B1(ram[3435]), .B2(n958), .ZN(
        n7676) );
  MOAI22 U16606 ( .A1(n28181), .A2(n957), .B1(ram[3436]), .B2(n958), .ZN(
        n7677) );
  MOAI22 U16607 ( .A1(n27946), .A2(n957), .B1(ram[3437]), .B2(n958), .ZN(
        n7678) );
  MOAI22 U16608 ( .A1(n27711), .A2(n957), .B1(ram[3438]), .B2(n958), .ZN(
        n7679) );
  MOAI22 U16609 ( .A1(n27476), .A2(n957), .B1(ram[3439]), .B2(n958), .ZN(
        n7680) );
  MOAI22 U16610 ( .A1(n29121), .A2(n959), .B1(ram[3440]), .B2(n960), .ZN(
        n7681) );
  MOAI22 U16611 ( .A1(n28886), .A2(n959), .B1(ram[3441]), .B2(n960), .ZN(
        n7682) );
  MOAI22 U16612 ( .A1(n28651), .A2(n959), .B1(ram[3442]), .B2(n960), .ZN(
        n7683) );
  MOAI22 U16613 ( .A1(n28416), .A2(n959), .B1(ram[3443]), .B2(n960), .ZN(
        n7684) );
  MOAI22 U16614 ( .A1(n28181), .A2(n959), .B1(ram[3444]), .B2(n960), .ZN(
        n7685) );
  MOAI22 U16615 ( .A1(n27946), .A2(n959), .B1(ram[3445]), .B2(n960), .ZN(
        n7686) );
  MOAI22 U16616 ( .A1(n27711), .A2(n959), .B1(ram[3446]), .B2(n960), .ZN(
        n7687) );
  MOAI22 U16617 ( .A1(n27476), .A2(n959), .B1(ram[3447]), .B2(n960), .ZN(
        n7688) );
  MOAI22 U16618 ( .A1(n29121), .A2(n961), .B1(ram[3448]), .B2(n962), .ZN(
        n7689) );
  MOAI22 U16619 ( .A1(n28886), .A2(n961), .B1(ram[3449]), .B2(n962), .ZN(
        n7690) );
  MOAI22 U16620 ( .A1(n28651), .A2(n961), .B1(ram[3450]), .B2(n962), .ZN(
        n7691) );
  MOAI22 U16621 ( .A1(n28416), .A2(n961), .B1(ram[3451]), .B2(n962), .ZN(
        n7692) );
  MOAI22 U16622 ( .A1(n28181), .A2(n961), .B1(ram[3452]), .B2(n962), .ZN(
        n7693) );
  MOAI22 U16623 ( .A1(n27946), .A2(n961), .B1(ram[3453]), .B2(n962), .ZN(
        n7694) );
  MOAI22 U16624 ( .A1(n27711), .A2(n961), .B1(ram[3454]), .B2(n962), .ZN(
        n7695) );
  MOAI22 U16625 ( .A1(n27476), .A2(n961), .B1(ram[3455]), .B2(n962), .ZN(
        n7696) );
  MOAI22 U16626 ( .A1(n29121), .A2(n963), .B1(ram[3456]), .B2(n964), .ZN(
        n7697) );
  MOAI22 U16627 ( .A1(n28886), .A2(n963), .B1(ram[3457]), .B2(n964), .ZN(
        n7698) );
  MOAI22 U16628 ( .A1(n28651), .A2(n963), .B1(ram[3458]), .B2(n964), .ZN(
        n7699) );
  MOAI22 U16629 ( .A1(n28416), .A2(n963), .B1(ram[3459]), .B2(n964), .ZN(
        n7700) );
  MOAI22 U16630 ( .A1(n28181), .A2(n963), .B1(ram[3460]), .B2(n964), .ZN(
        n7701) );
  MOAI22 U16631 ( .A1(n27946), .A2(n963), .B1(ram[3461]), .B2(n964), .ZN(
        n7702) );
  MOAI22 U16632 ( .A1(n27711), .A2(n963), .B1(ram[3462]), .B2(n964), .ZN(
        n7703) );
  MOAI22 U16633 ( .A1(n27476), .A2(n963), .B1(ram[3463]), .B2(n964), .ZN(
        n7704) );
  MOAI22 U16634 ( .A1(n29121), .A2(n965), .B1(ram[3464]), .B2(n966), .ZN(
        n7705) );
  MOAI22 U16635 ( .A1(n28886), .A2(n965), .B1(ram[3465]), .B2(n966), .ZN(
        n7706) );
  MOAI22 U16636 ( .A1(n28651), .A2(n965), .B1(ram[3466]), .B2(n966), .ZN(
        n7707) );
  MOAI22 U16637 ( .A1(n28416), .A2(n965), .B1(ram[3467]), .B2(n966), .ZN(
        n7708) );
  MOAI22 U16638 ( .A1(n28181), .A2(n965), .B1(ram[3468]), .B2(n966), .ZN(
        n7709) );
  MOAI22 U16639 ( .A1(n27946), .A2(n965), .B1(ram[3469]), .B2(n966), .ZN(
        n7710) );
  MOAI22 U16640 ( .A1(n27711), .A2(n965), .B1(ram[3470]), .B2(n966), .ZN(
        n7711) );
  MOAI22 U16641 ( .A1(n27476), .A2(n965), .B1(ram[3471]), .B2(n966), .ZN(
        n7712) );
  MOAI22 U16642 ( .A1(n29121), .A2(n967), .B1(ram[3472]), .B2(n968), .ZN(
        n7713) );
  MOAI22 U16643 ( .A1(n28886), .A2(n967), .B1(ram[3473]), .B2(n968), .ZN(
        n7714) );
  MOAI22 U16644 ( .A1(n28651), .A2(n967), .B1(ram[3474]), .B2(n968), .ZN(
        n7715) );
  MOAI22 U16645 ( .A1(n28416), .A2(n967), .B1(ram[3475]), .B2(n968), .ZN(
        n7716) );
  MOAI22 U16646 ( .A1(n28181), .A2(n967), .B1(ram[3476]), .B2(n968), .ZN(
        n7717) );
  MOAI22 U16647 ( .A1(n27946), .A2(n967), .B1(ram[3477]), .B2(n968), .ZN(
        n7718) );
  MOAI22 U16648 ( .A1(n27711), .A2(n967), .B1(ram[3478]), .B2(n968), .ZN(
        n7719) );
  MOAI22 U16649 ( .A1(n27476), .A2(n967), .B1(ram[3479]), .B2(n968), .ZN(
        n7720) );
  MOAI22 U16650 ( .A1(n29121), .A2(n969), .B1(ram[3480]), .B2(n970), .ZN(
        n7721) );
  MOAI22 U16651 ( .A1(n28886), .A2(n969), .B1(ram[3481]), .B2(n970), .ZN(
        n7722) );
  MOAI22 U16652 ( .A1(n28651), .A2(n969), .B1(ram[3482]), .B2(n970), .ZN(
        n7723) );
  MOAI22 U16653 ( .A1(n28416), .A2(n969), .B1(ram[3483]), .B2(n970), .ZN(
        n7724) );
  MOAI22 U16654 ( .A1(n28181), .A2(n969), .B1(ram[3484]), .B2(n970), .ZN(
        n7725) );
  MOAI22 U16655 ( .A1(n27946), .A2(n969), .B1(ram[3485]), .B2(n970), .ZN(
        n7726) );
  MOAI22 U16656 ( .A1(n27711), .A2(n969), .B1(ram[3486]), .B2(n970), .ZN(
        n7727) );
  MOAI22 U16657 ( .A1(n27476), .A2(n969), .B1(ram[3487]), .B2(n970), .ZN(
        n7728) );
  MOAI22 U16658 ( .A1(n29121), .A2(n971), .B1(ram[3488]), .B2(n972), .ZN(
        n7729) );
  MOAI22 U16659 ( .A1(n28886), .A2(n971), .B1(ram[3489]), .B2(n972), .ZN(
        n7730) );
  MOAI22 U16660 ( .A1(n28651), .A2(n971), .B1(ram[3490]), .B2(n972), .ZN(
        n7731) );
  MOAI22 U16661 ( .A1(n28416), .A2(n971), .B1(ram[3491]), .B2(n972), .ZN(
        n7732) );
  MOAI22 U16662 ( .A1(n28181), .A2(n971), .B1(ram[3492]), .B2(n972), .ZN(
        n7733) );
  MOAI22 U16663 ( .A1(n27946), .A2(n971), .B1(ram[3493]), .B2(n972), .ZN(
        n7734) );
  MOAI22 U16664 ( .A1(n27711), .A2(n971), .B1(ram[3494]), .B2(n972), .ZN(
        n7735) );
  MOAI22 U16665 ( .A1(n27476), .A2(n971), .B1(ram[3495]), .B2(n972), .ZN(
        n7736) );
  MOAI22 U16666 ( .A1(n29121), .A2(n973), .B1(ram[3496]), .B2(n974), .ZN(
        n7737) );
  MOAI22 U16667 ( .A1(n28886), .A2(n973), .B1(ram[3497]), .B2(n974), .ZN(
        n7738) );
  MOAI22 U16668 ( .A1(n28651), .A2(n973), .B1(ram[3498]), .B2(n974), .ZN(
        n7739) );
  MOAI22 U16669 ( .A1(n28416), .A2(n973), .B1(ram[3499]), .B2(n974), .ZN(
        n7740) );
  MOAI22 U16670 ( .A1(n28181), .A2(n973), .B1(ram[3500]), .B2(n974), .ZN(
        n7741) );
  MOAI22 U16671 ( .A1(n27946), .A2(n973), .B1(ram[3501]), .B2(n974), .ZN(
        n7742) );
  MOAI22 U16672 ( .A1(n27711), .A2(n973), .B1(ram[3502]), .B2(n974), .ZN(
        n7743) );
  MOAI22 U16673 ( .A1(n27476), .A2(n973), .B1(ram[3503]), .B2(n974), .ZN(
        n7744) );
  MOAI22 U16674 ( .A1(n29121), .A2(n975), .B1(ram[3504]), .B2(n976), .ZN(
        n7745) );
  MOAI22 U16675 ( .A1(n28886), .A2(n975), .B1(ram[3505]), .B2(n976), .ZN(
        n7746) );
  MOAI22 U16676 ( .A1(n28651), .A2(n975), .B1(ram[3506]), .B2(n976), .ZN(
        n7747) );
  MOAI22 U16677 ( .A1(n28416), .A2(n975), .B1(ram[3507]), .B2(n976), .ZN(
        n7748) );
  MOAI22 U16678 ( .A1(n28181), .A2(n975), .B1(ram[3508]), .B2(n976), .ZN(
        n7749) );
  MOAI22 U16679 ( .A1(n27946), .A2(n975), .B1(ram[3509]), .B2(n976), .ZN(
        n7750) );
  MOAI22 U16680 ( .A1(n27711), .A2(n975), .B1(ram[3510]), .B2(n976), .ZN(
        n7751) );
  MOAI22 U16681 ( .A1(n27476), .A2(n975), .B1(ram[3511]), .B2(n976), .ZN(
        n7752) );
  MOAI22 U16682 ( .A1(n29121), .A2(n977), .B1(ram[3512]), .B2(n978), .ZN(
        n7753) );
  MOAI22 U16683 ( .A1(n28886), .A2(n977), .B1(ram[3513]), .B2(n978), .ZN(
        n7754) );
  MOAI22 U16684 ( .A1(n28651), .A2(n977), .B1(ram[3514]), .B2(n978), .ZN(
        n7755) );
  MOAI22 U16685 ( .A1(n28416), .A2(n977), .B1(ram[3515]), .B2(n978), .ZN(
        n7756) );
  MOAI22 U16686 ( .A1(n28181), .A2(n977), .B1(ram[3516]), .B2(n978), .ZN(
        n7757) );
  MOAI22 U16687 ( .A1(n27946), .A2(n977), .B1(ram[3517]), .B2(n978), .ZN(
        n7758) );
  MOAI22 U16688 ( .A1(n27711), .A2(n977), .B1(ram[3518]), .B2(n978), .ZN(
        n7759) );
  MOAI22 U16689 ( .A1(n27476), .A2(n977), .B1(ram[3519]), .B2(n978), .ZN(
        n7760) );
  MOAI22 U16690 ( .A1(n29121), .A2(n979), .B1(ram[3520]), .B2(n980), .ZN(
        n7761) );
  MOAI22 U16691 ( .A1(n28886), .A2(n979), .B1(ram[3521]), .B2(n980), .ZN(
        n7762) );
  MOAI22 U16692 ( .A1(n28651), .A2(n979), .B1(ram[3522]), .B2(n980), .ZN(
        n7763) );
  MOAI22 U16693 ( .A1(n28416), .A2(n979), .B1(ram[3523]), .B2(n980), .ZN(
        n7764) );
  MOAI22 U16694 ( .A1(n28181), .A2(n979), .B1(ram[3524]), .B2(n980), .ZN(
        n7765) );
  MOAI22 U16695 ( .A1(n27946), .A2(n979), .B1(ram[3525]), .B2(n980), .ZN(
        n7766) );
  MOAI22 U16696 ( .A1(n27711), .A2(n979), .B1(ram[3526]), .B2(n980), .ZN(
        n7767) );
  MOAI22 U16697 ( .A1(n27476), .A2(n979), .B1(ram[3527]), .B2(n980), .ZN(
        n7768) );
  MOAI22 U16698 ( .A1(n29121), .A2(n981), .B1(ram[3528]), .B2(n982), .ZN(
        n7769) );
  MOAI22 U16699 ( .A1(n28886), .A2(n981), .B1(ram[3529]), .B2(n982), .ZN(
        n7770) );
  MOAI22 U16700 ( .A1(n28651), .A2(n981), .B1(ram[3530]), .B2(n982), .ZN(
        n7771) );
  MOAI22 U16701 ( .A1(n28416), .A2(n981), .B1(ram[3531]), .B2(n982), .ZN(
        n7772) );
  MOAI22 U16702 ( .A1(n28181), .A2(n981), .B1(ram[3532]), .B2(n982), .ZN(
        n7773) );
  MOAI22 U16703 ( .A1(n27946), .A2(n981), .B1(ram[3533]), .B2(n982), .ZN(
        n7774) );
  MOAI22 U16704 ( .A1(n27711), .A2(n981), .B1(ram[3534]), .B2(n982), .ZN(
        n7775) );
  MOAI22 U16705 ( .A1(n27476), .A2(n981), .B1(ram[3535]), .B2(n982), .ZN(
        n7776) );
  MOAI22 U16706 ( .A1(n29122), .A2(n983), .B1(ram[3536]), .B2(n984), .ZN(
        n7777) );
  MOAI22 U16707 ( .A1(n28887), .A2(n983), .B1(ram[3537]), .B2(n984), .ZN(
        n7778) );
  MOAI22 U16708 ( .A1(n28652), .A2(n983), .B1(ram[3538]), .B2(n984), .ZN(
        n7779) );
  MOAI22 U16709 ( .A1(n28417), .A2(n983), .B1(ram[3539]), .B2(n984), .ZN(
        n7780) );
  MOAI22 U16710 ( .A1(n28182), .A2(n983), .B1(ram[3540]), .B2(n984), .ZN(
        n7781) );
  MOAI22 U16711 ( .A1(n27947), .A2(n983), .B1(ram[3541]), .B2(n984), .ZN(
        n7782) );
  MOAI22 U16712 ( .A1(n27712), .A2(n983), .B1(ram[3542]), .B2(n984), .ZN(
        n7783) );
  MOAI22 U16713 ( .A1(n27477), .A2(n983), .B1(ram[3543]), .B2(n984), .ZN(
        n7784) );
  MOAI22 U16714 ( .A1(n29122), .A2(n985), .B1(ram[3544]), .B2(n986), .ZN(
        n7785) );
  MOAI22 U16715 ( .A1(n28887), .A2(n985), .B1(ram[3545]), .B2(n986), .ZN(
        n7786) );
  MOAI22 U16716 ( .A1(n28652), .A2(n985), .B1(ram[3546]), .B2(n986), .ZN(
        n7787) );
  MOAI22 U16717 ( .A1(n28417), .A2(n985), .B1(ram[3547]), .B2(n986), .ZN(
        n7788) );
  MOAI22 U16718 ( .A1(n28182), .A2(n985), .B1(ram[3548]), .B2(n986), .ZN(
        n7789) );
  MOAI22 U16719 ( .A1(n27947), .A2(n985), .B1(ram[3549]), .B2(n986), .ZN(
        n7790) );
  MOAI22 U16720 ( .A1(n27712), .A2(n985), .B1(ram[3550]), .B2(n986), .ZN(
        n7791) );
  MOAI22 U16721 ( .A1(n27477), .A2(n985), .B1(ram[3551]), .B2(n986), .ZN(
        n7792) );
  MOAI22 U16722 ( .A1(n29122), .A2(n987), .B1(ram[3552]), .B2(n988), .ZN(
        n7793) );
  MOAI22 U16723 ( .A1(n28887), .A2(n987), .B1(ram[3553]), .B2(n988), .ZN(
        n7794) );
  MOAI22 U16724 ( .A1(n28652), .A2(n987), .B1(ram[3554]), .B2(n988), .ZN(
        n7795) );
  MOAI22 U16725 ( .A1(n28417), .A2(n987), .B1(ram[3555]), .B2(n988), .ZN(
        n7796) );
  MOAI22 U16726 ( .A1(n28182), .A2(n987), .B1(ram[3556]), .B2(n988), .ZN(
        n7797) );
  MOAI22 U16727 ( .A1(n27947), .A2(n987), .B1(ram[3557]), .B2(n988), .ZN(
        n7798) );
  MOAI22 U16728 ( .A1(n27712), .A2(n987), .B1(ram[3558]), .B2(n988), .ZN(
        n7799) );
  MOAI22 U16729 ( .A1(n27477), .A2(n987), .B1(ram[3559]), .B2(n988), .ZN(
        n7800) );
  MOAI22 U16730 ( .A1(n29122), .A2(n989), .B1(ram[3560]), .B2(n990), .ZN(
        n7801) );
  MOAI22 U16731 ( .A1(n28887), .A2(n989), .B1(ram[3561]), .B2(n990), .ZN(
        n7802) );
  MOAI22 U16732 ( .A1(n28652), .A2(n989), .B1(ram[3562]), .B2(n990), .ZN(
        n7803) );
  MOAI22 U16733 ( .A1(n28417), .A2(n989), .B1(ram[3563]), .B2(n990), .ZN(
        n7804) );
  MOAI22 U16734 ( .A1(n28182), .A2(n989), .B1(ram[3564]), .B2(n990), .ZN(
        n7805) );
  MOAI22 U16735 ( .A1(n27947), .A2(n989), .B1(ram[3565]), .B2(n990), .ZN(
        n7806) );
  MOAI22 U16736 ( .A1(n27712), .A2(n989), .B1(ram[3566]), .B2(n990), .ZN(
        n7807) );
  MOAI22 U16737 ( .A1(n27477), .A2(n989), .B1(ram[3567]), .B2(n990), .ZN(
        n7808) );
  MOAI22 U16738 ( .A1(n29122), .A2(n991), .B1(ram[3568]), .B2(n992), .ZN(
        n7809) );
  MOAI22 U16739 ( .A1(n28887), .A2(n991), .B1(ram[3569]), .B2(n992), .ZN(
        n7810) );
  MOAI22 U16740 ( .A1(n28652), .A2(n991), .B1(ram[3570]), .B2(n992), .ZN(
        n7811) );
  MOAI22 U16741 ( .A1(n28417), .A2(n991), .B1(ram[3571]), .B2(n992), .ZN(
        n7812) );
  MOAI22 U16742 ( .A1(n28182), .A2(n991), .B1(ram[3572]), .B2(n992), .ZN(
        n7813) );
  MOAI22 U16743 ( .A1(n27947), .A2(n991), .B1(ram[3573]), .B2(n992), .ZN(
        n7814) );
  MOAI22 U16744 ( .A1(n27712), .A2(n991), .B1(ram[3574]), .B2(n992), .ZN(
        n7815) );
  MOAI22 U16745 ( .A1(n27477), .A2(n991), .B1(ram[3575]), .B2(n992), .ZN(
        n7816) );
  MOAI22 U16746 ( .A1(n29122), .A2(n993), .B1(ram[3576]), .B2(n994), .ZN(
        n7817) );
  MOAI22 U16747 ( .A1(n28887), .A2(n993), .B1(ram[3577]), .B2(n994), .ZN(
        n7818) );
  MOAI22 U16748 ( .A1(n28652), .A2(n993), .B1(ram[3578]), .B2(n994), .ZN(
        n7819) );
  MOAI22 U16749 ( .A1(n28417), .A2(n993), .B1(ram[3579]), .B2(n994), .ZN(
        n7820) );
  MOAI22 U16750 ( .A1(n28182), .A2(n993), .B1(ram[3580]), .B2(n994), .ZN(
        n7821) );
  MOAI22 U16751 ( .A1(n27947), .A2(n993), .B1(ram[3581]), .B2(n994), .ZN(
        n7822) );
  MOAI22 U16752 ( .A1(n27712), .A2(n993), .B1(ram[3582]), .B2(n994), .ZN(
        n7823) );
  MOAI22 U16753 ( .A1(n27477), .A2(n993), .B1(ram[3583]), .B2(n994), .ZN(
        n7824) );
  MOAI22 U16754 ( .A1(n29122), .A2(n996), .B1(ram[3584]), .B2(n997), .ZN(
        n7825) );
  MOAI22 U16755 ( .A1(n28887), .A2(n996), .B1(ram[3585]), .B2(n997), .ZN(
        n7826) );
  MOAI22 U16756 ( .A1(n28652), .A2(n996), .B1(ram[3586]), .B2(n997), .ZN(
        n7827) );
  MOAI22 U16757 ( .A1(n28417), .A2(n996), .B1(ram[3587]), .B2(n997), .ZN(
        n7828) );
  MOAI22 U16758 ( .A1(n28182), .A2(n996), .B1(ram[3588]), .B2(n997), .ZN(
        n7829) );
  MOAI22 U16759 ( .A1(n27947), .A2(n996), .B1(ram[3589]), .B2(n997), .ZN(
        n7830) );
  MOAI22 U16760 ( .A1(n27712), .A2(n996), .B1(ram[3590]), .B2(n997), .ZN(
        n7831) );
  MOAI22 U16761 ( .A1(n27477), .A2(n996), .B1(ram[3591]), .B2(n997), .ZN(
        n7832) );
  MOAI22 U16762 ( .A1(n29122), .A2(n999), .B1(ram[3592]), .B2(n1000), 
        .ZN(n7833) );
  MOAI22 U16763 ( .A1(n28887), .A2(n999), .B1(ram[3593]), .B2(n1000), 
        .ZN(n7834) );
  MOAI22 U16764 ( .A1(n28652), .A2(n999), .B1(ram[3594]), .B2(n1000), 
        .ZN(n7835) );
  MOAI22 U16765 ( .A1(n28417), .A2(n999), .B1(ram[3595]), .B2(n1000), 
        .ZN(n7836) );
  MOAI22 U16766 ( .A1(n28182), .A2(n999), .B1(ram[3596]), .B2(n1000), 
        .ZN(n7837) );
  MOAI22 U16767 ( .A1(n27947), .A2(n999), .B1(ram[3597]), .B2(n1000), 
        .ZN(n7838) );
  MOAI22 U16768 ( .A1(n27712), .A2(n999), .B1(ram[3598]), .B2(n1000), 
        .ZN(n7839) );
  MOAI22 U16769 ( .A1(n27477), .A2(n999), .B1(ram[3599]), .B2(n1000), 
        .ZN(n7840) );
  MOAI22 U16770 ( .A1(n29122), .A2(n1001), .B1(ram[3600]), .B2(n1002), 
        .ZN(n7841) );
  MOAI22 U16771 ( .A1(n28887), .A2(n1001), .B1(ram[3601]), .B2(n1002), 
        .ZN(n7842) );
  MOAI22 U16772 ( .A1(n28652), .A2(n1001), .B1(ram[3602]), .B2(n1002), 
        .ZN(n7843) );
  MOAI22 U16773 ( .A1(n28417), .A2(n1001), .B1(ram[3603]), .B2(n1002), 
        .ZN(n7844) );
  MOAI22 U16774 ( .A1(n28182), .A2(n1001), .B1(ram[3604]), .B2(n1002), 
        .ZN(n7845) );
  MOAI22 U16775 ( .A1(n27947), .A2(n1001), .B1(ram[3605]), .B2(n1002), 
        .ZN(n7846) );
  MOAI22 U16776 ( .A1(n27712), .A2(n1001), .B1(ram[3606]), .B2(n1002), 
        .ZN(n7847) );
  MOAI22 U16777 ( .A1(n27477), .A2(n1001), .B1(ram[3607]), .B2(n1002), 
        .ZN(n7848) );
  MOAI22 U16778 ( .A1(n29122), .A2(n1003), .B1(ram[3608]), .B2(n1004), 
        .ZN(n7849) );
  MOAI22 U16779 ( .A1(n28887), .A2(n1003), .B1(ram[3609]), .B2(n1004), 
        .ZN(n7850) );
  MOAI22 U16780 ( .A1(n28652), .A2(n1003), .B1(ram[3610]), .B2(n1004), 
        .ZN(n7851) );
  MOAI22 U16781 ( .A1(n28417), .A2(n1003), .B1(ram[3611]), .B2(n1004), 
        .ZN(n7852) );
  MOAI22 U16782 ( .A1(n28182), .A2(n1003), .B1(ram[3612]), .B2(n1004), 
        .ZN(n7853) );
  MOAI22 U16783 ( .A1(n27947), .A2(n1003), .B1(ram[3613]), .B2(n1004), 
        .ZN(n7854) );
  MOAI22 U16784 ( .A1(n27712), .A2(n1003), .B1(ram[3614]), .B2(n1004), 
        .ZN(n7855) );
  MOAI22 U16785 ( .A1(n27477), .A2(n1003), .B1(ram[3615]), .B2(n1004), 
        .ZN(n7856) );
  MOAI22 U16786 ( .A1(n29122), .A2(n1005), .B1(ram[3616]), .B2(n1006), 
        .ZN(n7857) );
  MOAI22 U16787 ( .A1(n28887), .A2(n1005), .B1(ram[3617]), .B2(n1006), 
        .ZN(n7858) );
  MOAI22 U16788 ( .A1(n28652), .A2(n1005), .B1(ram[3618]), .B2(n1006), 
        .ZN(n7859) );
  MOAI22 U16789 ( .A1(n28417), .A2(n1005), .B1(ram[3619]), .B2(n1006), 
        .ZN(n7860) );
  MOAI22 U16790 ( .A1(n28182), .A2(n1005), .B1(ram[3620]), .B2(n1006), 
        .ZN(n7861) );
  MOAI22 U16791 ( .A1(n27947), .A2(n1005), .B1(ram[3621]), .B2(n1006), 
        .ZN(n7862) );
  MOAI22 U16792 ( .A1(n27712), .A2(n1005), .B1(ram[3622]), .B2(n1006), 
        .ZN(n7863) );
  MOAI22 U16793 ( .A1(n27477), .A2(n1005), .B1(ram[3623]), .B2(n1006), 
        .ZN(n7864) );
  MOAI22 U16794 ( .A1(n29122), .A2(n1007), .B1(ram[3624]), .B2(n1008), 
        .ZN(n7865) );
  MOAI22 U16795 ( .A1(n28887), .A2(n1007), .B1(ram[3625]), .B2(n1008), 
        .ZN(n7866) );
  MOAI22 U16796 ( .A1(n28652), .A2(n1007), .B1(ram[3626]), .B2(n1008), 
        .ZN(n7867) );
  MOAI22 U16797 ( .A1(n28417), .A2(n1007), .B1(ram[3627]), .B2(n1008), 
        .ZN(n7868) );
  MOAI22 U16798 ( .A1(n28182), .A2(n1007), .B1(ram[3628]), .B2(n1008), 
        .ZN(n7869) );
  MOAI22 U16799 ( .A1(n27947), .A2(n1007), .B1(ram[3629]), .B2(n1008), 
        .ZN(n7870) );
  MOAI22 U16800 ( .A1(n27712), .A2(n1007), .B1(ram[3630]), .B2(n1008), 
        .ZN(n7871) );
  MOAI22 U16801 ( .A1(n27477), .A2(n1007), .B1(ram[3631]), .B2(n1008), 
        .ZN(n7872) );
  MOAI22 U16802 ( .A1(n29122), .A2(n1009), .B1(ram[3632]), .B2(n1010), 
        .ZN(n7873) );
  MOAI22 U16803 ( .A1(n28887), .A2(n1009), .B1(ram[3633]), .B2(n1010), 
        .ZN(n7874) );
  MOAI22 U16804 ( .A1(n28652), .A2(n1009), .B1(ram[3634]), .B2(n1010), 
        .ZN(n7875) );
  MOAI22 U16805 ( .A1(n28417), .A2(n1009), .B1(ram[3635]), .B2(n1010), 
        .ZN(n7876) );
  MOAI22 U16806 ( .A1(n28182), .A2(n1009), .B1(ram[3636]), .B2(n1010), 
        .ZN(n7877) );
  MOAI22 U16807 ( .A1(n27947), .A2(n1009), .B1(ram[3637]), .B2(n1010), 
        .ZN(n7878) );
  MOAI22 U16808 ( .A1(n27712), .A2(n1009), .B1(ram[3638]), .B2(n1010), 
        .ZN(n7879) );
  MOAI22 U16809 ( .A1(n27477), .A2(n1009), .B1(ram[3639]), .B2(n1010), 
        .ZN(n7880) );
  MOAI22 U16810 ( .A1(n29123), .A2(n1011), .B1(ram[3640]), .B2(n1012), 
        .ZN(n7881) );
  MOAI22 U16811 ( .A1(n28888), .A2(n1011), .B1(ram[3641]), .B2(n1012), 
        .ZN(n7882) );
  MOAI22 U16812 ( .A1(n28653), .A2(n1011), .B1(ram[3642]), .B2(n1012), 
        .ZN(n7883) );
  MOAI22 U16813 ( .A1(n28418), .A2(n1011), .B1(ram[3643]), .B2(n1012), 
        .ZN(n7884) );
  MOAI22 U16814 ( .A1(n28183), .A2(n1011), .B1(ram[3644]), .B2(n1012), 
        .ZN(n7885) );
  MOAI22 U16815 ( .A1(n27948), .A2(n1011), .B1(ram[3645]), .B2(n1012), 
        .ZN(n7886) );
  MOAI22 U16816 ( .A1(n27713), .A2(n1011), .B1(ram[3646]), .B2(n1012), 
        .ZN(n7887) );
  MOAI22 U16817 ( .A1(n27478), .A2(n1011), .B1(ram[3647]), .B2(n1012), 
        .ZN(n7888) );
  MOAI22 U16818 ( .A1(n29123), .A2(n1013), .B1(ram[3648]), .B2(n1014), 
        .ZN(n7889) );
  MOAI22 U16819 ( .A1(n28888), .A2(n1013), .B1(ram[3649]), .B2(n1014), 
        .ZN(n7890) );
  MOAI22 U16820 ( .A1(n28653), .A2(n1013), .B1(ram[3650]), .B2(n1014), 
        .ZN(n7891) );
  MOAI22 U16821 ( .A1(n28418), .A2(n1013), .B1(ram[3651]), .B2(n1014), 
        .ZN(n7892) );
  MOAI22 U16822 ( .A1(n28183), .A2(n1013), .B1(ram[3652]), .B2(n1014), 
        .ZN(n7893) );
  MOAI22 U16823 ( .A1(n27948), .A2(n1013), .B1(ram[3653]), .B2(n1014), 
        .ZN(n7894) );
  MOAI22 U16824 ( .A1(n27713), .A2(n1013), .B1(ram[3654]), .B2(n1014), 
        .ZN(n7895) );
  MOAI22 U16825 ( .A1(n27478), .A2(n1013), .B1(ram[3655]), .B2(n1014), 
        .ZN(n7896) );
  MOAI22 U16826 ( .A1(n29123), .A2(n1015), .B1(ram[3656]), .B2(n1016), 
        .ZN(n7897) );
  MOAI22 U16827 ( .A1(n28888), .A2(n1015), .B1(ram[3657]), .B2(n1016), 
        .ZN(n7898) );
  MOAI22 U16828 ( .A1(n28653), .A2(n1015), .B1(ram[3658]), .B2(n1016), 
        .ZN(n7899) );
  MOAI22 U16829 ( .A1(n28418), .A2(n1015), .B1(ram[3659]), .B2(n1016), 
        .ZN(n7900) );
  MOAI22 U16830 ( .A1(n28183), .A2(n1015), .B1(ram[3660]), .B2(n1016), 
        .ZN(n7901) );
  MOAI22 U16831 ( .A1(n27948), .A2(n1015), .B1(ram[3661]), .B2(n1016), 
        .ZN(n7902) );
  MOAI22 U16832 ( .A1(n27713), .A2(n1015), .B1(ram[3662]), .B2(n1016), 
        .ZN(n7903) );
  MOAI22 U16833 ( .A1(n27478), .A2(n1015), .B1(ram[3663]), .B2(n1016), 
        .ZN(n7904) );
  MOAI22 U16834 ( .A1(n29123), .A2(n1017), .B1(ram[3664]), .B2(n1018), 
        .ZN(n7905) );
  MOAI22 U16835 ( .A1(n28888), .A2(n1017), .B1(ram[3665]), .B2(n1018), 
        .ZN(n7906) );
  MOAI22 U16836 ( .A1(n28653), .A2(n1017), .B1(ram[3666]), .B2(n1018), 
        .ZN(n7907) );
  MOAI22 U16837 ( .A1(n28418), .A2(n1017), .B1(ram[3667]), .B2(n1018), 
        .ZN(n7908) );
  MOAI22 U16838 ( .A1(n28183), .A2(n1017), .B1(ram[3668]), .B2(n1018), 
        .ZN(n7909) );
  MOAI22 U16839 ( .A1(n27948), .A2(n1017), .B1(ram[3669]), .B2(n1018), 
        .ZN(n7910) );
  MOAI22 U16840 ( .A1(n27713), .A2(n1017), .B1(ram[3670]), .B2(n1018), 
        .ZN(n7911) );
  MOAI22 U16841 ( .A1(n27478), .A2(n1017), .B1(ram[3671]), .B2(n1018), 
        .ZN(n7912) );
  MOAI22 U16842 ( .A1(n29123), .A2(n1019), .B1(ram[3672]), .B2(n1020), 
        .ZN(n7913) );
  MOAI22 U16843 ( .A1(n28888), .A2(n1019), .B1(ram[3673]), .B2(n1020), 
        .ZN(n7914) );
  MOAI22 U16844 ( .A1(n28653), .A2(n1019), .B1(ram[3674]), .B2(n1020), 
        .ZN(n7915) );
  MOAI22 U16845 ( .A1(n28418), .A2(n1019), .B1(ram[3675]), .B2(n1020), 
        .ZN(n7916) );
  MOAI22 U16846 ( .A1(n28183), .A2(n1019), .B1(ram[3676]), .B2(n1020), 
        .ZN(n7917) );
  MOAI22 U16847 ( .A1(n27948), .A2(n1019), .B1(ram[3677]), .B2(n1020), 
        .ZN(n7918) );
  MOAI22 U16848 ( .A1(n27713), .A2(n1019), .B1(ram[3678]), .B2(n1020), 
        .ZN(n7919) );
  MOAI22 U16849 ( .A1(n27478), .A2(n1019), .B1(ram[3679]), .B2(n1020), 
        .ZN(n7920) );
  MOAI22 U16850 ( .A1(n29123), .A2(n1021), .B1(ram[3680]), .B2(n1022), 
        .ZN(n7921) );
  MOAI22 U16851 ( .A1(n28888), .A2(n1021), .B1(ram[3681]), .B2(n1022), 
        .ZN(n7922) );
  MOAI22 U16852 ( .A1(n28653), .A2(n1021), .B1(ram[3682]), .B2(n1022), 
        .ZN(n7923) );
  MOAI22 U16853 ( .A1(n28418), .A2(n1021), .B1(ram[3683]), .B2(n1022), 
        .ZN(n7924) );
  MOAI22 U16854 ( .A1(n28183), .A2(n1021), .B1(ram[3684]), .B2(n1022), 
        .ZN(n7925) );
  MOAI22 U16855 ( .A1(n27948), .A2(n1021), .B1(ram[3685]), .B2(n1022), 
        .ZN(n7926) );
  MOAI22 U16856 ( .A1(n27713), .A2(n1021), .B1(ram[3686]), .B2(n1022), 
        .ZN(n7927) );
  MOAI22 U16857 ( .A1(n27478), .A2(n1021), .B1(ram[3687]), .B2(n1022), 
        .ZN(n7928) );
  MOAI22 U16858 ( .A1(n29123), .A2(n1023), .B1(ram[3688]), .B2(n1024), 
        .ZN(n7929) );
  MOAI22 U16859 ( .A1(n28888), .A2(n1023), .B1(ram[3689]), .B2(n1024), 
        .ZN(n7930) );
  MOAI22 U16860 ( .A1(n28653), .A2(n1023), .B1(ram[3690]), .B2(n1024), 
        .ZN(n7931) );
  MOAI22 U16861 ( .A1(n28418), .A2(n1023), .B1(ram[3691]), .B2(n1024), 
        .ZN(n7932) );
  MOAI22 U16862 ( .A1(n28183), .A2(n1023), .B1(ram[3692]), .B2(n1024), 
        .ZN(n7933) );
  MOAI22 U16863 ( .A1(n27948), .A2(n1023), .B1(ram[3693]), .B2(n1024), 
        .ZN(n7934) );
  MOAI22 U16864 ( .A1(n27713), .A2(n1023), .B1(ram[3694]), .B2(n1024), 
        .ZN(n7935) );
  MOAI22 U16865 ( .A1(n27478), .A2(n1023), .B1(ram[3695]), .B2(n1024), 
        .ZN(n7936) );
  MOAI22 U16866 ( .A1(n29123), .A2(n1025), .B1(ram[3696]), .B2(n1026), 
        .ZN(n7937) );
  MOAI22 U16867 ( .A1(n28888), .A2(n1025), .B1(ram[3697]), .B2(n1026), 
        .ZN(n7938) );
  MOAI22 U16868 ( .A1(n28653), .A2(n1025), .B1(ram[3698]), .B2(n1026), 
        .ZN(n7939) );
  MOAI22 U16869 ( .A1(n28418), .A2(n1025), .B1(ram[3699]), .B2(n1026), 
        .ZN(n7940) );
  MOAI22 U16870 ( .A1(n28183), .A2(n1025), .B1(ram[3700]), .B2(n1026), 
        .ZN(n7941) );
  MOAI22 U16871 ( .A1(n27948), .A2(n1025), .B1(ram[3701]), .B2(n1026), 
        .ZN(n7942) );
  MOAI22 U16872 ( .A1(n27713), .A2(n1025), .B1(ram[3702]), .B2(n1026), 
        .ZN(n7943) );
  MOAI22 U16873 ( .A1(n27478), .A2(n1025), .B1(ram[3703]), .B2(n1026), 
        .ZN(n7944) );
  MOAI22 U16874 ( .A1(n29123), .A2(n1027), .B1(ram[3704]), .B2(n1028), 
        .ZN(n7945) );
  MOAI22 U16875 ( .A1(n28888), .A2(n1027), .B1(ram[3705]), .B2(n1028), 
        .ZN(n7946) );
  MOAI22 U16876 ( .A1(n28653), .A2(n1027), .B1(ram[3706]), .B2(n1028), 
        .ZN(n7947) );
  MOAI22 U16877 ( .A1(n28418), .A2(n1027), .B1(ram[3707]), .B2(n1028), 
        .ZN(n7948) );
  MOAI22 U16878 ( .A1(n28183), .A2(n1027), .B1(ram[3708]), .B2(n1028), 
        .ZN(n7949) );
  MOAI22 U16879 ( .A1(n27948), .A2(n1027), .B1(ram[3709]), .B2(n1028), 
        .ZN(n7950) );
  MOAI22 U16880 ( .A1(n27713), .A2(n1027), .B1(ram[3710]), .B2(n1028), 
        .ZN(n7951) );
  MOAI22 U16881 ( .A1(n27478), .A2(n1027), .B1(ram[3711]), .B2(n1028), 
        .ZN(n7952) );
  MOAI22 U16882 ( .A1(n29123), .A2(n1029), .B1(ram[3712]), .B2(n1030), 
        .ZN(n7953) );
  MOAI22 U16883 ( .A1(n28888), .A2(n1029), .B1(ram[3713]), .B2(n1030), 
        .ZN(n7954) );
  MOAI22 U16884 ( .A1(n28653), .A2(n1029), .B1(ram[3714]), .B2(n1030), 
        .ZN(n7955) );
  MOAI22 U16885 ( .A1(n28418), .A2(n1029), .B1(ram[3715]), .B2(n1030), 
        .ZN(n7956) );
  MOAI22 U16886 ( .A1(n28183), .A2(n1029), .B1(ram[3716]), .B2(n1030), 
        .ZN(n7957) );
  MOAI22 U16887 ( .A1(n27948), .A2(n1029), .B1(ram[3717]), .B2(n1030), 
        .ZN(n7958) );
  MOAI22 U16888 ( .A1(n27713), .A2(n1029), .B1(ram[3718]), .B2(n1030), 
        .ZN(n7959) );
  MOAI22 U16889 ( .A1(n27478), .A2(n1029), .B1(ram[3719]), .B2(n1030), 
        .ZN(n7960) );
  MOAI22 U16890 ( .A1(n29123), .A2(n1031), .B1(ram[3720]), .B2(n1032), 
        .ZN(n7961) );
  MOAI22 U16891 ( .A1(n28888), .A2(n1031), .B1(ram[3721]), .B2(n1032), 
        .ZN(n7962) );
  MOAI22 U16892 ( .A1(n28653), .A2(n1031), .B1(ram[3722]), .B2(n1032), 
        .ZN(n7963) );
  MOAI22 U16893 ( .A1(n28418), .A2(n1031), .B1(ram[3723]), .B2(n1032), 
        .ZN(n7964) );
  MOAI22 U16894 ( .A1(n28183), .A2(n1031), .B1(ram[3724]), .B2(n1032), 
        .ZN(n7965) );
  MOAI22 U16895 ( .A1(n27948), .A2(n1031), .B1(ram[3725]), .B2(n1032), 
        .ZN(n7966) );
  MOAI22 U16896 ( .A1(n27713), .A2(n1031), .B1(ram[3726]), .B2(n1032), 
        .ZN(n7967) );
  MOAI22 U16897 ( .A1(n27478), .A2(n1031), .B1(ram[3727]), .B2(n1032), 
        .ZN(n7968) );
  MOAI22 U16898 ( .A1(n29123), .A2(n1033), .B1(ram[3728]), .B2(n1034), 
        .ZN(n7969) );
  MOAI22 U16899 ( .A1(n28888), .A2(n1033), .B1(ram[3729]), .B2(n1034), 
        .ZN(n7970) );
  MOAI22 U16900 ( .A1(n28653), .A2(n1033), .B1(ram[3730]), .B2(n1034), 
        .ZN(n7971) );
  MOAI22 U16901 ( .A1(n28418), .A2(n1033), .B1(ram[3731]), .B2(n1034), 
        .ZN(n7972) );
  MOAI22 U16902 ( .A1(n28183), .A2(n1033), .B1(ram[3732]), .B2(n1034), 
        .ZN(n7973) );
  MOAI22 U16903 ( .A1(n27948), .A2(n1033), .B1(ram[3733]), .B2(n1034), 
        .ZN(n7974) );
  MOAI22 U16904 ( .A1(n27713), .A2(n1033), .B1(ram[3734]), .B2(n1034), 
        .ZN(n7975) );
  MOAI22 U16905 ( .A1(n27478), .A2(n1033), .B1(ram[3735]), .B2(n1034), 
        .ZN(n7976) );
  MOAI22 U16906 ( .A1(n29123), .A2(n1035), .B1(ram[3736]), .B2(n1036), 
        .ZN(n7977) );
  MOAI22 U16907 ( .A1(n28888), .A2(n1035), .B1(ram[3737]), .B2(n1036), 
        .ZN(n7978) );
  MOAI22 U16908 ( .A1(n28653), .A2(n1035), .B1(ram[3738]), .B2(n1036), 
        .ZN(n7979) );
  MOAI22 U16909 ( .A1(n28418), .A2(n1035), .B1(ram[3739]), .B2(n1036), 
        .ZN(n7980) );
  MOAI22 U16910 ( .A1(n28183), .A2(n1035), .B1(ram[3740]), .B2(n1036), 
        .ZN(n7981) );
  MOAI22 U16911 ( .A1(n27948), .A2(n1035), .B1(ram[3741]), .B2(n1036), 
        .ZN(n7982) );
  MOAI22 U16912 ( .A1(n27713), .A2(n1035), .B1(ram[3742]), .B2(n1036), 
        .ZN(n7983) );
  MOAI22 U16913 ( .A1(n27478), .A2(n1035), .B1(ram[3743]), .B2(n1036), 
        .ZN(n7984) );
  MOAI22 U16914 ( .A1(n29124), .A2(n1037), .B1(ram[3744]), .B2(n1038), 
        .ZN(n7985) );
  MOAI22 U16915 ( .A1(n28889), .A2(n1037), .B1(ram[3745]), .B2(n1038), 
        .ZN(n7986) );
  MOAI22 U16916 ( .A1(n28654), .A2(n1037), .B1(ram[3746]), .B2(n1038), 
        .ZN(n7987) );
  MOAI22 U16917 ( .A1(n28419), .A2(n1037), .B1(ram[3747]), .B2(n1038), 
        .ZN(n7988) );
  MOAI22 U16918 ( .A1(n28184), .A2(n1037), .B1(ram[3748]), .B2(n1038), 
        .ZN(n7989) );
  MOAI22 U16919 ( .A1(n27949), .A2(n1037), .B1(ram[3749]), .B2(n1038), 
        .ZN(n7990) );
  MOAI22 U16920 ( .A1(n27714), .A2(n1037), .B1(ram[3750]), .B2(n1038), 
        .ZN(n7991) );
  MOAI22 U16921 ( .A1(n27479), .A2(n1037), .B1(ram[3751]), .B2(n1038), 
        .ZN(n7992) );
  MOAI22 U16922 ( .A1(n29124), .A2(n1039), .B1(ram[3752]), .B2(n1040), 
        .ZN(n7993) );
  MOAI22 U16923 ( .A1(n28889), .A2(n1039), .B1(ram[3753]), .B2(n1040), 
        .ZN(n7994) );
  MOAI22 U16924 ( .A1(n28654), .A2(n1039), .B1(ram[3754]), .B2(n1040), 
        .ZN(n7995) );
  MOAI22 U16925 ( .A1(n28419), .A2(n1039), .B1(ram[3755]), .B2(n1040), 
        .ZN(n7996) );
  MOAI22 U16926 ( .A1(n28184), .A2(n1039), .B1(ram[3756]), .B2(n1040), 
        .ZN(n7997) );
  MOAI22 U16927 ( .A1(n27949), .A2(n1039), .B1(ram[3757]), .B2(n1040), 
        .ZN(n7998) );
  MOAI22 U16928 ( .A1(n27714), .A2(n1039), .B1(ram[3758]), .B2(n1040), 
        .ZN(n7999) );
  MOAI22 U16929 ( .A1(n27479), .A2(n1039), .B1(ram[3759]), .B2(n1040), 
        .ZN(n8000) );
  MOAI22 U16930 ( .A1(n29124), .A2(n1041), .B1(ram[3760]), .B2(n1042), 
        .ZN(n8001) );
  MOAI22 U16931 ( .A1(n28889), .A2(n1041), .B1(ram[3761]), .B2(n1042), 
        .ZN(n8002) );
  MOAI22 U16932 ( .A1(n28654), .A2(n1041), .B1(ram[3762]), .B2(n1042), 
        .ZN(n8003) );
  MOAI22 U16933 ( .A1(n28419), .A2(n1041), .B1(ram[3763]), .B2(n1042), 
        .ZN(n8004) );
  MOAI22 U16934 ( .A1(n28184), .A2(n1041), .B1(ram[3764]), .B2(n1042), 
        .ZN(n8005) );
  MOAI22 U16935 ( .A1(n27949), .A2(n1041), .B1(ram[3765]), .B2(n1042), 
        .ZN(n8006) );
  MOAI22 U16936 ( .A1(n27714), .A2(n1041), .B1(ram[3766]), .B2(n1042), 
        .ZN(n8007) );
  MOAI22 U16937 ( .A1(n27479), .A2(n1041), .B1(ram[3767]), .B2(n1042), 
        .ZN(n8008) );
  MOAI22 U16938 ( .A1(n29124), .A2(n1043), .B1(ram[3768]), .B2(n1044), 
        .ZN(n8009) );
  MOAI22 U16939 ( .A1(n28889), .A2(n1043), .B1(ram[3769]), .B2(n1044), 
        .ZN(n8010) );
  MOAI22 U16940 ( .A1(n28654), .A2(n1043), .B1(ram[3770]), .B2(n1044), 
        .ZN(n8011) );
  MOAI22 U16941 ( .A1(n28419), .A2(n1043), .B1(ram[3771]), .B2(n1044), 
        .ZN(n8012) );
  MOAI22 U16942 ( .A1(n28184), .A2(n1043), .B1(ram[3772]), .B2(n1044), 
        .ZN(n8013) );
  MOAI22 U16943 ( .A1(n27949), .A2(n1043), .B1(ram[3773]), .B2(n1044), 
        .ZN(n8014) );
  MOAI22 U16944 ( .A1(n27714), .A2(n1043), .B1(ram[3774]), .B2(n1044), 
        .ZN(n8015) );
  MOAI22 U16945 ( .A1(n27479), .A2(n1043), .B1(ram[3775]), .B2(n1044), 
        .ZN(n8016) );
  MOAI22 U16946 ( .A1(n29124), .A2(n1045), .B1(ram[3776]), .B2(n1046), 
        .ZN(n8017) );
  MOAI22 U16947 ( .A1(n28889), .A2(n1045), .B1(ram[3777]), .B2(n1046), 
        .ZN(n8018) );
  MOAI22 U16948 ( .A1(n28654), .A2(n1045), .B1(ram[3778]), .B2(n1046), 
        .ZN(n8019) );
  MOAI22 U16949 ( .A1(n28419), .A2(n1045), .B1(ram[3779]), .B2(n1046), 
        .ZN(n8020) );
  MOAI22 U16950 ( .A1(n28184), .A2(n1045), .B1(ram[3780]), .B2(n1046), 
        .ZN(n8021) );
  MOAI22 U16951 ( .A1(n27949), .A2(n1045), .B1(ram[3781]), .B2(n1046), 
        .ZN(n8022) );
  MOAI22 U16952 ( .A1(n27714), .A2(n1045), .B1(ram[3782]), .B2(n1046), 
        .ZN(n8023) );
  MOAI22 U16953 ( .A1(n27479), .A2(n1045), .B1(ram[3783]), .B2(n1046), 
        .ZN(n8024) );
  MOAI22 U16954 ( .A1(n29124), .A2(n1047), .B1(ram[3784]), .B2(n1048), 
        .ZN(n8025) );
  MOAI22 U16955 ( .A1(n28889), .A2(n1047), .B1(ram[3785]), .B2(n1048), 
        .ZN(n8026) );
  MOAI22 U16956 ( .A1(n28654), .A2(n1047), .B1(ram[3786]), .B2(n1048), 
        .ZN(n8027) );
  MOAI22 U16957 ( .A1(n28419), .A2(n1047), .B1(ram[3787]), .B2(n1048), 
        .ZN(n8028) );
  MOAI22 U16958 ( .A1(n28184), .A2(n1047), .B1(ram[3788]), .B2(n1048), 
        .ZN(n8029) );
  MOAI22 U16959 ( .A1(n27949), .A2(n1047), .B1(ram[3789]), .B2(n1048), 
        .ZN(n8030) );
  MOAI22 U16960 ( .A1(n27714), .A2(n1047), .B1(ram[3790]), .B2(n1048), 
        .ZN(n8031) );
  MOAI22 U16961 ( .A1(n27479), .A2(n1047), .B1(ram[3791]), .B2(n1048), 
        .ZN(n8032) );
  MOAI22 U16962 ( .A1(n29124), .A2(n1049), .B1(ram[3792]), .B2(n1050), 
        .ZN(n8033) );
  MOAI22 U16963 ( .A1(n28889), .A2(n1049), .B1(ram[3793]), .B2(n1050), 
        .ZN(n8034) );
  MOAI22 U16964 ( .A1(n28654), .A2(n1049), .B1(ram[3794]), .B2(n1050), 
        .ZN(n8035) );
  MOAI22 U16965 ( .A1(n28419), .A2(n1049), .B1(ram[3795]), .B2(n1050), 
        .ZN(n8036) );
  MOAI22 U16966 ( .A1(n28184), .A2(n1049), .B1(ram[3796]), .B2(n1050), 
        .ZN(n8037) );
  MOAI22 U16967 ( .A1(n27949), .A2(n1049), .B1(ram[3797]), .B2(n1050), 
        .ZN(n8038) );
  MOAI22 U16968 ( .A1(n27714), .A2(n1049), .B1(ram[3798]), .B2(n1050), 
        .ZN(n8039) );
  MOAI22 U16969 ( .A1(n27479), .A2(n1049), .B1(ram[3799]), .B2(n1050), 
        .ZN(n8040) );
  MOAI22 U16970 ( .A1(n29124), .A2(n1051), .B1(ram[3800]), .B2(n1052), 
        .ZN(n8041) );
  MOAI22 U16971 ( .A1(n28889), .A2(n1051), .B1(ram[3801]), .B2(n1052), 
        .ZN(n8042) );
  MOAI22 U16972 ( .A1(n28654), .A2(n1051), .B1(ram[3802]), .B2(n1052), 
        .ZN(n8043) );
  MOAI22 U16973 ( .A1(n28419), .A2(n1051), .B1(ram[3803]), .B2(n1052), 
        .ZN(n8044) );
  MOAI22 U16974 ( .A1(n28184), .A2(n1051), .B1(ram[3804]), .B2(n1052), 
        .ZN(n8045) );
  MOAI22 U16975 ( .A1(n27949), .A2(n1051), .B1(ram[3805]), .B2(n1052), 
        .ZN(n8046) );
  MOAI22 U16976 ( .A1(n27714), .A2(n1051), .B1(ram[3806]), .B2(n1052), 
        .ZN(n8047) );
  MOAI22 U16977 ( .A1(n27479), .A2(n1051), .B1(ram[3807]), .B2(n1052), 
        .ZN(n8048) );
  MOAI22 U16978 ( .A1(n29124), .A2(n1053), .B1(ram[3808]), .B2(n1054), 
        .ZN(n8049) );
  MOAI22 U16979 ( .A1(n28889), .A2(n1053), .B1(ram[3809]), .B2(n1054), 
        .ZN(n8050) );
  MOAI22 U16980 ( .A1(n28654), .A2(n1053), .B1(ram[3810]), .B2(n1054), 
        .ZN(n8051) );
  MOAI22 U16981 ( .A1(n28419), .A2(n1053), .B1(ram[3811]), .B2(n1054), 
        .ZN(n8052) );
  MOAI22 U16982 ( .A1(n28184), .A2(n1053), .B1(ram[3812]), .B2(n1054), 
        .ZN(n8053) );
  MOAI22 U16983 ( .A1(n27949), .A2(n1053), .B1(ram[3813]), .B2(n1054), 
        .ZN(n8054) );
  MOAI22 U16984 ( .A1(n27714), .A2(n1053), .B1(ram[3814]), .B2(n1054), 
        .ZN(n8055) );
  MOAI22 U16985 ( .A1(n27479), .A2(n1053), .B1(ram[3815]), .B2(n1054), 
        .ZN(n8056) );
  MOAI22 U16986 ( .A1(n29124), .A2(n1055), .B1(ram[3816]), .B2(n1056), 
        .ZN(n8057) );
  MOAI22 U16987 ( .A1(n28889), .A2(n1055), .B1(ram[3817]), .B2(n1056), 
        .ZN(n8058) );
  MOAI22 U16988 ( .A1(n28654), .A2(n1055), .B1(ram[3818]), .B2(n1056), 
        .ZN(n8059) );
  MOAI22 U16989 ( .A1(n28419), .A2(n1055), .B1(ram[3819]), .B2(n1056), 
        .ZN(n8060) );
  MOAI22 U16990 ( .A1(n28184), .A2(n1055), .B1(ram[3820]), .B2(n1056), 
        .ZN(n8061) );
  MOAI22 U16991 ( .A1(n27949), .A2(n1055), .B1(ram[3821]), .B2(n1056), 
        .ZN(n8062) );
  MOAI22 U16992 ( .A1(n27714), .A2(n1055), .B1(ram[3822]), .B2(n1056), 
        .ZN(n8063) );
  MOAI22 U16993 ( .A1(n27479), .A2(n1055), .B1(ram[3823]), .B2(n1056), 
        .ZN(n8064) );
  MOAI22 U16994 ( .A1(n29124), .A2(n1057), .B1(ram[3824]), .B2(n1058), 
        .ZN(n8065) );
  MOAI22 U16995 ( .A1(n28889), .A2(n1057), .B1(ram[3825]), .B2(n1058), 
        .ZN(n8066) );
  MOAI22 U16996 ( .A1(n28654), .A2(n1057), .B1(ram[3826]), .B2(n1058), 
        .ZN(n8067) );
  MOAI22 U16997 ( .A1(n28419), .A2(n1057), .B1(ram[3827]), .B2(n1058), 
        .ZN(n8068) );
  MOAI22 U16998 ( .A1(n28184), .A2(n1057), .B1(ram[3828]), .B2(n1058), 
        .ZN(n8069) );
  MOAI22 U16999 ( .A1(n27949), .A2(n1057), .B1(ram[3829]), .B2(n1058), 
        .ZN(n8070) );
  MOAI22 U17000 ( .A1(n27714), .A2(n1057), .B1(ram[3830]), .B2(n1058), 
        .ZN(n8071) );
  MOAI22 U17001 ( .A1(n27479), .A2(n1057), .B1(ram[3831]), .B2(n1058), 
        .ZN(n8072) );
  MOAI22 U17002 ( .A1(n29124), .A2(n1059), .B1(ram[3832]), .B2(n1060), 
        .ZN(n8073) );
  MOAI22 U17003 ( .A1(n28889), .A2(n1059), .B1(ram[3833]), .B2(n1060), 
        .ZN(n8074) );
  MOAI22 U17004 ( .A1(n28654), .A2(n1059), .B1(ram[3834]), .B2(n1060), 
        .ZN(n8075) );
  MOAI22 U17005 ( .A1(n28419), .A2(n1059), .B1(ram[3835]), .B2(n1060), 
        .ZN(n8076) );
  MOAI22 U17006 ( .A1(n28184), .A2(n1059), .B1(ram[3836]), .B2(n1060), 
        .ZN(n8077) );
  MOAI22 U17007 ( .A1(n27949), .A2(n1059), .B1(ram[3837]), .B2(n1060), 
        .ZN(n8078) );
  MOAI22 U17008 ( .A1(n27714), .A2(n1059), .B1(ram[3838]), .B2(n1060), 
        .ZN(n8079) );
  MOAI22 U17009 ( .A1(n27479), .A2(n1059), .B1(ram[3839]), .B2(n1060), 
        .ZN(n8080) );
  MOAI22 U17010 ( .A1(n29124), .A2(n1061), .B1(ram[3840]), .B2(n1062), 
        .ZN(n8081) );
  MOAI22 U17011 ( .A1(n28889), .A2(n1061), .B1(ram[3841]), .B2(n1062), 
        .ZN(n8082) );
  MOAI22 U17012 ( .A1(n28654), .A2(n1061), .B1(ram[3842]), .B2(n1062), 
        .ZN(n8083) );
  MOAI22 U17013 ( .A1(n28419), .A2(n1061), .B1(ram[3843]), .B2(n1062), 
        .ZN(n8084) );
  MOAI22 U17014 ( .A1(n28184), .A2(n1061), .B1(ram[3844]), .B2(n1062), 
        .ZN(n8085) );
  MOAI22 U17015 ( .A1(n27949), .A2(n1061), .B1(ram[3845]), .B2(n1062), 
        .ZN(n8086) );
  MOAI22 U17016 ( .A1(n27714), .A2(n1061), .B1(ram[3846]), .B2(n1062), 
        .ZN(n8087) );
  MOAI22 U17017 ( .A1(n27479), .A2(n1061), .B1(ram[3847]), .B2(n1062), 
        .ZN(n8088) );
  MOAI22 U17018 ( .A1(n29125), .A2(n1063), .B1(ram[3848]), .B2(n1064), 
        .ZN(n8089) );
  MOAI22 U17019 ( .A1(n28890), .A2(n1063), .B1(ram[3849]), .B2(n1064), 
        .ZN(n8090) );
  MOAI22 U17020 ( .A1(n28655), .A2(n1063), .B1(ram[3850]), .B2(n1064), 
        .ZN(n8091) );
  MOAI22 U17021 ( .A1(n28420), .A2(n1063), .B1(ram[3851]), .B2(n1064), 
        .ZN(n8092) );
  MOAI22 U17022 ( .A1(n28185), .A2(n1063), .B1(ram[3852]), .B2(n1064), 
        .ZN(n8093) );
  MOAI22 U17023 ( .A1(n27950), .A2(n1063), .B1(ram[3853]), .B2(n1064), 
        .ZN(n8094) );
  MOAI22 U17024 ( .A1(n27715), .A2(n1063), .B1(ram[3854]), .B2(n1064), 
        .ZN(n8095) );
  MOAI22 U17025 ( .A1(n27480), .A2(n1063), .B1(ram[3855]), .B2(n1064), 
        .ZN(n8096) );
  MOAI22 U17026 ( .A1(n29125), .A2(n1065), .B1(ram[3856]), .B2(n1066), 
        .ZN(n8097) );
  MOAI22 U17027 ( .A1(n28890), .A2(n1065), .B1(ram[3857]), .B2(n1066), 
        .ZN(n8098) );
  MOAI22 U17028 ( .A1(n28655), .A2(n1065), .B1(ram[3858]), .B2(n1066), 
        .ZN(n8099) );
  MOAI22 U17029 ( .A1(n28420), .A2(n1065), .B1(ram[3859]), .B2(n1066), 
        .ZN(n8100) );
  MOAI22 U17030 ( .A1(n28185), .A2(n1065), .B1(ram[3860]), .B2(n1066), 
        .ZN(n8101) );
  MOAI22 U17031 ( .A1(n27950), .A2(n1065), .B1(ram[3861]), .B2(n1066), 
        .ZN(n8102) );
  MOAI22 U17032 ( .A1(n27715), .A2(n1065), .B1(ram[3862]), .B2(n1066), 
        .ZN(n8103) );
  MOAI22 U17033 ( .A1(n27480), .A2(n1065), .B1(ram[3863]), .B2(n1066), 
        .ZN(n8104) );
  MOAI22 U17034 ( .A1(n29125), .A2(n1067), .B1(ram[3864]), .B2(n1068), 
        .ZN(n8105) );
  MOAI22 U17035 ( .A1(n28890), .A2(n1067), .B1(ram[3865]), .B2(n1068), 
        .ZN(n8106) );
  MOAI22 U17036 ( .A1(n28655), .A2(n1067), .B1(ram[3866]), .B2(n1068), 
        .ZN(n8107) );
  MOAI22 U17037 ( .A1(n28420), .A2(n1067), .B1(ram[3867]), .B2(n1068), 
        .ZN(n8108) );
  MOAI22 U17038 ( .A1(n28185), .A2(n1067), .B1(ram[3868]), .B2(n1068), 
        .ZN(n8109) );
  MOAI22 U17039 ( .A1(n27950), .A2(n1067), .B1(ram[3869]), .B2(n1068), 
        .ZN(n8110) );
  MOAI22 U17040 ( .A1(n27715), .A2(n1067), .B1(ram[3870]), .B2(n1068), 
        .ZN(n8111) );
  MOAI22 U17041 ( .A1(n27480), .A2(n1067), .B1(ram[3871]), .B2(n1068), 
        .ZN(n8112) );
  MOAI22 U17042 ( .A1(n29125), .A2(n1069), .B1(ram[3872]), .B2(n1070), 
        .ZN(n8113) );
  MOAI22 U17043 ( .A1(n28890), .A2(n1069), .B1(ram[3873]), .B2(n1070), 
        .ZN(n8114) );
  MOAI22 U17044 ( .A1(n28655), .A2(n1069), .B1(ram[3874]), .B2(n1070), 
        .ZN(n8115) );
  MOAI22 U17045 ( .A1(n28420), .A2(n1069), .B1(ram[3875]), .B2(n1070), 
        .ZN(n8116) );
  MOAI22 U17046 ( .A1(n28185), .A2(n1069), .B1(ram[3876]), .B2(n1070), 
        .ZN(n8117) );
  MOAI22 U17047 ( .A1(n27950), .A2(n1069), .B1(ram[3877]), .B2(n1070), 
        .ZN(n8118) );
  MOAI22 U17048 ( .A1(n27715), .A2(n1069), .B1(ram[3878]), .B2(n1070), 
        .ZN(n8119) );
  MOAI22 U17049 ( .A1(n27480), .A2(n1069), .B1(ram[3879]), .B2(n1070), 
        .ZN(n8120) );
  MOAI22 U17050 ( .A1(n29125), .A2(n1071), .B1(ram[3880]), .B2(n1072), 
        .ZN(n8121) );
  MOAI22 U17051 ( .A1(n28890), .A2(n1071), .B1(ram[3881]), .B2(n1072), 
        .ZN(n8122) );
  MOAI22 U17052 ( .A1(n28655), .A2(n1071), .B1(ram[3882]), .B2(n1072), 
        .ZN(n8123) );
  MOAI22 U17053 ( .A1(n28420), .A2(n1071), .B1(ram[3883]), .B2(n1072), 
        .ZN(n8124) );
  MOAI22 U17054 ( .A1(n28185), .A2(n1071), .B1(ram[3884]), .B2(n1072), 
        .ZN(n8125) );
  MOAI22 U17055 ( .A1(n27950), .A2(n1071), .B1(ram[3885]), .B2(n1072), 
        .ZN(n8126) );
  MOAI22 U17056 ( .A1(n27715), .A2(n1071), .B1(ram[3886]), .B2(n1072), 
        .ZN(n8127) );
  MOAI22 U17057 ( .A1(n27480), .A2(n1071), .B1(ram[3887]), .B2(n1072), 
        .ZN(n8128) );
  MOAI22 U17058 ( .A1(n29125), .A2(n1073), .B1(ram[3888]), .B2(n1074), 
        .ZN(n8129) );
  MOAI22 U17059 ( .A1(n28890), .A2(n1073), .B1(ram[3889]), .B2(n1074), 
        .ZN(n8130) );
  MOAI22 U17060 ( .A1(n28655), .A2(n1073), .B1(ram[3890]), .B2(n1074), 
        .ZN(n8131) );
  MOAI22 U17061 ( .A1(n28420), .A2(n1073), .B1(ram[3891]), .B2(n1074), 
        .ZN(n8132) );
  MOAI22 U17062 ( .A1(n28185), .A2(n1073), .B1(ram[3892]), .B2(n1074), 
        .ZN(n8133) );
  MOAI22 U17063 ( .A1(n27950), .A2(n1073), .B1(ram[3893]), .B2(n1074), 
        .ZN(n8134) );
  MOAI22 U17064 ( .A1(n27715), .A2(n1073), .B1(ram[3894]), .B2(n1074), 
        .ZN(n8135) );
  MOAI22 U17065 ( .A1(n27480), .A2(n1073), .B1(ram[3895]), .B2(n1074), 
        .ZN(n8136) );
  MOAI22 U17066 ( .A1(n29125), .A2(n1075), .B1(ram[3896]), .B2(n1076), 
        .ZN(n8137) );
  MOAI22 U17067 ( .A1(n28890), .A2(n1075), .B1(ram[3897]), .B2(n1076), 
        .ZN(n8138) );
  MOAI22 U17068 ( .A1(n28655), .A2(n1075), .B1(ram[3898]), .B2(n1076), 
        .ZN(n8139) );
  MOAI22 U17069 ( .A1(n28420), .A2(n1075), .B1(ram[3899]), .B2(n1076), 
        .ZN(n8140) );
  MOAI22 U17070 ( .A1(n28185), .A2(n1075), .B1(ram[3900]), .B2(n1076), 
        .ZN(n8141) );
  MOAI22 U17071 ( .A1(n27950), .A2(n1075), .B1(ram[3901]), .B2(n1076), 
        .ZN(n8142) );
  MOAI22 U17072 ( .A1(n27715), .A2(n1075), .B1(ram[3902]), .B2(n1076), 
        .ZN(n8143) );
  MOAI22 U17073 ( .A1(n27480), .A2(n1075), .B1(ram[3903]), .B2(n1076), 
        .ZN(n8144) );
  MOAI22 U17074 ( .A1(n29125), .A2(n1077), .B1(ram[3904]), .B2(n1078), 
        .ZN(n8145) );
  MOAI22 U17075 ( .A1(n28890), .A2(n1077), .B1(ram[3905]), .B2(n1078), 
        .ZN(n8146) );
  MOAI22 U17076 ( .A1(n28655), .A2(n1077), .B1(ram[3906]), .B2(n1078), 
        .ZN(n8147) );
  MOAI22 U17077 ( .A1(n28420), .A2(n1077), .B1(ram[3907]), .B2(n1078), 
        .ZN(n8148) );
  MOAI22 U17078 ( .A1(n28185), .A2(n1077), .B1(ram[3908]), .B2(n1078), 
        .ZN(n8149) );
  MOAI22 U17079 ( .A1(n27950), .A2(n1077), .B1(ram[3909]), .B2(n1078), 
        .ZN(n8150) );
  MOAI22 U17080 ( .A1(n27715), .A2(n1077), .B1(ram[3910]), .B2(n1078), 
        .ZN(n8151) );
  MOAI22 U17081 ( .A1(n27480), .A2(n1077), .B1(ram[3911]), .B2(n1078), 
        .ZN(n8152) );
  MOAI22 U17082 ( .A1(n29125), .A2(n1079), .B1(ram[3912]), .B2(n1080), 
        .ZN(n8153) );
  MOAI22 U17083 ( .A1(n28890), .A2(n1079), .B1(ram[3913]), .B2(n1080), 
        .ZN(n8154) );
  MOAI22 U17084 ( .A1(n28655), .A2(n1079), .B1(ram[3914]), .B2(n1080), 
        .ZN(n8155) );
  MOAI22 U17085 ( .A1(n28420), .A2(n1079), .B1(ram[3915]), .B2(n1080), 
        .ZN(n8156) );
  MOAI22 U17086 ( .A1(n28185), .A2(n1079), .B1(ram[3916]), .B2(n1080), 
        .ZN(n8157) );
  MOAI22 U17087 ( .A1(n27950), .A2(n1079), .B1(ram[3917]), .B2(n1080), 
        .ZN(n8158) );
  MOAI22 U17088 ( .A1(n27715), .A2(n1079), .B1(ram[3918]), .B2(n1080), 
        .ZN(n8159) );
  MOAI22 U17089 ( .A1(n27480), .A2(n1079), .B1(ram[3919]), .B2(n1080), 
        .ZN(n8160) );
  MOAI22 U17090 ( .A1(n29125), .A2(n1081), .B1(ram[3920]), .B2(n1082), 
        .ZN(n8161) );
  MOAI22 U17091 ( .A1(n28890), .A2(n1081), .B1(ram[3921]), .B2(n1082), 
        .ZN(n8162) );
  MOAI22 U17092 ( .A1(n28655), .A2(n1081), .B1(ram[3922]), .B2(n1082), 
        .ZN(n8163) );
  MOAI22 U17093 ( .A1(n28420), .A2(n1081), .B1(ram[3923]), .B2(n1082), 
        .ZN(n8164) );
  MOAI22 U17094 ( .A1(n28185), .A2(n1081), .B1(ram[3924]), .B2(n1082), 
        .ZN(n8165) );
  MOAI22 U17095 ( .A1(n27950), .A2(n1081), .B1(ram[3925]), .B2(n1082), 
        .ZN(n8166) );
  MOAI22 U17096 ( .A1(n27715), .A2(n1081), .B1(ram[3926]), .B2(n1082), 
        .ZN(n8167) );
  MOAI22 U17097 ( .A1(n27480), .A2(n1081), .B1(ram[3927]), .B2(n1082), 
        .ZN(n8168) );
  MOAI22 U17098 ( .A1(n29125), .A2(n1083), .B1(ram[3928]), .B2(n1084), 
        .ZN(n8169) );
  MOAI22 U17099 ( .A1(n28890), .A2(n1083), .B1(ram[3929]), .B2(n1084), 
        .ZN(n8170) );
  MOAI22 U17100 ( .A1(n28655), .A2(n1083), .B1(ram[3930]), .B2(n1084), 
        .ZN(n8171) );
  MOAI22 U17101 ( .A1(n28420), .A2(n1083), .B1(ram[3931]), .B2(n1084), 
        .ZN(n8172) );
  MOAI22 U17102 ( .A1(n28185), .A2(n1083), .B1(ram[3932]), .B2(n1084), 
        .ZN(n8173) );
  MOAI22 U17103 ( .A1(n27950), .A2(n1083), .B1(ram[3933]), .B2(n1084), 
        .ZN(n8174) );
  MOAI22 U17104 ( .A1(n27715), .A2(n1083), .B1(ram[3934]), .B2(n1084), 
        .ZN(n8175) );
  MOAI22 U17105 ( .A1(n27480), .A2(n1083), .B1(ram[3935]), .B2(n1084), 
        .ZN(n8176) );
  MOAI22 U17106 ( .A1(n29125), .A2(n1085), .B1(ram[3936]), .B2(n1086), 
        .ZN(n8177) );
  MOAI22 U17107 ( .A1(n28890), .A2(n1085), .B1(ram[3937]), .B2(n1086), 
        .ZN(n8178) );
  MOAI22 U17108 ( .A1(n28655), .A2(n1085), .B1(ram[3938]), .B2(n1086), 
        .ZN(n8179) );
  MOAI22 U17109 ( .A1(n28420), .A2(n1085), .B1(ram[3939]), .B2(n1086), 
        .ZN(n8180) );
  MOAI22 U17110 ( .A1(n28185), .A2(n1085), .B1(ram[3940]), .B2(n1086), 
        .ZN(n8181) );
  MOAI22 U17111 ( .A1(n27950), .A2(n1085), .B1(ram[3941]), .B2(n1086), 
        .ZN(n8182) );
  MOAI22 U17112 ( .A1(n27715), .A2(n1085), .B1(ram[3942]), .B2(n1086), 
        .ZN(n8183) );
  MOAI22 U17113 ( .A1(n27480), .A2(n1085), .B1(ram[3943]), .B2(n1086), 
        .ZN(n8184) );
  MOAI22 U17114 ( .A1(n29125), .A2(n1087), .B1(ram[3944]), .B2(n1088), 
        .ZN(n8185) );
  MOAI22 U17115 ( .A1(n28890), .A2(n1087), .B1(ram[3945]), .B2(n1088), 
        .ZN(n8186) );
  MOAI22 U17116 ( .A1(n28655), .A2(n1087), .B1(ram[3946]), .B2(n1088), 
        .ZN(n8187) );
  MOAI22 U17117 ( .A1(n28420), .A2(n1087), .B1(ram[3947]), .B2(n1088), 
        .ZN(n8188) );
  MOAI22 U17118 ( .A1(n28185), .A2(n1087), .B1(ram[3948]), .B2(n1088), 
        .ZN(n8189) );
  MOAI22 U17119 ( .A1(n27950), .A2(n1087), .B1(ram[3949]), .B2(n1088), 
        .ZN(n8190) );
  MOAI22 U17120 ( .A1(n27715), .A2(n1087), .B1(ram[3950]), .B2(n1088), 
        .ZN(n8191) );
  MOAI22 U17121 ( .A1(n27480), .A2(n1087), .B1(ram[3951]), .B2(n1088), 
        .ZN(n8192) );
  MOAI22 U17122 ( .A1(n29126), .A2(n1089), .B1(ram[3952]), .B2(n1090), 
        .ZN(n8193) );
  MOAI22 U17123 ( .A1(n28891), .A2(n1089), .B1(ram[3953]), .B2(n1090), 
        .ZN(n8194) );
  MOAI22 U17124 ( .A1(n28656), .A2(n1089), .B1(ram[3954]), .B2(n1090), 
        .ZN(n8195) );
  MOAI22 U17125 ( .A1(n28421), .A2(n1089), .B1(ram[3955]), .B2(n1090), 
        .ZN(n8196) );
  MOAI22 U17126 ( .A1(n28186), .A2(n1089), .B1(ram[3956]), .B2(n1090), 
        .ZN(n8197) );
  MOAI22 U17127 ( .A1(n27951), .A2(n1089), .B1(ram[3957]), .B2(n1090), 
        .ZN(n8198) );
  MOAI22 U17128 ( .A1(n27716), .A2(n1089), .B1(ram[3958]), .B2(n1090), 
        .ZN(n8199) );
  MOAI22 U17129 ( .A1(n27481), .A2(n1089), .B1(ram[3959]), .B2(n1090), 
        .ZN(n8200) );
  MOAI22 U17130 ( .A1(n29126), .A2(n1091), .B1(ram[3960]), .B2(n1092), 
        .ZN(n8201) );
  MOAI22 U17131 ( .A1(n28891), .A2(n1091), .B1(ram[3961]), .B2(n1092), 
        .ZN(n8202) );
  MOAI22 U17132 ( .A1(n28656), .A2(n1091), .B1(ram[3962]), .B2(n1092), 
        .ZN(n8203) );
  MOAI22 U17133 ( .A1(n28421), .A2(n1091), .B1(ram[3963]), .B2(n1092), 
        .ZN(n8204) );
  MOAI22 U17134 ( .A1(n28186), .A2(n1091), .B1(ram[3964]), .B2(n1092), 
        .ZN(n8205) );
  MOAI22 U17135 ( .A1(n27951), .A2(n1091), .B1(ram[3965]), .B2(n1092), 
        .ZN(n8206) );
  MOAI22 U17136 ( .A1(n27716), .A2(n1091), .B1(ram[3966]), .B2(n1092), 
        .ZN(n8207) );
  MOAI22 U17137 ( .A1(n27481), .A2(n1091), .B1(ram[3967]), .B2(n1092), 
        .ZN(n8208) );
  MOAI22 U17138 ( .A1(n29126), .A2(n1093), .B1(ram[3968]), .B2(n1094), 
        .ZN(n8209) );
  MOAI22 U17139 ( .A1(n28891), .A2(n1093), .B1(ram[3969]), .B2(n1094), 
        .ZN(n8210) );
  MOAI22 U17140 ( .A1(n28656), .A2(n1093), .B1(ram[3970]), .B2(n1094), 
        .ZN(n8211) );
  MOAI22 U17141 ( .A1(n28421), .A2(n1093), .B1(ram[3971]), .B2(n1094), 
        .ZN(n8212) );
  MOAI22 U17142 ( .A1(n28186), .A2(n1093), .B1(ram[3972]), .B2(n1094), 
        .ZN(n8213) );
  MOAI22 U17143 ( .A1(n27951), .A2(n1093), .B1(ram[3973]), .B2(n1094), 
        .ZN(n8214) );
  MOAI22 U17144 ( .A1(n27716), .A2(n1093), .B1(ram[3974]), .B2(n1094), 
        .ZN(n8215) );
  MOAI22 U17145 ( .A1(n27481), .A2(n1093), .B1(ram[3975]), .B2(n1094), 
        .ZN(n8216) );
  MOAI22 U17146 ( .A1(n29126), .A2(n1095), .B1(ram[3976]), .B2(n1096), 
        .ZN(n8217) );
  MOAI22 U17147 ( .A1(n28891), .A2(n1095), .B1(ram[3977]), .B2(n1096), 
        .ZN(n8218) );
  MOAI22 U17148 ( .A1(n28656), .A2(n1095), .B1(ram[3978]), .B2(n1096), 
        .ZN(n8219) );
  MOAI22 U17149 ( .A1(n28421), .A2(n1095), .B1(ram[3979]), .B2(n1096), 
        .ZN(n8220) );
  MOAI22 U17150 ( .A1(n28186), .A2(n1095), .B1(ram[3980]), .B2(n1096), 
        .ZN(n8221) );
  MOAI22 U17151 ( .A1(n27951), .A2(n1095), .B1(ram[3981]), .B2(n1096), 
        .ZN(n8222) );
  MOAI22 U17152 ( .A1(n27716), .A2(n1095), .B1(ram[3982]), .B2(n1096), 
        .ZN(n8223) );
  MOAI22 U17153 ( .A1(n27481), .A2(n1095), .B1(ram[3983]), .B2(n1096), 
        .ZN(n8224) );
  MOAI22 U17154 ( .A1(n29126), .A2(n1097), .B1(ram[3984]), .B2(n1098), 
        .ZN(n8225) );
  MOAI22 U17155 ( .A1(n28891), .A2(n1097), .B1(ram[3985]), .B2(n1098), 
        .ZN(n8226) );
  MOAI22 U17156 ( .A1(n28656), .A2(n1097), .B1(ram[3986]), .B2(n1098), 
        .ZN(n8227) );
  MOAI22 U17157 ( .A1(n28421), .A2(n1097), .B1(ram[3987]), .B2(n1098), 
        .ZN(n8228) );
  MOAI22 U17158 ( .A1(n28186), .A2(n1097), .B1(ram[3988]), .B2(n1098), 
        .ZN(n8229) );
  MOAI22 U17159 ( .A1(n27951), .A2(n1097), .B1(ram[3989]), .B2(n1098), 
        .ZN(n8230) );
  MOAI22 U17160 ( .A1(n27716), .A2(n1097), .B1(ram[3990]), .B2(n1098), 
        .ZN(n8231) );
  MOAI22 U17161 ( .A1(n27481), .A2(n1097), .B1(ram[3991]), .B2(n1098), 
        .ZN(n8232) );
  MOAI22 U17162 ( .A1(n29126), .A2(n1099), .B1(ram[3992]), .B2(n1100), 
        .ZN(n8233) );
  MOAI22 U17163 ( .A1(n28891), .A2(n1099), .B1(ram[3993]), .B2(n1100), 
        .ZN(n8234) );
  MOAI22 U17164 ( .A1(n28656), .A2(n1099), .B1(ram[3994]), .B2(n1100), 
        .ZN(n8235) );
  MOAI22 U17165 ( .A1(n28421), .A2(n1099), .B1(ram[3995]), .B2(n1100), 
        .ZN(n8236) );
  MOAI22 U17166 ( .A1(n28186), .A2(n1099), .B1(ram[3996]), .B2(n1100), 
        .ZN(n8237) );
  MOAI22 U17167 ( .A1(n27951), .A2(n1099), .B1(ram[3997]), .B2(n1100), 
        .ZN(n8238) );
  MOAI22 U17168 ( .A1(n27716), .A2(n1099), .B1(ram[3998]), .B2(n1100), 
        .ZN(n8239) );
  MOAI22 U17169 ( .A1(n27481), .A2(n1099), .B1(ram[3999]), .B2(n1100), 
        .ZN(n8240) );
  MOAI22 U17170 ( .A1(n29126), .A2(n1101), .B1(ram[4000]), .B2(n1102), 
        .ZN(n8241) );
  MOAI22 U17171 ( .A1(n28891), .A2(n1101), .B1(ram[4001]), .B2(n1102), 
        .ZN(n8242) );
  MOAI22 U17172 ( .A1(n28656), .A2(n1101), .B1(ram[4002]), .B2(n1102), 
        .ZN(n8243) );
  MOAI22 U17173 ( .A1(n28421), .A2(n1101), .B1(ram[4003]), .B2(n1102), 
        .ZN(n8244) );
  MOAI22 U17174 ( .A1(n28186), .A2(n1101), .B1(ram[4004]), .B2(n1102), 
        .ZN(n8245) );
  MOAI22 U17175 ( .A1(n27951), .A2(n1101), .B1(ram[4005]), .B2(n1102), 
        .ZN(n8246) );
  MOAI22 U17176 ( .A1(n27716), .A2(n1101), .B1(ram[4006]), .B2(n1102), 
        .ZN(n8247) );
  MOAI22 U17177 ( .A1(n27481), .A2(n1101), .B1(ram[4007]), .B2(n1102), 
        .ZN(n8248) );
  MOAI22 U17178 ( .A1(n29126), .A2(n1103), .B1(ram[4008]), .B2(n1104), 
        .ZN(n8249) );
  MOAI22 U17179 ( .A1(n28891), .A2(n1103), .B1(ram[4009]), .B2(n1104), 
        .ZN(n8250) );
  MOAI22 U17180 ( .A1(n28656), .A2(n1103), .B1(ram[4010]), .B2(n1104), 
        .ZN(n8251) );
  MOAI22 U17181 ( .A1(n28421), .A2(n1103), .B1(ram[4011]), .B2(n1104), 
        .ZN(n8252) );
  MOAI22 U17182 ( .A1(n28186), .A2(n1103), .B1(ram[4012]), .B2(n1104), 
        .ZN(n8253) );
  MOAI22 U17183 ( .A1(n27951), .A2(n1103), .B1(ram[4013]), .B2(n1104), 
        .ZN(n8254) );
  MOAI22 U17184 ( .A1(n27716), .A2(n1103), .B1(ram[4014]), .B2(n1104), 
        .ZN(n8255) );
  MOAI22 U17185 ( .A1(n27481), .A2(n1103), .B1(ram[4015]), .B2(n1104), 
        .ZN(n8256) );
  MOAI22 U17186 ( .A1(n29126), .A2(n1105), .B1(ram[4016]), .B2(n1106), 
        .ZN(n8257) );
  MOAI22 U17187 ( .A1(n28891), .A2(n1105), .B1(ram[4017]), .B2(n1106), 
        .ZN(n8258) );
  MOAI22 U17188 ( .A1(n28656), .A2(n1105), .B1(ram[4018]), .B2(n1106), 
        .ZN(n8259) );
  MOAI22 U17189 ( .A1(n28421), .A2(n1105), .B1(ram[4019]), .B2(n1106), 
        .ZN(n8260) );
  MOAI22 U17190 ( .A1(n28186), .A2(n1105), .B1(ram[4020]), .B2(n1106), 
        .ZN(n8261) );
  MOAI22 U17191 ( .A1(n27951), .A2(n1105), .B1(ram[4021]), .B2(n1106), 
        .ZN(n8262) );
  MOAI22 U17192 ( .A1(n27716), .A2(n1105), .B1(ram[4022]), .B2(n1106), 
        .ZN(n8263) );
  MOAI22 U17193 ( .A1(n27481), .A2(n1105), .B1(ram[4023]), .B2(n1106), 
        .ZN(n8264) );
  MOAI22 U17194 ( .A1(n29126), .A2(n1107), .B1(ram[4024]), .B2(n1108), 
        .ZN(n8265) );
  MOAI22 U17195 ( .A1(n28891), .A2(n1107), .B1(ram[4025]), .B2(n1108), 
        .ZN(n8266) );
  MOAI22 U17196 ( .A1(n28656), .A2(n1107), .B1(ram[4026]), .B2(n1108), 
        .ZN(n8267) );
  MOAI22 U17197 ( .A1(n28421), .A2(n1107), .B1(ram[4027]), .B2(n1108), 
        .ZN(n8268) );
  MOAI22 U17198 ( .A1(n28186), .A2(n1107), .B1(ram[4028]), .B2(n1108), 
        .ZN(n8269) );
  MOAI22 U17199 ( .A1(n27951), .A2(n1107), .B1(ram[4029]), .B2(n1108), 
        .ZN(n8270) );
  MOAI22 U17200 ( .A1(n27716), .A2(n1107), .B1(ram[4030]), .B2(n1108), 
        .ZN(n8271) );
  MOAI22 U17201 ( .A1(n27481), .A2(n1107), .B1(ram[4031]), .B2(n1108), 
        .ZN(n8272) );
  MOAI22 U17202 ( .A1(n29126), .A2(n1109), .B1(ram[4032]), .B2(n1110), 
        .ZN(n8273) );
  MOAI22 U17203 ( .A1(n28891), .A2(n1109), .B1(ram[4033]), .B2(n1110), 
        .ZN(n8274) );
  MOAI22 U17204 ( .A1(n28656), .A2(n1109), .B1(ram[4034]), .B2(n1110), 
        .ZN(n8275) );
  MOAI22 U17205 ( .A1(n28421), .A2(n1109), .B1(ram[4035]), .B2(n1110), 
        .ZN(n8276) );
  MOAI22 U17206 ( .A1(n28186), .A2(n1109), .B1(ram[4036]), .B2(n1110), 
        .ZN(n8277) );
  MOAI22 U17207 ( .A1(n27951), .A2(n1109), .B1(ram[4037]), .B2(n1110), 
        .ZN(n8278) );
  MOAI22 U17208 ( .A1(n27716), .A2(n1109), .B1(ram[4038]), .B2(n1110), 
        .ZN(n8279) );
  MOAI22 U17209 ( .A1(n27481), .A2(n1109), .B1(ram[4039]), .B2(n1110), 
        .ZN(n8280) );
  MOAI22 U17210 ( .A1(n29126), .A2(n1111), .B1(ram[4040]), .B2(n1112), 
        .ZN(n8281) );
  MOAI22 U17211 ( .A1(n28891), .A2(n1111), .B1(ram[4041]), .B2(n1112), 
        .ZN(n8282) );
  MOAI22 U17212 ( .A1(n28656), .A2(n1111), .B1(ram[4042]), .B2(n1112), 
        .ZN(n8283) );
  MOAI22 U17213 ( .A1(n28421), .A2(n1111), .B1(ram[4043]), .B2(n1112), 
        .ZN(n8284) );
  MOAI22 U17214 ( .A1(n28186), .A2(n1111), .B1(ram[4044]), .B2(n1112), 
        .ZN(n8285) );
  MOAI22 U17215 ( .A1(n27951), .A2(n1111), .B1(ram[4045]), .B2(n1112), 
        .ZN(n8286) );
  MOAI22 U17216 ( .A1(n27716), .A2(n1111), .B1(ram[4046]), .B2(n1112), 
        .ZN(n8287) );
  MOAI22 U17217 ( .A1(n27481), .A2(n1111), .B1(ram[4047]), .B2(n1112), 
        .ZN(n8288) );
  MOAI22 U17218 ( .A1(n29126), .A2(n1113), .B1(ram[4048]), .B2(n1114), 
        .ZN(n8289) );
  MOAI22 U17219 ( .A1(n28891), .A2(n1113), .B1(ram[4049]), .B2(n1114), 
        .ZN(n8290) );
  MOAI22 U17220 ( .A1(n28656), .A2(n1113), .B1(ram[4050]), .B2(n1114), 
        .ZN(n8291) );
  MOAI22 U17221 ( .A1(n28421), .A2(n1113), .B1(ram[4051]), .B2(n1114), 
        .ZN(n8292) );
  MOAI22 U17222 ( .A1(n28186), .A2(n1113), .B1(ram[4052]), .B2(n1114), 
        .ZN(n8293) );
  MOAI22 U17223 ( .A1(n27951), .A2(n1113), .B1(ram[4053]), .B2(n1114), 
        .ZN(n8294) );
  MOAI22 U17224 ( .A1(n27716), .A2(n1113), .B1(ram[4054]), .B2(n1114), 
        .ZN(n8295) );
  MOAI22 U17225 ( .A1(n27481), .A2(n1113), .B1(ram[4055]), .B2(n1114), 
        .ZN(n8296) );
  MOAI22 U17226 ( .A1(n29127), .A2(n1115), .B1(ram[4056]), .B2(n1116), 
        .ZN(n8297) );
  MOAI22 U17227 ( .A1(n28892), .A2(n1115), .B1(ram[4057]), .B2(n1116), 
        .ZN(n8298) );
  MOAI22 U17228 ( .A1(n28657), .A2(n1115), .B1(ram[4058]), .B2(n1116), 
        .ZN(n8299) );
  MOAI22 U17229 ( .A1(n28422), .A2(n1115), .B1(ram[4059]), .B2(n1116), 
        .ZN(n8300) );
  MOAI22 U17230 ( .A1(n28187), .A2(n1115), .B1(ram[4060]), .B2(n1116), 
        .ZN(n8301) );
  MOAI22 U17231 ( .A1(n27952), .A2(n1115), .B1(ram[4061]), .B2(n1116), 
        .ZN(n8302) );
  MOAI22 U17232 ( .A1(n27717), .A2(n1115), .B1(ram[4062]), .B2(n1116), 
        .ZN(n8303) );
  MOAI22 U17233 ( .A1(n27482), .A2(n1115), .B1(ram[4063]), .B2(n1116), 
        .ZN(n8304) );
  MOAI22 U17234 ( .A1(n29127), .A2(n1117), .B1(ram[4064]), .B2(n1118), 
        .ZN(n8305) );
  MOAI22 U17235 ( .A1(n28892), .A2(n1117), .B1(ram[4065]), .B2(n1118), 
        .ZN(n8306) );
  MOAI22 U17236 ( .A1(n28657), .A2(n1117), .B1(ram[4066]), .B2(n1118), 
        .ZN(n8307) );
  MOAI22 U17237 ( .A1(n28422), .A2(n1117), .B1(ram[4067]), .B2(n1118), 
        .ZN(n8308) );
  MOAI22 U17238 ( .A1(n28187), .A2(n1117), .B1(ram[4068]), .B2(n1118), 
        .ZN(n8309) );
  MOAI22 U17239 ( .A1(n27952), .A2(n1117), .B1(ram[4069]), .B2(n1118), 
        .ZN(n8310) );
  MOAI22 U17240 ( .A1(n27717), .A2(n1117), .B1(ram[4070]), .B2(n1118), 
        .ZN(n8311) );
  MOAI22 U17241 ( .A1(n27482), .A2(n1117), .B1(ram[4071]), .B2(n1118), 
        .ZN(n8312) );
  MOAI22 U17242 ( .A1(n29127), .A2(n1119), .B1(ram[4072]), .B2(n1120), 
        .ZN(n8313) );
  MOAI22 U17243 ( .A1(n28892), .A2(n1119), .B1(ram[4073]), .B2(n1120), 
        .ZN(n8314) );
  MOAI22 U17244 ( .A1(n28657), .A2(n1119), .B1(ram[4074]), .B2(n1120), 
        .ZN(n8315) );
  MOAI22 U17245 ( .A1(n28422), .A2(n1119), .B1(ram[4075]), .B2(n1120), 
        .ZN(n8316) );
  MOAI22 U17246 ( .A1(n28187), .A2(n1119), .B1(ram[4076]), .B2(n1120), 
        .ZN(n8317) );
  MOAI22 U17247 ( .A1(n27952), .A2(n1119), .B1(ram[4077]), .B2(n1120), 
        .ZN(n8318) );
  MOAI22 U17248 ( .A1(n27717), .A2(n1119), .B1(ram[4078]), .B2(n1120), 
        .ZN(n8319) );
  MOAI22 U17249 ( .A1(n27482), .A2(n1119), .B1(ram[4079]), .B2(n1120), 
        .ZN(n8320) );
  MOAI22 U17250 ( .A1(n29127), .A2(n1121), .B1(ram[4080]), .B2(n1122), 
        .ZN(n8321) );
  MOAI22 U17251 ( .A1(n28892), .A2(n1121), .B1(ram[4081]), .B2(n1122), 
        .ZN(n8322) );
  MOAI22 U17252 ( .A1(n28657), .A2(n1121), .B1(ram[4082]), .B2(n1122), 
        .ZN(n8323) );
  MOAI22 U17253 ( .A1(n28422), .A2(n1121), .B1(ram[4083]), .B2(n1122), 
        .ZN(n8324) );
  MOAI22 U17254 ( .A1(n28187), .A2(n1121), .B1(ram[4084]), .B2(n1122), 
        .ZN(n8325) );
  MOAI22 U17255 ( .A1(n27952), .A2(n1121), .B1(ram[4085]), .B2(n1122), 
        .ZN(n8326) );
  MOAI22 U17256 ( .A1(n27717), .A2(n1121), .B1(ram[4086]), .B2(n1122), 
        .ZN(n8327) );
  MOAI22 U17257 ( .A1(n27482), .A2(n1121), .B1(ram[4087]), .B2(n1122), 
        .ZN(n8328) );
  MOAI22 U17258 ( .A1(n29127), .A2(n1126), .B1(ram[4096]), .B2(n1127), 
        .ZN(n8337) );
  MOAI22 U17259 ( .A1(n28892), .A2(n1126), .B1(ram[4097]), .B2(n1127), 
        .ZN(n8338) );
  MOAI22 U17260 ( .A1(n28657), .A2(n1126), .B1(ram[4098]), .B2(n1127), 
        .ZN(n8339) );
  MOAI22 U17261 ( .A1(n28422), .A2(n1126), .B1(ram[4099]), .B2(n1127), 
        .ZN(n8340) );
  MOAI22 U17262 ( .A1(n28187), .A2(n1126), .B1(ram[4100]), .B2(n1127), 
        .ZN(n8341) );
  MOAI22 U17263 ( .A1(n27952), .A2(n1126), .B1(ram[4101]), .B2(n1127), 
        .ZN(n8342) );
  MOAI22 U17264 ( .A1(n27717), .A2(n1126), .B1(ram[4102]), .B2(n1127), 
        .ZN(n8343) );
  MOAI22 U17265 ( .A1(n27482), .A2(n1126), .B1(ram[4103]), .B2(n1127), 
        .ZN(n8344) );
  MOAI22 U17266 ( .A1(n29127), .A2(n1129), .B1(ram[4104]), .B2(n1130), 
        .ZN(n8345) );
  MOAI22 U17267 ( .A1(n28892), .A2(n1129), .B1(ram[4105]), .B2(n1130), 
        .ZN(n8346) );
  MOAI22 U17268 ( .A1(n28657), .A2(n1129), .B1(ram[4106]), .B2(n1130), 
        .ZN(n8347) );
  MOAI22 U17269 ( .A1(n28422), .A2(n1129), .B1(ram[4107]), .B2(n1130), 
        .ZN(n8348) );
  MOAI22 U17270 ( .A1(n28187), .A2(n1129), .B1(ram[4108]), .B2(n1130), 
        .ZN(n8349) );
  MOAI22 U17271 ( .A1(n27952), .A2(n1129), .B1(ram[4109]), .B2(n1130), 
        .ZN(n8350) );
  MOAI22 U17272 ( .A1(n27717), .A2(n1129), .B1(ram[4110]), .B2(n1130), 
        .ZN(n8351) );
  MOAI22 U17273 ( .A1(n27482), .A2(n1129), .B1(ram[4111]), .B2(n1130), 
        .ZN(n8352) );
  MOAI22 U17274 ( .A1(n29127), .A2(n1131), .B1(ram[4112]), .B2(n1132), 
        .ZN(n8353) );
  MOAI22 U17275 ( .A1(n28892), .A2(n1131), .B1(ram[4113]), .B2(n1132), 
        .ZN(n8354) );
  MOAI22 U17276 ( .A1(n28657), .A2(n1131), .B1(ram[4114]), .B2(n1132), 
        .ZN(n8355) );
  MOAI22 U17277 ( .A1(n28422), .A2(n1131), .B1(ram[4115]), .B2(n1132), 
        .ZN(n8356) );
  MOAI22 U17278 ( .A1(n28187), .A2(n1131), .B1(ram[4116]), .B2(n1132), 
        .ZN(n8357) );
  MOAI22 U17279 ( .A1(n27952), .A2(n1131), .B1(ram[4117]), .B2(n1132), 
        .ZN(n8358) );
  MOAI22 U17280 ( .A1(n27717), .A2(n1131), .B1(ram[4118]), .B2(n1132), 
        .ZN(n8359) );
  MOAI22 U17281 ( .A1(n27482), .A2(n1131), .B1(ram[4119]), .B2(n1132), 
        .ZN(n8360) );
  MOAI22 U17282 ( .A1(n29127), .A2(n1133), .B1(ram[4120]), .B2(n1134), 
        .ZN(n8361) );
  MOAI22 U17283 ( .A1(n28892), .A2(n1133), .B1(ram[4121]), .B2(n1134), 
        .ZN(n8362) );
  MOAI22 U17284 ( .A1(n28657), .A2(n1133), .B1(ram[4122]), .B2(n1134), 
        .ZN(n8363) );
  MOAI22 U17285 ( .A1(n28422), .A2(n1133), .B1(ram[4123]), .B2(n1134), 
        .ZN(n8364) );
  MOAI22 U17286 ( .A1(n28187), .A2(n1133), .B1(ram[4124]), .B2(n1134), 
        .ZN(n8365) );
  MOAI22 U17287 ( .A1(n27952), .A2(n1133), .B1(ram[4125]), .B2(n1134), 
        .ZN(n8366) );
  MOAI22 U17288 ( .A1(n27717), .A2(n1133), .B1(ram[4126]), .B2(n1134), 
        .ZN(n8367) );
  MOAI22 U17289 ( .A1(n27482), .A2(n1133), .B1(ram[4127]), .B2(n1134), 
        .ZN(n8368) );
  MOAI22 U17290 ( .A1(n29127), .A2(n1135), .B1(ram[4128]), .B2(n1136), 
        .ZN(n8369) );
  MOAI22 U17291 ( .A1(n28892), .A2(n1135), .B1(ram[4129]), .B2(n1136), 
        .ZN(n8370) );
  MOAI22 U17292 ( .A1(n28657), .A2(n1135), .B1(ram[4130]), .B2(n1136), 
        .ZN(n8371) );
  MOAI22 U17293 ( .A1(n28422), .A2(n1135), .B1(ram[4131]), .B2(n1136), 
        .ZN(n8372) );
  MOAI22 U17294 ( .A1(n28187), .A2(n1135), .B1(ram[4132]), .B2(n1136), 
        .ZN(n8373) );
  MOAI22 U17295 ( .A1(n27952), .A2(n1135), .B1(ram[4133]), .B2(n1136), 
        .ZN(n8374) );
  MOAI22 U17296 ( .A1(n27717), .A2(n1135), .B1(ram[4134]), .B2(n1136), 
        .ZN(n8375) );
  MOAI22 U17297 ( .A1(n27482), .A2(n1135), .B1(ram[4135]), .B2(n1136), 
        .ZN(n8376) );
  MOAI22 U17298 ( .A1(n29127), .A2(n1137), .B1(ram[4136]), .B2(n1138), 
        .ZN(n8377) );
  MOAI22 U17299 ( .A1(n28892), .A2(n1137), .B1(ram[4137]), .B2(n1138), 
        .ZN(n8378) );
  MOAI22 U17300 ( .A1(n28657), .A2(n1137), .B1(ram[4138]), .B2(n1138), 
        .ZN(n8379) );
  MOAI22 U17301 ( .A1(n28422), .A2(n1137), .B1(ram[4139]), .B2(n1138), 
        .ZN(n8380) );
  MOAI22 U17302 ( .A1(n28187), .A2(n1137), .B1(ram[4140]), .B2(n1138), 
        .ZN(n8381) );
  MOAI22 U17303 ( .A1(n27952), .A2(n1137), .B1(ram[4141]), .B2(n1138), 
        .ZN(n8382) );
  MOAI22 U17304 ( .A1(n27717), .A2(n1137), .B1(ram[4142]), .B2(n1138), 
        .ZN(n8383) );
  MOAI22 U17305 ( .A1(n27482), .A2(n1137), .B1(ram[4143]), .B2(n1138), 
        .ZN(n8384) );
  MOAI22 U17306 ( .A1(n29127), .A2(n1139), .B1(ram[4144]), .B2(n1140), 
        .ZN(n8385) );
  MOAI22 U17307 ( .A1(n28892), .A2(n1139), .B1(ram[4145]), .B2(n1140), 
        .ZN(n8386) );
  MOAI22 U17308 ( .A1(n28657), .A2(n1139), .B1(ram[4146]), .B2(n1140), 
        .ZN(n8387) );
  MOAI22 U17309 ( .A1(n28422), .A2(n1139), .B1(ram[4147]), .B2(n1140), 
        .ZN(n8388) );
  MOAI22 U17310 ( .A1(n28187), .A2(n1139), .B1(ram[4148]), .B2(n1140), 
        .ZN(n8389) );
  MOAI22 U17311 ( .A1(n27952), .A2(n1139), .B1(ram[4149]), .B2(n1140), 
        .ZN(n8390) );
  MOAI22 U17312 ( .A1(n27717), .A2(n1139), .B1(ram[4150]), .B2(n1140), 
        .ZN(n8391) );
  MOAI22 U17313 ( .A1(n27482), .A2(n1139), .B1(ram[4151]), .B2(n1140), 
        .ZN(n8392) );
  MOAI22 U17314 ( .A1(n29127), .A2(n1141), .B1(ram[4152]), .B2(n1142), 
        .ZN(n8393) );
  MOAI22 U17315 ( .A1(n28892), .A2(n1141), .B1(ram[4153]), .B2(n1142), 
        .ZN(n8394) );
  MOAI22 U17316 ( .A1(n28657), .A2(n1141), .B1(ram[4154]), .B2(n1142), 
        .ZN(n8395) );
  MOAI22 U17317 ( .A1(n28422), .A2(n1141), .B1(ram[4155]), .B2(n1142), 
        .ZN(n8396) );
  MOAI22 U17318 ( .A1(n28187), .A2(n1141), .B1(ram[4156]), .B2(n1142), 
        .ZN(n8397) );
  MOAI22 U17319 ( .A1(n27952), .A2(n1141), .B1(ram[4157]), .B2(n1142), 
        .ZN(n8398) );
  MOAI22 U17320 ( .A1(n27717), .A2(n1141), .B1(ram[4158]), .B2(n1142), 
        .ZN(n8399) );
  MOAI22 U17321 ( .A1(n27482), .A2(n1141), .B1(ram[4159]), .B2(n1142), 
        .ZN(n8400) );
  MOAI22 U17322 ( .A1(n29128), .A2(n1143), .B1(ram[4160]), .B2(n1144), 
        .ZN(n8401) );
  MOAI22 U17323 ( .A1(n28893), .A2(n1143), .B1(ram[4161]), .B2(n1144), 
        .ZN(n8402) );
  MOAI22 U17324 ( .A1(n28658), .A2(n1143), .B1(ram[4162]), .B2(n1144), 
        .ZN(n8403) );
  MOAI22 U17325 ( .A1(n28423), .A2(n1143), .B1(ram[4163]), .B2(n1144), 
        .ZN(n8404) );
  MOAI22 U17326 ( .A1(n28188), .A2(n1143), .B1(ram[4164]), .B2(n1144), 
        .ZN(n8405) );
  MOAI22 U17327 ( .A1(n27953), .A2(n1143), .B1(ram[4165]), .B2(n1144), 
        .ZN(n8406) );
  MOAI22 U17328 ( .A1(n27718), .A2(n1143), .B1(ram[4166]), .B2(n1144), 
        .ZN(n8407) );
  MOAI22 U17329 ( .A1(n27483), .A2(n1143), .B1(ram[4167]), .B2(n1144), 
        .ZN(n8408) );
  MOAI22 U17330 ( .A1(n29128), .A2(n1145), .B1(ram[4168]), .B2(n1146), 
        .ZN(n8409) );
  MOAI22 U17331 ( .A1(n28893), .A2(n1145), .B1(ram[4169]), .B2(n1146), 
        .ZN(n8410) );
  MOAI22 U17332 ( .A1(n28658), .A2(n1145), .B1(ram[4170]), .B2(n1146), 
        .ZN(n8411) );
  MOAI22 U17333 ( .A1(n28423), .A2(n1145), .B1(ram[4171]), .B2(n1146), 
        .ZN(n8412) );
  MOAI22 U17334 ( .A1(n28188), .A2(n1145), .B1(ram[4172]), .B2(n1146), 
        .ZN(n8413) );
  MOAI22 U17335 ( .A1(n27953), .A2(n1145), .B1(ram[4173]), .B2(n1146), 
        .ZN(n8414) );
  MOAI22 U17336 ( .A1(n27718), .A2(n1145), .B1(ram[4174]), .B2(n1146), 
        .ZN(n8415) );
  MOAI22 U17337 ( .A1(n27483), .A2(n1145), .B1(ram[4175]), .B2(n1146), 
        .ZN(n8416) );
  MOAI22 U17338 ( .A1(n29128), .A2(n1147), .B1(ram[4176]), .B2(n1148), 
        .ZN(n8417) );
  MOAI22 U17339 ( .A1(n28893), .A2(n1147), .B1(ram[4177]), .B2(n1148), 
        .ZN(n8418) );
  MOAI22 U17340 ( .A1(n28658), .A2(n1147), .B1(ram[4178]), .B2(n1148), 
        .ZN(n8419) );
  MOAI22 U17341 ( .A1(n28423), .A2(n1147), .B1(ram[4179]), .B2(n1148), 
        .ZN(n8420) );
  MOAI22 U17342 ( .A1(n28188), .A2(n1147), .B1(ram[4180]), .B2(n1148), 
        .ZN(n8421) );
  MOAI22 U17343 ( .A1(n27953), .A2(n1147), .B1(ram[4181]), .B2(n1148), 
        .ZN(n8422) );
  MOAI22 U17344 ( .A1(n27718), .A2(n1147), .B1(ram[4182]), .B2(n1148), 
        .ZN(n8423) );
  MOAI22 U17345 ( .A1(n27483), .A2(n1147), .B1(ram[4183]), .B2(n1148), 
        .ZN(n8424) );
  MOAI22 U17346 ( .A1(n29128), .A2(n1149), .B1(ram[4184]), .B2(n1150), 
        .ZN(n8425) );
  MOAI22 U17347 ( .A1(n28893), .A2(n1149), .B1(ram[4185]), .B2(n1150), 
        .ZN(n8426) );
  MOAI22 U17348 ( .A1(n28658), .A2(n1149), .B1(ram[4186]), .B2(n1150), 
        .ZN(n8427) );
  MOAI22 U17349 ( .A1(n28423), .A2(n1149), .B1(ram[4187]), .B2(n1150), 
        .ZN(n8428) );
  MOAI22 U17350 ( .A1(n28188), .A2(n1149), .B1(ram[4188]), .B2(n1150), 
        .ZN(n8429) );
  MOAI22 U17351 ( .A1(n27953), .A2(n1149), .B1(ram[4189]), .B2(n1150), 
        .ZN(n8430) );
  MOAI22 U17352 ( .A1(n27718), .A2(n1149), .B1(ram[4190]), .B2(n1150), 
        .ZN(n8431) );
  MOAI22 U17353 ( .A1(n27483), .A2(n1149), .B1(ram[4191]), .B2(n1150), 
        .ZN(n8432) );
  MOAI22 U17354 ( .A1(n29128), .A2(n1151), .B1(ram[4192]), .B2(n1152), 
        .ZN(n8433) );
  MOAI22 U17355 ( .A1(n28893), .A2(n1151), .B1(ram[4193]), .B2(n1152), 
        .ZN(n8434) );
  MOAI22 U17356 ( .A1(n28658), .A2(n1151), .B1(ram[4194]), .B2(n1152), 
        .ZN(n8435) );
  MOAI22 U17357 ( .A1(n28423), .A2(n1151), .B1(ram[4195]), .B2(n1152), 
        .ZN(n8436) );
  MOAI22 U17358 ( .A1(n28188), .A2(n1151), .B1(ram[4196]), .B2(n1152), 
        .ZN(n8437) );
  MOAI22 U17359 ( .A1(n27953), .A2(n1151), .B1(ram[4197]), .B2(n1152), 
        .ZN(n8438) );
  MOAI22 U17360 ( .A1(n27718), .A2(n1151), .B1(ram[4198]), .B2(n1152), 
        .ZN(n8439) );
  MOAI22 U17361 ( .A1(n27483), .A2(n1151), .B1(ram[4199]), .B2(n1152), 
        .ZN(n8440) );
  MOAI22 U17362 ( .A1(n29128), .A2(n1153), .B1(ram[4200]), .B2(n1154), 
        .ZN(n8441) );
  MOAI22 U17363 ( .A1(n28893), .A2(n1153), .B1(ram[4201]), .B2(n1154), 
        .ZN(n8442) );
  MOAI22 U17364 ( .A1(n28658), .A2(n1153), .B1(ram[4202]), .B2(n1154), 
        .ZN(n8443) );
  MOAI22 U17365 ( .A1(n28423), .A2(n1153), .B1(ram[4203]), .B2(n1154), 
        .ZN(n8444) );
  MOAI22 U17366 ( .A1(n28188), .A2(n1153), .B1(ram[4204]), .B2(n1154), 
        .ZN(n8445) );
  MOAI22 U17367 ( .A1(n27953), .A2(n1153), .B1(ram[4205]), .B2(n1154), 
        .ZN(n8446) );
  MOAI22 U17368 ( .A1(n27718), .A2(n1153), .B1(ram[4206]), .B2(n1154), 
        .ZN(n8447) );
  MOAI22 U17369 ( .A1(n27483), .A2(n1153), .B1(ram[4207]), .B2(n1154), 
        .ZN(n8448) );
  MOAI22 U17370 ( .A1(n29128), .A2(n1155), .B1(ram[4208]), .B2(n1156), 
        .ZN(n8449) );
  MOAI22 U17371 ( .A1(n28893), .A2(n1155), .B1(ram[4209]), .B2(n1156), 
        .ZN(n8450) );
  MOAI22 U17372 ( .A1(n28658), .A2(n1155), .B1(ram[4210]), .B2(n1156), 
        .ZN(n8451) );
  MOAI22 U17373 ( .A1(n28423), .A2(n1155), .B1(ram[4211]), .B2(n1156), 
        .ZN(n8452) );
  MOAI22 U17374 ( .A1(n28188), .A2(n1155), .B1(ram[4212]), .B2(n1156), 
        .ZN(n8453) );
  MOAI22 U17375 ( .A1(n27953), .A2(n1155), .B1(ram[4213]), .B2(n1156), 
        .ZN(n8454) );
  MOAI22 U17376 ( .A1(n27718), .A2(n1155), .B1(ram[4214]), .B2(n1156), 
        .ZN(n8455) );
  MOAI22 U17377 ( .A1(n27483), .A2(n1155), .B1(ram[4215]), .B2(n1156), 
        .ZN(n8456) );
  MOAI22 U17378 ( .A1(n29128), .A2(n1157), .B1(ram[4216]), .B2(n1158), 
        .ZN(n8457) );
  MOAI22 U17379 ( .A1(n28893), .A2(n1157), .B1(ram[4217]), .B2(n1158), 
        .ZN(n8458) );
  MOAI22 U17380 ( .A1(n28658), .A2(n1157), .B1(ram[4218]), .B2(n1158), 
        .ZN(n8459) );
  MOAI22 U17381 ( .A1(n28423), .A2(n1157), .B1(ram[4219]), .B2(n1158), 
        .ZN(n8460) );
  MOAI22 U17382 ( .A1(n28188), .A2(n1157), .B1(ram[4220]), .B2(n1158), 
        .ZN(n8461) );
  MOAI22 U17383 ( .A1(n27953), .A2(n1157), .B1(ram[4221]), .B2(n1158), 
        .ZN(n8462) );
  MOAI22 U17384 ( .A1(n27718), .A2(n1157), .B1(ram[4222]), .B2(n1158), 
        .ZN(n8463) );
  MOAI22 U17385 ( .A1(n27483), .A2(n1157), .B1(ram[4223]), .B2(n1158), 
        .ZN(n8464) );
  MOAI22 U17386 ( .A1(n29128), .A2(n1159), .B1(ram[4224]), .B2(n1160), 
        .ZN(n8465) );
  MOAI22 U17387 ( .A1(n28893), .A2(n1159), .B1(ram[4225]), .B2(n1160), 
        .ZN(n8466) );
  MOAI22 U17388 ( .A1(n28658), .A2(n1159), .B1(ram[4226]), .B2(n1160), 
        .ZN(n8467) );
  MOAI22 U17389 ( .A1(n28423), .A2(n1159), .B1(ram[4227]), .B2(n1160), 
        .ZN(n8468) );
  MOAI22 U17390 ( .A1(n28188), .A2(n1159), .B1(ram[4228]), .B2(n1160), 
        .ZN(n8469) );
  MOAI22 U17391 ( .A1(n27953), .A2(n1159), .B1(ram[4229]), .B2(n1160), 
        .ZN(n8470) );
  MOAI22 U17392 ( .A1(n27718), .A2(n1159), .B1(ram[4230]), .B2(n1160), 
        .ZN(n8471) );
  MOAI22 U17393 ( .A1(n27483), .A2(n1159), .B1(ram[4231]), .B2(n1160), 
        .ZN(n8472) );
  MOAI22 U17394 ( .A1(n29128), .A2(n1161), .B1(ram[4232]), .B2(n1162), 
        .ZN(n8473) );
  MOAI22 U17395 ( .A1(n28893), .A2(n1161), .B1(ram[4233]), .B2(n1162), 
        .ZN(n8474) );
  MOAI22 U17396 ( .A1(n28658), .A2(n1161), .B1(ram[4234]), .B2(n1162), 
        .ZN(n8475) );
  MOAI22 U17397 ( .A1(n28423), .A2(n1161), .B1(ram[4235]), .B2(n1162), 
        .ZN(n8476) );
  MOAI22 U17398 ( .A1(n28188), .A2(n1161), .B1(ram[4236]), .B2(n1162), 
        .ZN(n8477) );
  MOAI22 U17399 ( .A1(n27953), .A2(n1161), .B1(ram[4237]), .B2(n1162), 
        .ZN(n8478) );
  MOAI22 U17400 ( .A1(n27718), .A2(n1161), .B1(ram[4238]), .B2(n1162), 
        .ZN(n8479) );
  MOAI22 U17401 ( .A1(n27483), .A2(n1161), .B1(ram[4239]), .B2(n1162), 
        .ZN(n8480) );
  MOAI22 U17402 ( .A1(n29128), .A2(n1163), .B1(ram[4240]), .B2(n1164), 
        .ZN(n8481) );
  MOAI22 U17403 ( .A1(n28893), .A2(n1163), .B1(ram[4241]), .B2(n1164), 
        .ZN(n8482) );
  MOAI22 U17404 ( .A1(n28658), .A2(n1163), .B1(ram[4242]), .B2(n1164), 
        .ZN(n8483) );
  MOAI22 U17405 ( .A1(n28423), .A2(n1163), .B1(ram[4243]), .B2(n1164), 
        .ZN(n8484) );
  MOAI22 U17406 ( .A1(n28188), .A2(n1163), .B1(ram[4244]), .B2(n1164), 
        .ZN(n8485) );
  MOAI22 U17407 ( .A1(n27953), .A2(n1163), .B1(ram[4245]), .B2(n1164), 
        .ZN(n8486) );
  MOAI22 U17408 ( .A1(n27718), .A2(n1163), .B1(ram[4246]), .B2(n1164), 
        .ZN(n8487) );
  MOAI22 U17409 ( .A1(n27483), .A2(n1163), .B1(ram[4247]), .B2(n1164), 
        .ZN(n8488) );
  MOAI22 U17410 ( .A1(n29128), .A2(n1165), .B1(ram[4248]), .B2(n1166), 
        .ZN(n8489) );
  MOAI22 U17411 ( .A1(n28893), .A2(n1165), .B1(ram[4249]), .B2(n1166), 
        .ZN(n8490) );
  MOAI22 U17412 ( .A1(n28658), .A2(n1165), .B1(ram[4250]), .B2(n1166), 
        .ZN(n8491) );
  MOAI22 U17413 ( .A1(n28423), .A2(n1165), .B1(ram[4251]), .B2(n1166), 
        .ZN(n8492) );
  MOAI22 U17414 ( .A1(n28188), .A2(n1165), .B1(ram[4252]), .B2(n1166), 
        .ZN(n8493) );
  MOAI22 U17415 ( .A1(n27953), .A2(n1165), .B1(ram[4253]), .B2(n1166), 
        .ZN(n8494) );
  MOAI22 U17416 ( .A1(n27718), .A2(n1165), .B1(ram[4254]), .B2(n1166), 
        .ZN(n8495) );
  MOAI22 U17417 ( .A1(n27483), .A2(n1165), .B1(ram[4255]), .B2(n1166), 
        .ZN(n8496) );
  MOAI22 U17418 ( .A1(n29128), .A2(n1167), .B1(ram[4256]), .B2(n1168), 
        .ZN(n8497) );
  MOAI22 U17419 ( .A1(n28893), .A2(n1167), .B1(ram[4257]), .B2(n1168), 
        .ZN(n8498) );
  MOAI22 U17420 ( .A1(n28658), .A2(n1167), .B1(ram[4258]), .B2(n1168), 
        .ZN(n8499) );
  MOAI22 U17421 ( .A1(n28423), .A2(n1167), .B1(ram[4259]), .B2(n1168), 
        .ZN(n8500) );
  MOAI22 U17422 ( .A1(n28188), .A2(n1167), .B1(ram[4260]), .B2(n1168), 
        .ZN(n8501) );
  MOAI22 U17423 ( .A1(n27953), .A2(n1167), .B1(ram[4261]), .B2(n1168), 
        .ZN(n8502) );
  MOAI22 U17424 ( .A1(n27718), .A2(n1167), .B1(ram[4262]), .B2(n1168), 
        .ZN(n8503) );
  MOAI22 U17425 ( .A1(n27483), .A2(n1167), .B1(ram[4263]), .B2(n1168), 
        .ZN(n8504) );
  MOAI22 U17426 ( .A1(n29129), .A2(n1169), .B1(ram[4264]), .B2(n1170), 
        .ZN(n8505) );
  MOAI22 U17427 ( .A1(n28894), .A2(n1169), .B1(ram[4265]), .B2(n1170), 
        .ZN(n8506) );
  MOAI22 U17428 ( .A1(n28659), .A2(n1169), .B1(ram[4266]), .B2(n1170), 
        .ZN(n8507) );
  MOAI22 U17429 ( .A1(n28424), .A2(n1169), .B1(ram[4267]), .B2(n1170), 
        .ZN(n8508) );
  MOAI22 U17430 ( .A1(n28189), .A2(n1169), .B1(ram[4268]), .B2(n1170), 
        .ZN(n8509) );
  MOAI22 U17431 ( .A1(n27954), .A2(n1169), .B1(ram[4269]), .B2(n1170), 
        .ZN(n8510) );
  MOAI22 U17432 ( .A1(n27719), .A2(n1169), .B1(ram[4270]), .B2(n1170), 
        .ZN(n8511) );
  MOAI22 U17433 ( .A1(n27484), .A2(n1169), .B1(ram[4271]), .B2(n1170), 
        .ZN(n8512) );
  MOAI22 U17434 ( .A1(n29129), .A2(n1171), .B1(ram[4272]), .B2(n1172), 
        .ZN(n8513) );
  MOAI22 U17435 ( .A1(n28894), .A2(n1171), .B1(ram[4273]), .B2(n1172), 
        .ZN(n8514) );
  MOAI22 U17436 ( .A1(n28659), .A2(n1171), .B1(ram[4274]), .B2(n1172), 
        .ZN(n8515) );
  MOAI22 U17437 ( .A1(n28424), .A2(n1171), .B1(ram[4275]), .B2(n1172), 
        .ZN(n8516) );
  MOAI22 U17438 ( .A1(n28189), .A2(n1171), .B1(ram[4276]), .B2(n1172), 
        .ZN(n8517) );
  MOAI22 U17439 ( .A1(n27954), .A2(n1171), .B1(ram[4277]), .B2(n1172), 
        .ZN(n8518) );
  MOAI22 U17440 ( .A1(n27719), .A2(n1171), .B1(ram[4278]), .B2(n1172), 
        .ZN(n8519) );
  MOAI22 U17441 ( .A1(n27484), .A2(n1171), .B1(ram[4279]), .B2(n1172), 
        .ZN(n8520) );
  MOAI22 U17442 ( .A1(n29129), .A2(n1173), .B1(ram[4280]), .B2(n1174), 
        .ZN(n8521) );
  MOAI22 U17443 ( .A1(n28894), .A2(n1173), .B1(ram[4281]), .B2(n1174), 
        .ZN(n8522) );
  MOAI22 U17444 ( .A1(n28659), .A2(n1173), .B1(ram[4282]), .B2(n1174), 
        .ZN(n8523) );
  MOAI22 U17445 ( .A1(n28424), .A2(n1173), .B1(ram[4283]), .B2(n1174), 
        .ZN(n8524) );
  MOAI22 U17446 ( .A1(n28189), .A2(n1173), .B1(ram[4284]), .B2(n1174), 
        .ZN(n8525) );
  MOAI22 U17447 ( .A1(n27954), .A2(n1173), .B1(ram[4285]), .B2(n1174), 
        .ZN(n8526) );
  MOAI22 U17448 ( .A1(n27719), .A2(n1173), .B1(ram[4286]), .B2(n1174), 
        .ZN(n8527) );
  MOAI22 U17449 ( .A1(n27484), .A2(n1173), .B1(ram[4287]), .B2(n1174), 
        .ZN(n8528) );
  MOAI22 U17450 ( .A1(n29129), .A2(n1175), .B1(ram[4288]), .B2(n1176), 
        .ZN(n8529) );
  MOAI22 U17451 ( .A1(n28894), .A2(n1175), .B1(ram[4289]), .B2(n1176), 
        .ZN(n8530) );
  MOAI22 U17452 ( .A1(n28659), .A2(n1175), .B1(ram[4290]), .B2(n1176), 
        .ZN(n8531) );
  MOAI22 U17453 ( .A1(n28424), .A2(n1175), .B1(ram[4291]), .B2(n1176), 
        .ZN(n8532) );
  MOAI22 U17454 ( .A1(n28189), .A2(n1175), .B1(ram[4292]), .B2(n1176), 
        .ZN(n8533) );
  MOAI22 U17455 ( .A1(n27954), .A2(n1175), .B1(ram[4293]), .B2(n1176), 
        .ZN(n8534) );
  MOAI22 U17456 ( .A1(n27719), .A2(n1175), .B1(ram[4294]), .B2(n1176), 
        .ZN(n8535) );
  MOAI22 U17457 ( .A1(n27484), .A2(n1175), .B1(ram[4295]), .B2(n1176), 
        .ZN(n8536) );
  MOAI22 U17458 ( .A1(n29129), .A2(n1177), .B1(ram[4296]), .B2(n1178), 
        .ZN(n8537) );
  MOAI22 U17459 ( .A1(n28894), .A2(n1177), .B1(ram[4297]), .B2(n1178), 
        .ZN(n8538) );
  MOAI22 U17460 ( .A1(n28659), .A2(n1177), .B1(ram[4298]), .B2(n1178), 
        .ZN(n8539) );
  MOAI22 U17461 ( .A1(n28424), .A2(n1177), .B1(ram[4299]), .B2(n1178), 
        .ZN(n8540) );
  MOAI22 U17462 ( .A1(n28189), .A2(n1177), .B1(ram[4300]), .B2(n1178), 
        .ZN(n8541) );
  MOAI22 U17463 ( .A1(n27954), .A2(n1177), .B1(ram[4301]), .B2(n1178), 
        .ZN(n8542) );
  MOAI22 U17464 ( .A1(n27719), .A2(n1177), .B1(ram[4302]), .B2(n1178), 
        .ZN(n8543) );
  MOAI22 U17465 ( .A1(n27484), .A2(n1177), .B1(ram[4303]), .B2(n1178), 
        .ZN(n8544) );
  MOAI22 U17466 ( .A1(n29129), .A2(n1179), .B1(ram[4304]), .B2(n1180), 
        .ZN(n8545) );
  MOAI22 U17467 ( .A1(n28894), .A2(n1179), .B1(ram[4305]), .B2(n1180), 
        .ZN(n8546) );
  MOAI22 U17468 ( .A1(n28659), .A2(n1179), .B1(ram[4306]), .B2(n1180), 
        .ZN(n8547) );
  MOAI22 U17469 ( .A1(n28424), .A2(n1179), .B1(ram[4307]), .B2(n1180), 
        .ZN(n8548) );
  MOAI22 U17470 ( .A1(n28189), .A2(n1179), .B1(ram[4308]), .B2(n1180), 
        .ZN(n8549) );
  MOAI22 U17471 ( .A1(n27954), .A2(n1179), .B1(ram[4309]), .B2(n1180), 
        .ZN(n8550) );
  MOAI22 U17472 ( .A1(n27719), .A2(n1179), .B1(ram[4310]), .B2(n1180), 
        .ZN(n8551) );
  MOAI22 U17473 ( .A1(n27484), .A2(n1179), .B1(ram[4311]), .B2(n1180), 
        .ZN(n8552) );
  MOAI22 U17474 ( .A1(n29129), .A2(n1181), .B1(ram[4312]), .B2(n1182), 
        .ZN(n8553) );
  MOAI22 U17475 ( .A1(n28894), .A2(n1181), .B1(ram[4313]), .B2(n1182), 
        .ZN(n8554) );
  MOAI22 U17476 ( .A1(n28659), .A2(n1181), .B1(ram[4314]), .B2(n1182), 
        .ZN(n8555) );
  MOAI22 U17477 ( .A1(n28424), .A2(n1181), .B1(ram[4315]), .B2(n1182), 
        .ZN(n8556) );
  MOAI22 U17478 ( .A1(n28189), .A2(n1181), .B1(ram[4316]), .B2(n1182), 
        .ZN(n8557) );
  MOAI22 U17479 ( .A1(n27954), .A2(n1181), .B1(ram[4317]), .B2(n1182), 
        .ZN(n8558) );
  MOAI22 U17480 ( .A1(n27719), .A2(n1181), .B1(ram[4318]), .B2(n1182), 
        .ZN(n8559) );
  MOAI22 U17481 ( .A1(n27484), .A2(n1181), .B1(ram[4319]), .B2(n1182), 
        .ZN(n8560) );
  MOAI22 U17482 ( .A1(n29129), .A2(n1183), .B1(ram[4320]), .B2(n1184), 
        .ZN(n8561) );
  MOAI22 U17483 ( .A1(n28894), .A2(n1183), .B1(ram[4321]), .B2(n1184), 
        .ZN(n8562) );
  MOAI22 U17484 ( .A1(n28659), .A2(n1183), .B1(ram[4322]), .B2(n1184), 
        .ZN(n8563) );
  MOAI22 U17485 ( .A1(n28424), .A2(n1183), .B1(ram[4323]), .B2(n1184), 
        .ZN(n8564) );
  MOAI22 U17486 ( .A1(n28189), .A2(n1183), .B1(ram[4324]), .B2(n1184), 
        .ZN(n8565) );
  MOAI22 U17487 ( .A1(n27954), .A2(n1183), .B1(ram[4325]), .B2(n1184), 
        .ZN(n8566) );
  MOAI22 U17488 ( .A1(n27719), .A2(n1183), .B1(ram[4326]), .B2(n1184), 
        .ZN(n8567) );
  MOAI22 U17489 ( .A1(n27484), .A2(n1183), .B1(ram[4327]), .B2(n1184), 
        .ZN(n8568) );
  MOAI22 U17490 ( .A1(n29129), .A2(n1185), .B1(ram[4328]), .B2(n1186), 
        .ZN(n8569) );
  MOAI22 U17491 ( .A1(n28894), .A2(n1185), .B1(ram[4329]), .B2(n1186), 
        .ZN(n8570) );
  MOAI22 U17492 ( .A1(n28659), .A2(n1185), .B1(ram[4330]), .B2(n1186), 
        .ZN(n8571) );
  MOAI22 U17493 ( .A1(n28424), .A2(n1185), .B1(ram[4331]), .B2(n1186), 
        .ZN(n8572) );
  MOAI22 U17494 ( .A1(n28189), .A2(n1185), .B1(ram[4332]), .B2(n1186), 
        .ZN(n8573) );
  MOAI22 U17495 ( .A1(n27954), .A2(n1185), .B1(ram[4333]), .B2(n1186), 
        .ZN(n8574) );
  MOAI22 U17496 ( .A1(n27719), .A2(n1185), .B1(ram[4334]), .B2(n1186), 
        .ZN(n8575) );
  MOAI22 U17497 ( .A1(n27484), .A2(n1185), .B1(ram[4335]), .B2(n1186), 
        .ZN(n8576) );
  MOAI22 U17498 ( .A1(n29129), .A2(n1187), .B1(ram[4336]), .B2(n1188), 
        .ZN(n8577) );
  MOAI22 U17499 ( .A1(n28894), .A2(n1187), .B1(ram[4337]), .B2(n1188), 
        .ZN(n8578) );
  MOAI22 U17500 ( .A1(n28659), .A2(n1187), .B1(ram[4338]), .B2(n1188), 
        .ZN(n8579) );
  MOAI22 U17501 ( .A1(n28424), .A2(n1187), .B1(ram[4339]), .B2(n1188), 
        .ZN(n8580) );
  MOAI22 U17502 ( .A1(n28189), .A2(n1187), .B1(ram[4340]), .B2(n1188), 
        .ZN(n8581) );
  MOAI22 U17503 ( .A1(n27954), .A2(n1187), .B1(ram[4341]), .B2(n1188), 
        .ZN(n8582) );
  MOAI22 U17504 ( .A1(n27719), .A2(n1187), .B1(ram[4342]), .B2(n1188), 
        .ZN(n8583) );
  MOAI22 U17505 ( .A1(n27484), .A2(n1187), .B1(ram[4343]), .B2(n1188), 
        .ZN(n8584) );
  MOAI22 U17506 ( .A1(n29129), .A2(n1189), .B1(ram[4344]), .B2(n1190), 
        .ZN(n8585) );
  MOAI22 U17507 ( .A1(n28894), .A2(n1189), .B1(ram[4345]), .B2(n1190), 
        .ZN(n8586) );
  MOAI22 U17508 ( .A1(n28659), .A2(n1189), .B1(ram[4346]), .B2(n1190), 
        .ZN(n8587) );
  MOAI22 U17509 ( .A1(n28424), .A2(n1189), .B1(ram[4347]), .B2(n1190), 
        .ZN(n8588) );
  MOAI22 U17510 ( .A1(n28189), .A2(n1189), .B1(ram[4348]), .B2(n1190), 
        .ZN(n8589) );
  MOAI22 U17511 ( .A1(n27954), .A2(n1189), .B1(ram[4349]), .B2(n1190), 
        .ZN(n8590) );
  MOAI22 U17512 ( .A1(n27719), .A2(n1189), .B1(ram[4350]), .B2(n1190), 
        .ZN(n8591) );
  MOAI22 U17513 ( .A1(n27484), .A2(n1189), .B1(ram[4351]), .B2(n1190), 
        .ZN(n8592) );
  MOAI22 U17514 ( .A1(n29129), .A2(n1191), .B1(ram[4352]), .B2(n1192), 
        .ZN(n8593) );
  MOAI22 U17515 ( .A1(n28894), .A2(n1191), .B1(ram[4353]), .B2(n1192), 
        .ZN(n8594) );
  MOAI22 U17516 ( .A1(n28659), .A2(n1191), .B1(ram[4354]), .B2(n1192), 
        .ZN(n8595) );
  MOAI22 U17517 ( .A1(n28424), .A2(n1191), .B1(ram[4355]), .B2(n1192), 
        .ZN(n8596) );
  MOAI22 U17518 ( .A1(n28189), .A2(n1191), .B1(ram[4356]), .B2(n1192), 
        .ZN(n8597) );
  MOAI22 U17519 ( .A1(n27954), .A2(n1191), .B1(ram[4357]), .B2(n1192), 
        .ZN(n8598) );
  MOAI22 U17520 ( .A1(n27719), .A2(n1191), .B1(ram[4358]), .B2(n1192), 
        .ZN(n8599) );
  MOAI22 U17521 ( .A1(n27484), .A2(n1191), .B1(ram[4359]), .B2(n1192), 
        .ZN(n8600) );
  MOAI22 U17522 ( .A1(n29129), .A2(n1193), .B1(ram[4360]), .B2(n1194), 
        .ZN(n8601) );
  MOAI22 U17523 ( .A1(n28894), .A2(n1193), .B1(ram[4361]), .B2(n1194), 
        .ZN(n8602) );
  MOAI22 U17524 ( .A1(n28659), .A2(n1193), .B1(ram[4362]), .B2(n1194), 
        .ZN(n8603) );
  MOAI22 U17525 ( .A1(n28424), .A2(n1193), .B1(ram[4363]), .B2(n1194), 
        .ZN(n8604) );
  MOAI22 U17526 ( .A1(n28189), .A2(n1193), .B1(ram[4364]), .B2(n1194), 
        .ZN(n8605) );
  MOAI22 U17527 ( .A1(n27954), .A2(n1193), .B1(ram[4365]), .B2(n1194), 
        .ZN(n8606) );
  MOAI22 U17528 ( .A1(n27719), .A2(n1193), .B1(ram[4366]), .B2(n1194), 
        .ZN(n8607) );
  MOAI22 U17529 ( .A1(n27484), .A2(n1193), .B1(ram[4367]), .B2(n1194), 
        .ZN(n8608) );
  MOAI22 U17530 ( .A1(n29130), .A2(n1195), .B1(ram[4368]), .B2(n1196), 
        .ZN(n8609) );
  MOAI22 U17531 ( .A1(n28895), .A2(n1195), .B1(ram[4369]), .B2(n1196), 
        .ZN(n8610) );
  MOAI22 U17532 ( .A1(n28660), .A2(n1195), .B1(ram[4370]), .B2(n1196), 
        .ZN(n8611) );
  MOAI22 U17533 ( .A1(n28425), .A2(n1195), .B1(ram[4371]), .B2(n1196), 
        .ZN(n8612) );
  MOAI22 U17534 ( .A1(n28190), .A2(n1195), .B1(ram[4372]), .B2(n1196), 
        .ZN(n8613) );
  MOAI22 U17535 ( .A1(n27955), .A2(n1195), .B1(ram[4373]), .B2(n1196), 
        .ZN(n8614) );
  MOAI22 U17536 ( .A1(n27720), .A2(n1195), .B1(ram[4374]), .B2(n1196), 
        .ZN(n8615) );
  MOAI22 U17537 ( .A1(n27485), .A2(n1195), .B1(ram[4375]), .B2(n1196), 
        .ZN(n8616) );
  MOAI22 U17538 ( .A1(n29130), .A2(n1197), .B1(ram[4376]), .B2(n1198), 
        .ZN(n8617) );
  MOAI22 U17539 ( .A1(n28895), .A2(n1197), .B1(ram[4377]), .B2(n1198), 
        .ZN(n8618) );
  MOAI22 U17540 ( .A1(n28660), .A2(n1197), .B1(ram[4378]), .B2(n1198), 
        .ZN(n8619) );
  MOAI22 U17541 ( .A1(n28425), .A2(n1197), .B1(ram[4379]), .B2(n1198), 
        .ZN(n8620) );
  MOAI22 U17542 ( .A1(n28190), .A2(n1197), .B1(ram[4380]), .B2(n1198), 
        .ZN(n8621) );
  MOAI22 U17543 ( .A1(n27955), .A2(n1197), .B1(ram[4381]), .B2(n1198), 
        .ZN(n8622) );
  MOAI22 U17544 ( .A1(n27720), .A2(n1197), .B1(ram[4382]), .B2(n1198), 
        .ZN(n8623) );
  MOAI22 U17545 ( .A1(n27485), .A2(n1197), .B1(ram[4383]), .B2(n1198), 
        .ZN(n8624) );
  MOAI22 U17546 ( .A1(n29130), .A2(n1199), .B1(ram[4384]), .B2(n1200), 
        .ZN(n8625) );
  MOAI22 U17547 ( .A1(n28895), .A2(n1199), .B1(ram[4385]), .B2(n1200), 
        .ZN(n8626) );
  MOAI22 U17548 ( .A1(n28660), .A2(n1199), .B1(ram[4386]), .B2(n1200), 
        .ZN(n8627) );
  MOAI22 U17549 ( .A1(n28425), .A2(n1199), .B1(ram[4387]), .B2(n1200), 
        .ZN(n8628) );
  MOAI22 U17550 ( .A1(n28190), .A2(n1199), .B1(ram[4388]), .B2(n1200), 
        .ZN(n8629) );
  MOAI22 U17551 ( .A1(n27955), .A2(n1199), .B1(ram[4389]), .B2(n1200), 
        .ZN(n8630) );
  MOAI22 U17552 ( .A1(n27720), .A2(n1199), .B1(ram[4390]), .B2(n1200), 
        .ZN(n8631) );
  MOAI22 U17553 ( .A1(n27485), .A2(n1199), .B1(ram[4391]), .B2(n1200), 
        .ZN(n8632) );
  MOAI22 U17554 ( .A1(n29130), .A2(n1201), .B1(ram[4392]), .B2(n1202), 
        .ZN(n8633) );
  MOAI22 U17555 ( .A1(n28895), .A2(n1201), .B1(ram[4393]), .B2(n1202), 
        .ZN(n8634) );
  MOAI22 U17556 ( .A1(n28660), .A2(n1201), .B1(ram[4394]), .B2(n1202), 
        .ZN(n8635) );
  MOAI22 U17557 ( .A1(n28425), .A2(n1201), .B1(ram[4395]), .B2(n1202), 
        .ZN(n8636) );
  MOAI22 U17558 ( .A1(n28190), .A2(n1201), .B1(ram[4396]), .B2(n1202), 
        .ZN(n8637) );
  MOAI22 U17559 ( .A1(n27955), .A2(n1201), .B1(ram[4397]), .B2(n1202), 
        .ZN(n8638) );
  MOAI22 U17560 ( .A1(n27720), .A2(n1201), .B1(ram[4398]), .B2(n1202), 
        .ZN(n8639) );
  MOAI22 U17561 ( .A1(n27485), .A2(n1201), .B1(ram[4399]), .B2(n1202), 
        .ZN(n8640) );
  MOAI22 U17562 ( .A1(n29130), .A2(n1203), .B1(ram[4400]), .B2(n1204), 
        .ZN(n8641) );
  MOAI22 U17563 ( .A1(n28895), .A2(n1203), .B1(ram[4401]), .B2(n1204), 
        .ZN(n8642) );
  MOAI22 U17564 ( .A1(n28660), .A2(n1203), .B1(ram[4402]), .B2(n1204), 
        .ZN(n8643) );
  MOAI22 U17565 ( .A1(n28425), .A2(n1203), .B1(ram[4403]), .B2(n1204), 
        .ZN(n8644) );
  MOAI22 U17566 ( .A1(n28190), .A2(n1203), .B1(ram[4404]), .B2(n1204), 
        .ZN(n8645) );
  MOAI22 U17567 ( .A1(n27955), .A2(n1203), .B1(ram[4405]), .B2(n1204), 
        .ZN(n8646) );
  MOAI22 U17568 ( .A1(n27720), .A2(n1203), .B1(ram[4406]), .B2(n1204), 
        .ZN(n8647) );
  MOAI22 U17569 ( .A1(n27485), .A2(n1203), .B1(ram[4407]), .B2(n1204), 
        .ZN(n8648) );
  MOAI22 U17570 ( .A1(n29130), .A2(n1205), .B1(ram[4408]), .B2(n1206), 
        .ZN(n8649) );
  MOAI22 U17571 ( .A1(n28895), .A2(n1205), .B1(ram[4409]), .B2(n1206), 
        .ZN(n8650) );
  MOAI22 U17572 ( .A1(n28660), .A2(n1205), .B1(ram[4410]), .B2(n1206), 
        .ZN(n8651) );
  MOAI22 U17573 ( .A1(n28425), .A2(n1205), .B1(ram[4411]), .B2(n1206), 
        .ZN(n8652) );
  MOAI22 U17574 ( .A1(n28190), .A2(n1205), .B1(ram[4412]), .B2(n1206), 
        .ZN(n8653) );
  MOAI22 U17575 ( .A1(n27955), .A2(n1205), .B1(ram[4413]), .B2(n1206), 
        .ZN(n8654) );
  MOAI22 U17576 ( .A1(n27720), .A2(n1205), .B1(ram[4414]), .B2(n1206), 
        .ZN(n8655) );
  MOAI22 U17577 ( .A1(n27485), .A2(n1205), .B1(ram[4415]), .B2(n1206), 
        .ZN(n8656) );
  MOAI22 U17578 ( .A1(n29130), .A2(n1207), .B1(ram[4416]), .B2(n1208), 
        .ZN(n8657) );
  MOAI22 U17579 ( .A1(n28895), .A2(n1207), .B1(ram[4417]), .B2(n1208), 
        .ZN(n8658) );
  MOAI22 U17580 ( .A1(n28660), .A2(n1207), .B1(ram[4418]), .B2(n1208), 
        .ZN(n8659) );
  MOAI22 U17581 ( .A1(n28425), .A2(n1207), .B1(ram[4419]), .B2(n1208), 
        .ZN(n8660) );
  MOAI22 U17582 ( .A1(n28190), .A2(n1207), .B1(ram[4420]), .B2(n1208), 
        .ZN(n8661) );
  MOAI22 U17583 ( .A1(n27955), .A2(n1207), .B1(ram[4421]), .B2(n1208), 
        .ZN(n8662) );
  MOAI22 U17584 ( .A1(n27720), .A2(n1207), .B1(ram[4422]), .B2(n1208), 
        .ZN(n8663) );
  MOAI22 U17585 ( .A1(n27485), .A2(n1207), .B1(ram[4423]), .B2(n1208), 
        .ZN(n8664) );
  MOAI22 U17586 ( .A1(n29130), .A2(n1209), .B1(ram[4424]), .B2(n1210), 
        .ZN(n8665) );
  MOAI22 U17587 ( .A1(n28895), .A2(n1209), .B1(ram[4425]), .B2(n1210), 
        .ZN(n8666) );
  MOAI22 U17588 ( .A1(n28660), .A2(n1209), .B1(ram[4426]), .B2(n1210), 
        .ZN(n8667) );
  MOAI22 U17589 ( .A1(n28425), .A2(n1209), .B1(ram[4427]), .B2(n1210), 
        .ZN(n8668) );
  MOAI22 U17590 ( .A1(n28190), .A2(n1209), .B1(ram[4428]), .B2(n1210), 
        .ZN(n8669) );
  MOAI22 U17591 ( .A1(n27955), .A2(n1209), .B1(ram[4429]), .B2(n1210), 
        .ZN(n8670) );
  MOAI22 U17592 ( .A1(n27720), .A2(n1209), .B1(ram[4430]), .B2(n1210), 
        .ZN(n8671) );
  MOAI22 U17593 ( .A1(n27485), .A2(n1209), .B1(ram[4431]), .B2(n1210), 
        .ZN(n8672) );
  MOAI22 U17594 ( .A1(n29130), .A2(n1211), .B1(ram[4432]), .B2(n1212), 
        .ZN(n8673) );
  MOAI22 U17595 ( .A1(n28895), .A2(n1211), .B1(ram[4433]), .B2(n1212), 
        .ZN(n8674) );
  MOAI22 U17596 ( .A1(n28660), .A2(n1211), .B1(ram[4434]), .B2(n1212), 
        .ZN(n8675) );
  MOAI22 U17597 ( .A1(n28425), .A2(n1211), .B1(ram[4435]), .B2(n1212), 
        .ZN(n8676) );
  MOAI22 U17598 ( .A1(n28190), .A2(n1211), .B1(ram[4436]), .B2(n1212), 
        .ZN(n8677) );
  MOAI22 U17599 ( .A1(n27955), .A2(n1211), .B1(ram[4437]), .B2(n1212), 
        .ZN(n8678) );
  MOAI22 U17600 ( .A1(n27720), .A2(n1211), .B1(ram[4438]), .B2(n1212), 
        .ZN(n8679) );
  MOAI22 U17601 ( .A1(n27485), .A2(n1211), .B1(ram[4439]), .B2(n1212), 
        .ZN(n8680) );
  MOAI22 U17602 ( .A1(n29130), .A2(n1213), .B1(ram[4440]), .B2(n1214), 
        .ZN(n8681) );
  MOAI22 U17603 ( .A1(n28895), .A2(n1213), .B1(ram[4441]), .B2(n1214), 
        .ZN(n8682) );
  MOAI22 U17604 ( .A1(n28660), .A2(n1213), .B1(ram[4442]), .B2(n1214), 
        .ZN(n8683) );
  MOAI22 U17605 ( .A1(n28425), .A2(n1213), .B1(ram[4443]), .B2(n1214), 
        .ZN(n8684) );
  MOAI22 U17606 ( .A1(n28190), .A2(n1213), .B1(ram[4444]), .B2(n1214), 
        .ZN(n8685) );
  MOAI22 U17607 ( .A1(n27955), .A2(n1213), .B1(ram[4445]), .B2(n1214), 
        .ZN(n8686) );
  MOAI22 U17608 ( .A1(n27720), .A2(n1213), .B1(ram[4446]), .B2(n1214), 
        .ZN(n8687) );
  MOAI22 U17609 ( .A1(n27485), .A2(n1213), .B1(ram[4447]), .B2(n1214), 
        .ZN(n8688) );
  MOAI22 U17610 ( .A1(n29130), .A2(n1215), .B1(ram[4448]), .B2(n1216), 
        .ZN(n8689) );
  MOAI22 U17611 ( .A1(n28895), .A2(n1215), .B1(ram[4449]), .B2(n1216), 
        .ZN(n8690) );
  MOAI22 U17612 ( .A1(n28660), .A2(n1215), .B1(ram[4450]), .B2(n1216), 
        .ZN(n8691) );
  MOAI22 U17613 ( .A1(n28425), .A2(n1215), .B1(ram[4451]), .B2(n1216), 
        .ZN(n8692) );
  MOAI22 U17614 ( .A1(n28190), .A2(n1215), .B1(ram[4452]), .B2(n1216), 
        .ZN(n8693) );
  MOAI22 U17615 ( .A1(n27955), .A2(n1215), .B1(ram[4453]), .B2(n1216), 
        .ZN(n8694) );
  MOAI22 U17616 ( .A1(n27720), .A2(n1215), .B1(ram[4454]), .B2(n1216), 
        .ZN(n8695) );
  MOAI22 U17617 ( .A1(n27485), .A2(n1215), .B1(ram[4455]), .B2(n1216), 
        .ZN(n8696) );
  MOAI22 U17618 ( .A1(n29130), .A2(n1217), .B1(ram[4456]), .B2(n1218), 
        .ZN(n8697) );
  MOAI22 U17619 ( .A1(n28895), .A2(n1217), .B1(ram[4457]), .B2(n1218), 
        .ZN(n8698) );
  MOAI22 U17620 ( .A1(n28660), .A2(n1217), .B1(ram[4458]), .B2(n1218), 
        .ZN(n8699) );
  MOAI22 U17621 ( .A1(n28425), .A2(n1217), .B1(ram[4459]), .B2(n1218), 
        .ZN(n8700) );
  MOAI22 U17622 ( .A1(n28190), .A2(n1217), .B1(ram[4460]), .B2(n1218), 
        .ZN(n8701) );
  MOAI22 U17623 ( .A1(n27955), .A2(n1217), .B1(ram[4461]), .B2(n1218), 
        .ZN(n8702) );
  MOAI22 U17624 ( .A1(n27720), .A2(n1217), .B1(ram[4462]), .B2(n1218), 
        .ZN(n8703) );
  MOAI22 U17625 ( .A1(n27485), .A2(n1217), .B1(ram[4463]), .B2(n1218), 
        .ZN(n8704) );
  MOAI22 U17626 ( .A1(n29130), .A2(n1219), .B1(ram[4464]), .B2(n1220), 
        .ZN(n8705) );
  MOAI22 U17627 ( .A1(n28895), .A2(n1219), .B1(ram[4465]), .B2(n1220), 
        .ZN(n8706) );
  MOAI22 U17628 ( .A1(n28660), .A2(n1219), .B1(ram[4466]), .B2(n1220), 
        .ZN(n8707) );
  MOAI22 U17629 ( .A1(n28425), .A2(n1219), .B1(ram[4467]), .B2(n1220), 
        .ZN(n8708) );
  MOAI22 U17630 ( .A1(n28190), .A2(n1219), .B1(ram[4468]), .B2(n1220), 
        .ZN(n8709) );
  MOAI22 U17631 ( .A1(n27955), .A2(n1219), .B1(ram[4469]), .B2(n1220), 
        .ZN(n8710) );
  MOAI22 U17632 ( .A1(n27720), .A2(n1219), .B1(ram[4470]), .B2(n1220), 
        .ZN(n8711) );
  MOAI22 U17633 ( .A1(n27485), .A2(n1219), .B1(ram[4471]), .B2(n1220), 
        .ZN(n8712) );
  MOAI22 U17634 ( .A1(n29131), .A2(n1221), .B1(ram[4472]), .B2(n1222), 
        .ZN(n8713) );
  MOAI22 U17635 ( .A1(n28896), .A2(n1221), .B1(ram[4473]), .B2(n1222), 
        .ZN(n8714) );
  MOAI22 U17636 ( .A1(n28661), .A2(n1221), .B1(ram[4474]), .B2(n1222), 
        .ZN(n8715) );
  MOAI22 U17637 ( .A1(n28426), .A2(n1221), .B1(ram[4475]), .B2(n1222), 
        .ZN(n8716) );
  MOAI22 U17638 ( .A1(n28191), .A2(n1221), .B1(ram[4476]), .B2(n1222), 
        .ZN(n8717) );
  MOAI22 U17639 ( .A1(n27956), .A2(n1221), .B1(ram[4477]), .B2(n1222), 
        .ZN(n8718) );
  MOAI22 U17640 ( .A1(n27721), .A2(n1221), .B1(ram[4478]), .B2(n1222), 
        .ZN(n8719) );
  MOAI22 U17641 ( .A1(n27486), .A2(n1221), .B1(ram[4479]), .B2(n1222), 
        .ZN(n8720) );
  MOAI22 U17642 ( .A1(n29131), .A2(n1223), .B1(ram[4480]), .B2(n1224), 
        .ZN(n8721) );
  MOAI22 U17643 ( .A1(n28896), .A2(n1223), .B1(ram[4481]), .B2(n1224), 
        .ZN(n8722) );
  MOAI22 U17644 ( .A1(n28661), .A2(n1223), .B1(ram[4482]), .B2(n1224), 
        .ZN(n8723) );
  MOAI22 U17645 ( .A1(n28426), .A2(n1223), .B1(ram[4483]), .B2(n1224), 
        .ZN(n8724) );
  MOAI22 U17646 ( .A1(n28191), .A2(n1223), .B1(ram[4484]), .B2(n1224), 
        .ZN(n8725) );
  MOAI22 U17647 ( .A1(n27956), .A2(n1223), .B1(ram[4485]), .B2(n1224), 
        .ZN(n8726) );
  MOAI22 U17648 ( .A1(n27721), .A2(n1223), .B1(ram[4486]), .B2(n1224), 
        .ZN(n8727) );
  MOAI22 U17649 ( .A1(n27486), .A2(n1223), .B1(ram[4487]), .B2(n1224), 
        .ZN(n8728) );
  MOAI22 U17650 ( .A1(n29131), .A2(n1225), .B1(ram[4488]), .B2(n1226), 
        .ZN(n8729) );
  MOAI22 U17651 ( .A1(n28896), .A2(n1225), .B1(ram[4489]), .B2(n1226), 
        .ZN(n8730) );
  MOAI22 U17652 ( .A1(n28661), .A2(n1225), .B1(ram[4490]), .B2(n1226), 
        .ZN(n8731) );
  MOAI22 U17653 ( .A1(n28426), .A2(n1225), .B1(ram[4491]), .B2(n1226), 
        .ZN(n8732) );
  MOAI22 U17654 ( .A1(n28191), .A2(n1225), .B1(ram[4492]), .B2(n1226), 
        .ZN(n8733) );
  MOAI22 U17655 ( .A1(n27956), .A2(n1225), .B1(ram[4493]), .B2(n1226), 
        .ZN(n8734) );
  MOAI22 U17656 ( .A1(n27721), .A2(n1225), .B1(ram[4494]), .B2(n1226), 
        .ZN(n8735) );
  MOAI22 U17657 ( .A1(n27486), .A2(n1225), .B1(ram[4495]), .B2(n1226), 
        .ZN(n8736) );
  MOAI22 U17658 ( .A1(n29131), .A2(n1227), .B1(ram[4496]), .B2(n1228), 
        .ZN(n8737) );
  MOAI22 U17659 ( .A1(n28896), .A2(n1227), .B1(ram[4497]), .B2(n1228), 
        .ZN(n8738) );
  MOAI22 U17660 ( .A1(n28661), .A2(n1227), .B1(ram[4498]), .B2(n1228), 
        .ZN(n8739) );
  MOAI22 U17661 ( .A1(n28426), .A2(n1227), .B1(ram[4499]), .B2(n1228), 
        .ZN(n8740) );
  MOAI22 U17662 ( .A1(n28191), .A2(n1227), .B1(ram[4500]), .B2(n1228), 
        .ZN(n8741) );
  MOAI22 U17663 ( .A1(n27956), .A2(n1227), .B1(ram[4501]), .B2(n1228), 
        .ZN(n8742) );
  MOAI22 U17664 ( .A1(n27721), .A2(n1227), .B1(ram[4502]), .B2(n1228), 
        .ZN(n8743) );
  MOAI22 U17665 ( .A1(n27486), .A2(n1227), .B1(ram[4503]), .B2(n1228), 
        .ZN(n8744) );
  MOAI22 U17666 ( .A1(n29131), .A2(n1229), .B1(ram[4504]), .B2(n1230), 
        .ZN(n8745) );
  MOAI22 U17667 ( .A1(n28896), .A2(n1229), .B1(ram[4505]), .B2(n1230), 
        .ZN(n8746) );
  MOAI22 U17668 ( .A1(n28661), .A2(n1229), .B1(ram[4506]), .B2(n1230), 
        .ZN(n8747) );
  MOAI22 U17669 ( .A1(n28426), .A2(n1229), .B1(ram[4507]), .B2(n1230), 
        .ZN(n8748) );
  MOAI22 U17670 ( .A1(n28191), .A2(n1229), .B1(ram[4508]), .B2(n1230), 
        .ZN(n8749) );
  MOAI22 U17671 ( .A1(n27956), .A2(n1229), .B1(ram[4509]), .B2(n1230), 
        .ZN(n8750) );
  MOAI22 U17672 ( .A1(n27721), .A2(n1229), .B1(ram[4510]), .B2(n1230), 
        .ZN(n8751) );
  MOAI22 U17673 ( .A1(n27486), .A2(n1229), .B1(ram[4511]), .B2(n1230), 
        .ZN(n8752) );
  MOAI22 U17674 ( .A1(n29131), .A2(n1231), .B1(ram[4512]), .B2(n1232), 
        .ZN(n8753) );
  MOAI22 U17675 ( .A1(n28896), .A2(n1231), .B1(ram[4513]), .B2(n1232), 
        .ZN(n8754) );
  MOAI22 U17676 ( .A1(n28661), .A2(n1231), .B1(ram[4514]), .B2(n1232), 
        .ZN(n8755) );
  MOAI22 U17677 ( .A1(n28426), .A2(n1231), .B1(ram[4515]), .B2(n1232), 
        .ZN(n8756) );
  MOAI22 U17678 ( .A1(n28191), .A2(n1231), .B1(ram[4516]), .B2(n1232), 
        .ZN(n8757) );
  MOAI22 U17679 ( .A1(n27956), .A2(n1231), .B1(ram[4517]), .B2(n1232), 
        .ZN(n8758) );
  MOAI22 U17680 ( .A1(n27721), .A2(n1231), .B1(ram[4518]), .B2(n1232), 
        .ZN(n8759) );
  MOAI22 U17681 ( .A1(n27486), .A2(n1231), .B1(ram[4519]), .B2(n1232), 
        .ZN(n8760) );
  MOAI22 U17682 ( .A1(n29131), .A2(n1233), .B1(ram[4520]), .B2(n1234), 
        .ZN(n8761) );
  MOAI22 U17683 ( .A1(n28896), .A2(n1233), .B1(ram[4521]), .B2(n1234), 
        .ZN(n8762) );
  MOAI22 U17684 ( .A1(n28661), .A2(n1233), .B1(ram[4522]), .B2(n1234), 
        .ZN(n8763) );
  MOAI22 U17685 ( .A1(n28426), .A2(n1233), .B1(ram[4523]), .B2(n1234), 
        .ZN(n8764) );
  MOAI22 U17686 ( .A1(n28191), .A2(n1233), .B1(ram[4524]), .B2(n1234), 
        .ZN(n8765) );
  MOAI22 U17687 ( .A1(n27956), .A2(n1233), .B1(ram[4525]), .B2(n1234), 
        .ZN(n8766) );
  MOAI22 U17688 ( .A1(n27721), .A2(n1233), .B1(ram[4526]), .B2(n1234), 
        .ZN(n8767) );
  MOAI22 U17689 ( .A1(n27486), .A2(n1233), .B1(ram[4527]), .B2(n1234), 
        .ZN(n8768) );
  MOAI22 U17690 ( .A1(n29131), .A2(n1235), .B1(ram[4528]), .B2(n1236), 
        .ZN(n8769) );
  MOAI22 U17691 ( .A1(n28896), .A2(n1235), .B1(ram[4529]), .B2(n1236), 
        .ZN(n8770) );
  MOAI22 U17692 ( .A1(n28661), .A2(n1235), .B1(ram[4530]), .B2(n1236), 
        .ZN(n8771) );
  MOAI22 U17693 ( .A1(n28426), .A2(n1235), .B1(ram[4531]), .B2(n1236), 
        .ZN(n8772) );
  MOAI22 U17694 ( .A1(n28191), .A2(n1235), .B1(ram[4532]), .B2(n1236), 
        .ZN(n8773) );
  MOAI22 U17695 ( .A1(n27956), .A2(n1235), .B1(ram[4533]), .B2(n1236), 
        .ZN(n8774) );
  MOAI22 U17696 ( .A1(n27721), .A2(n1235), .B1(ram[4534]), .B2(n1236), 
        .ZN(n8775) );
  MOAI22 U17697 ( .A1(n27486), .A2(n1235), .B1(ram[4535]), .B2(n1236), 
        .ZN(n8776) );
  MOAI22 U17698 ( .A1(n29131), .A2(n1237), .B1(ram[4536]), .B2(n1238), 
        .ZN(n8777) );
  MOAI22 U17699 ( .A1(n28896), .A2(n1237), .B1(ram[4537]), .B2(n1238), 
        .ZN(n8778) );
  MOAI22 U17700 ( .A1(n28661), .A2(n1237), .B1(ram[4538]), .B2(n1238), 
        .ZN(n8779) );
  MOAI22 U17701 ( .A1(n28426), .A2(n1237), .B1(ram[4539]), .B2(n1238), 
        .ZN(n8780) );
  MOAI22 U17702 ( .A1(n28191), .A2(n1237), .B1(ram[4540]), .B2(n1238), 
        .ZN(n8781) );
  MOAI22 U17703 ( .A1(n27956), .A2(n1237), .B1(ram[4541]), .B2(n1238), 
        .ZN(n8782) );
  MOAI22 U17704 ( .A1(n27721), .A2(n1237), .B1(ram[4542]), .B2(n1238), 
        .ZN(n8783) );
  MOAI22 U17705 ( .A1(n27486), .A2(n1237), .B1(ram[4543]), .B2(n1238), 
        .ZN(n8784) );
  MOAI22 U17706 ( .A1(n29131), .A2(n1239), .B1(ram[4544]), .B2(n1240), 
        .ZN(n8785) );
  MOAI22 U17707 ( .A1(n28896), .A2(n1239), .B1(ram[4545]), .B2(n1240), 
        .ZN(n8786) );
  MOAI22 U17708 ( .A1(n28661), .A2(n1239), .B1(ram[4546]), .B2(n1240), 
        .ZN(n8787) );
  MOAI22 U17709 ( .A1(n28426), .A2(n1239), .B1(ram[4547]), .B2(n1240), 
        .ZN(n8788) );
  MOAI22 U17710 ( .A1(n28191), .A2(n1239), .B1(ram[4548]), .B2(n1240), 
        .ZN(n8789) );
  MOAI22 U17711 ( .A1(n27956), .A2(n1239), .B1(ram[4549]), .B2(n1240), 
        .ZN(n8790) );
  MOAI22 U17712 ( .A1(n27721), .A2(n1239), .B1(ram[4550]), .B2(n1240), 
        .ZN(n8791) );
  MOAI22 U17713 ( .A1(n27486), .A2(n1239), .B1(ram[4551]), .B2(n1240), 
        .ZN(n8792) );
  MOAI22 U17714 ( .A1(n29131), .A2(n1241), .B1(ram[4552]), .B2(n1242), 
        .ZN(n8793) );
  MOAI22 U17715 ( .A1(n28896), .A2(n1241), .B1(ram[4553]), .B2(n1242), 
        .ZN(n8794) );
  MOAI22 U17716 ( .A1(n28661), .A2(n1241), .B1(ram[4554]), .B2(n1242), 
        .ZN(n8795) );
  MOAI22 U17717 ( .A1(n28426), .A2(n1241), .B1(ram[4555]), .B2(n1242), 
        .ZN(n8796) );
  MOAI22 U17718 ( .A1(n28191), .A2(n1241), .B1(ram[4556]), .B2(n1242), 
        .ZN(n8797) );
  MOAI22 U17719 ( .A1(n27956), .A2(n1241), .B1(ram[4557]), .B2(n1242), 
        .ZN(n8798) );
  MOAI22 U17720 ( .A1(n27721), .A2(n1241), .B1(ram[4558]), .B2(n1242), 
        .ZN(n8799) );
  MOAI22 U17721 ( .A1(n27486), .A2(n1241), .B1(ram[4559]), .B2(n1242), 
        .ZN(n8800) );
  MOAI22 U17722 ( .A1(n29131), .A2(n1243), .B1(ram[4560]), .B2(n1244), 
        .ZN(n8801) );
  MOAI22 U17723 ( .A1(n28896), .A2(n1243), .B1(ram[4561]), .B2(n1244), 
        .ZN(n8802) );
  MOAI22 U17724 ( .A1(n28661), .A2(n1243), .B1(ram[4562]), .B2(n1244), 
        .ZN(n8803) );
  MOAI22 U17725 ( .A1(n28426), .A2(n1243), .B1(ram[4563]), .B2(n1244), 
        .ZN(n8804) );
  MOAI22 U17726 ( .A1(n28191), .A2(n1243), .B1(ram[4564]), .B2(n1244), 
        .ZN(n8805) );
  MOAI22 U17727 ( .A1(n27956), .A2(n1243), .B1(ram[4565]), .B2(n1244), 
        .ZN(n8806) );
  MOAI22 U17728 ( .A1(n27721), .A2(n1243), .B1(ram[4566]), .B2(n1244), 
        .ZN(n8807) );
  MOAI22 U17729 ( .A1(n27486), .A2(n1243), .B1(ram[4567]), .B2(n1244), 
        .ZN(n8808) );
  MOAI22 U17730 ( .A1(n29131), .A2(n1245), .B1(ram[4568]), .B2(n1246), 
        .ZN(n8809) );
  MOAI22 U17731 ( .A1(n28896), .A2(n1245), .B1(ram[4569]), .B2(n1246), 
        .ZN(n8810) );
  MOAI22 U17732 ( .A1(n28661), .A2(n1245), .B1(ram[4570]), .B2(n1246), 
        .ZN(n8811) );
  MOAI22 U17733 ( .A1(n28426), .A2(n1245), .B1(ram[4571]), .B2(n1246), 
        .ZN(n8812) );
  MOAI22 U17734 ( .A1(n28191), .A2(n1245), .B1(ram[4572]), .B2(n1246), 
        .ZN(n8813) );
  MOAI22 U17735 ( .A1(n27956), .A2(n1245), .B1(ram[4573]), .B2(n1246), 
        .ZN(n8814) );
  MOAI22 U17736 ( .A1(n27721), .A2(n1245), .B1(ram[4574]), .B2(n1246), 
        .ZN(n8815) );
  MOAI22 U17737 ( .A1(n27486), .A2(n1245), .B1(ram[4575]), .B2(n1246), 
        .ZN(n8816) );
  MOAI22 U17738 ( .A1(n29132), .A2(n1247), .B1(ram[4576]), .B2(n1248), 
        .ZN(n8817) );
  MOAI22 U17739 ( .A1(n28897), .A2(n1247), .B1(ram[4577]), .B2(n1248), 
        .ZN(n8818) );
  MOAI22 U17740 ( .A1(n28662), .A2(n1247), .B1(ram[4578]), .B2(n1248), 
        .ZN(n8819) );
  MOAI22 U17741 ( .A1(n28427), .A2(n1247), .B1(ram[4579]), .B2(n1248), 
        .ZN(n8820) );
  MOAI22 U17742 ( .A1(n28192), .A2(n1247), .B1(ram[4580]), .B2(n1248), 
        .ZN(n8821) );
  MOAI22 U17743 ( .A1(n27957), .A2(n1247), .B1(ram[4581]), .B2(n1248), 
        .ZN(n8822) );
  MOAI22 U17744 ( .A1(n27722), .A2(n1247), .B1(ram[4582]), .B2(n1248), 
        .ZN(n8823) );
  MOAI22 U17745 ( .A1(n27487), .A2(n1247), .B1(ram[4583]), .B2(n1248), 
        .ZN(n8824) );
  MOAI22 U17746 ( .A1(n29132), .A2(n1249), .B1(ram[4584]), .B2(n1250), 
        .ZN(n8825) );
  MOAI22 U17747 ( .A1(n28897), .A2(n1249), .B1(ram[4585]), .B2(n1250), 
        .ZN(n8826) );
  MOAI22 U17748 ( .A1(n28662), .A2(n1249), .B1(ram[4586]), .B2(n1250), 
        .ZN(n8827) );
  MOAI22 U17749 ( .A1(n28427), .A2(n1249), .B1(ram[4587]), .B2(n1250), 
        .ZN(n8828) );
  MOAI22 U17750 ( .A1(n28192), .A2(n1249), .B1(ram[4588]), .B2(n1250), 
        .ZN(n8829) );
  MOAI22 U17751 ( .A1(n27957), .A2(n1249), .B1(ram[4589]), .B2(n1250), 
        .ZN(n8830) );
  MOAI22 U17752 ( .A1(n27722), .A2(n1249), .B1(ram[4590]), .B2(n1250), 
        .ZN(n8831) );
  MOAI22 U17753 ( .A1(n27487), .A2(n1249), .B1(ram[4591]), .B2(n1250), 
        .ZN(n8832) );
  MOAI22 U17754 ( .A1(n29132), .A2(n1251), .B1(ram[4592]), .B2(n1252), 
        .ZN(n8833) );
  MOAI22 U17755 ( .A1(n28897), .A2(n1251), .B1(ram[4593]), .B2(n1252), 
        .ZN(n8834) );
  MOAI22 U17756 ( .A1(n28662), .A2(n1251), .B1(ram[4594]), .B2(n1252), 
        .ZN(n8835) );
  MOAI22 U17757 ( .A1(n28427), .A2(n1251), .B1(ram[4595]), .B2(n1252), 
        .ZN(n8836) );
  MOAI22 U17758 ( .A1(n28192), .A2(n1251), .B1(ram[4596]), .B2(n1252), 
        .ZN(n8837) );
  MOAI22 U17759 ( .A1(n27957), .A2(n1251), .B1(ram[4597]), .B2(n1252), 
        .ZN(n8838) );
  MOAI22 U17760 ( .A1(n27722), .A2(n1251), .B1(ram[4598]), .B2(n1252), 
        .ZN(n8839) );
  MOAI22 U17761 ( .A1(n27487), .A2(n1251), .B1(ram[4599]), .B2(n1252), 
        .ZN(n8840) );
  MOAI22 U17762 ( .A1(n29132), .A2(n1253), .B1(ram[4600]), .B2(n1254), 
        .ZN(n8841) );
  MOAI22 U17763 ( .A1(n28897), .A2(n1253), .B1(ram[4601]), .B2(n1254), 
        .ZN(n8842) );
  MOAI22 U17764 ( .A1(n28662), .A2(n1253), .B1(ram[4602]), .B2(n1254), 
        .ZN(n8843) );
  MOAI22 U17765 ( .A1(n28427), .A2(n1253), .B1(ram[4603]), .B2(n1254), 
        .ZN(n8844) );
  MOAI22 U17766 ( .A1(n28192), .A2(n1253), .B1(ram[4604]), .B2(n1254), 
        .ZN(n8845) );
  MOAI22 U17767 ( .A1(n27957), .A2(n1253), .B1(ram[4605]), .B2(n1254), 
        .ZN(n8846) );
  MOAI22 U17768 ( .A1(n27722), .A2(n1253), .B1(ram[4606]), .B2(n1254), 
        .ZN(n8847) );
  MOAI22 U17769 ( .A1(n27487), .A2(n1253), .B1(ram[4607]), .B2(n1254), 
        .ZN(n8848) );
  MOAI22 U17770 ( .A1(n29132), .A2(n1256), .B1(ram[4608]), .B2(n1257), 
        .ZN(n8849) );
  MOAI22 U17771 ( .A1(n28897), .A2(n1256), .B1(ram[4609]), .B2(n1257), 
        .ZN(n8850) );
  MOAI22 U17772 ( .A1(n28662), .A2(n1256), .B1(ram[4610]), .B2(n1257), 
        .ZN(n8851) );
  MOAI22 U17773 ( .A1(n28427), .A2(n1256), .B1(ram[4611]), .B2(n1257), 
        .ZN(n8852) );
  MOAI22 U17774 ( .A1(n28192), .A2(n1256), .B1(ram[4612]), .B2(n1257), 
        .ZN(n8853) );
  MOAI22 U17775 ( .A1(n27957), .A2(n1256), .B1(ram[4613]), .B2(n1257), 
        .ZN(n8854) );
  MOAI22 U17776 ( .A1(n27722), .A2(n1256), .B1(ram[4614]), .B2(n1257), 
        .ZN(n8855) );
  MOAI22 U17777 ( .A1(n27487), .A2(n1256), .B1(ram[4615]), .B2(n1257), 
        .ZN(n8856) );
  MOAI22 U17778 ( .A1(n29132), .A2(n1259), .B1(ram[4616]), .B2(n1260), 
        .ZN(n8857) );
  MOAI22 U17779 ( .A1(n28897), .A2(n1259), .B1(ram[4617]), .B2(n1260), 
        .ZN(n8858) );
  MOAI22 U17780 ( .A1(n28662), .A2(n1259), .B1(ram[4618]), .B2(n1260), 
        .ZN(n8859) );
  MOAI22 U17781 ( .A1(n28427), .A2(n1259), .B1(ram[4619]), .B2(n1260), 
        .ZN(n8860) );
  MOAI22 U17782 ( .A1(n28192), .A2(n1259), .B1(ram[4620]), .B2(n1260), 
        .ZN(n8861) );
  MOAI22 U17783 ( .A1(n27957), .A2(n1259), .B1(ram[4621]), .B2(n1260), 
        .ZN(n8862) );
  MOAI22 U17784 ( .A1(n27722), .A2(n1259), .B1(ram[4622]), .B2(n1260), 
        .ZN(n8863) );
  MOAI22 U17785 ( .A1(n27487), .A2(n1259), .B1(ram[4623]), .B2(n1260), 
        .ZN(n8864) );
  MOAI22 U17786 ( .A1(n29132), .A2(n1261), .B1(ram[4624]), .B2(n1262), 
        .ZN(n8865) );
  MOAI22 U17787 ( .A1(n28897), .A2(n1261), .B1(ram[4625]), .B2(n1262), 
        .ZN(n8866) );
  MOAI22 U17788 ( .A1(n28662), .A2(n1261), .B1(ram[4626]), .B2(n1262), 
        .ZN(n8867) );
  MOAI22 U17789 ( .A1(n28427), .A2(n1261), .B1(ram[4627]), .B2(n1262), 
        .ZN(n8868) );
  MOAI22 U17790 ( .A1(n28192), .A2(n1261), .B1(ram[4628]), .B2(n1262), 
        .ZN(n8869) );
  MOAI22 U17791 ( .A1(n27957), .A2(n1261), .B1(ram[4629]), .B2(n1262), 
        .ZN(n8870) );
  MOAI22 U17792 ( .A1(n27722), .A2(n1261), .B1(ram[4630]), .B2(n1262), 
        .ZN(n8871) );
  MOAI22 U17793 ( .A1(n27487), .A2(n1261), .B1(ram[4631]), .B2(n1262), 
        .ZN(n8872) );
  MOAI22 U17794 ( .A1(n29132), .A2(n1263), .B1(ram[4632]), .B2(n1264), 
        .ZN(n8873) );
  MOAI22 U17795 ( .A1(n28897), .A2(n1263), .B1(ram[4633]), .B2(n1264), 
        .ZN(n8874) );
  MOAI22 U17796 ( .A1(n28662), .A2(n1263), .B1(ram[4634]), .B2(n1264), 
        .ZN(n8875) );
  MOAI22 U17797 ( .A1(n28427), .A2(n1263), .B1(ram[4635]), .B2(n1264), 
        .ZN(n8876) );
  MOAI22 U17798 ( .A1(n28192), .A2(n1263), .B1(ram[4636]), .B2(n1264), 
        .ZN(n8877) );
  MOAI22 U17799 ( .A1(n27957), .A2(n1263), .B1(ram[4637]), .B2(n1264), 
        .ZN(n8878) );
  MOAI22 U17800 ( .A1(n27722), .A2(n1263), .B1(ram[4638]), .B2(n1264), 
        .ZN(n8879) );
  MOAI22 U17801 ( .A1(n27487), .A2(n1263), .B1(ram[4639]), .B2(n1264), 
        .ZN(n8880) );
  MOAI22 U17802 ( .A1(n29132), .A2(n1265), .B1(ram[4640]), .B2(n1266), 
        .ZN(n8881) );
  MOAI22 U17803 ( .A1(n28897), .A2(n1265), .B1(ram[4641]), .B2(n1266), 
        .ZN(n8882) );
  MOAI22 U17804 ( .A1(n28662), .A2(n1265), .B1(ram[4642]), .B2(n1266), 
        .ZN(n8883) );
  MOAI22 U17805 ( .A1(n28427), .A2(n1265), .B1(ram[4643]), .B2(n1266), 
        .ZN(n8884) );
  MOAI22 U17806 ( .A1(n28192), .A2(n1265), .B1(ram[4644]), .B2(n1266), 
        .ZN(n8885) );
  MOAI22 U17807 ( .A1(n27957), .A2(n1265), .B1(ram[4645]), .B2(n1266), 
        .ZN(n8886) );
  MOAI22 U17808 ( .A1(n27722), .A2(n1265), .B1(ram[4646]), .B2(n1266), 
        .ZN(n8887) );
  MOAI22 U17809 ( .A1(n27487), .A2(n1265), .B1(ram[4647]), .B2(n1266), 
        .ZN(n8888) );
  MOAI22 U17810 ( .A1(n29132), .A2(n1267), .B1(ram[4648]), .B2(n1268), 
        .ZN(n8889) );
  MOAI22 U17811 ( .A1(n28897), .A2(n1267), .B1(ram[4649]), .B2(n1268), 
        .ZN(n8890) );
  MOAI22 U17812 ( .A1(n28662), .A2(n1267), .B1(ram[4650]), .B2(n1268), 
        .ZN(n8891) );
  MOAI22 U17813 ( .A1(n28427), .A2(n1267), .B1(ram[4651]), .B2(n1268), 
        .ZN(n8892) );
  MOAI22 U17814 ( .A1(n28192), .A2(n1267), .B1(ram[4652]), .B2(n1268), 
        .ZN(n8893) );
  MOAI22 U17815 ( .A1(n27957), .A2(n1267), .B1(ram[4653]), .B2(n1268), 
        .ZN(n8894) );
  MOAI22 U17816 ( .A1(n27722), .A2(n1267), .B1(ram[4654]), .B2(n1268), 
        .ZN(n8895) );
  MOAI22 U17817 ( .A1(n27487), .A2(n1267), .B1(ram[4655]), .B2(n1268), 
        .ZN(n8896) );
  MOAI22 U17818 ( .A1(n29132), .A2(n1269), .B1(ram[4656]), .B2(n1270), 
        .ZN(n8897) );
  MOAI22 U17819 ( .A1(n28897), .A2(n1269), .B1(ram[4657]), .B2(n1270), 
        .ZN(n8898) );
  MOAI22 U17820 ( .A1(n28662), .A2(n1269), .B1(ram[4658]), .B2(n1270), 
        .ZN(n8899) );
  MOAI22 U17821 ( .A1(n28427), .A2(n1269), .B1(ram[4659]), .B2(n1270), 
        .ZN(n8900) );
  MOAI22 U17822 ( .A1(n28192), .A2(n1269), .B1(ram[4660]), .B2(n1270), 
        .ZN(n8901) );
  MOAI22 U17823 ( .A1(n27957), .A2(n1269), .B1(ram[4661]), .B2(n1270), 
        .ZN(n8902) );
  MOAI22 U17824 ( .A1(n27722), .A2(n1269), .B1(ram[4662]), .B2(n1270), 
        .ZN(n8903) );
  MOAI22 U17825 ( .A1(n27487), .A2(n1269), .B1(ram[4663]), .B2(n1270), 
        .ZN(n8904) );
  MOAI22 U17826 ( .A1(n29132), .A2(n1271), .B1(ram[4664]), .B2(n1272), 
        .ZN(n8905) );
  MOAI22 U17827 ( .A1(n28897), .A2(n1271), .B1(ram[4665]), .B2(n1272), 
        .ZN(n8906) );
  MOAI22 U17828 ( .A1(n28662), .A2(n1271), .B1(ram[4666]), .B2(n1272), 
        .ZN(n8907) );
  MOAI22 U17829 ( .A1(n28427), .A2(n1271), .B1(ram[4667]), .B2(n1272), 
        .ZN(n8908) );
  MOAI22 U17830 ( .A1(n28192), .A2(n1271), .B1(ram[4668]), .B2(n1272), 
        .ZN(n8909) );
  MOAI22 U17831 ( .A1(n27957), .A2(n1271), .B1(ram[4669]), .B2(n1272), 
        .ZN(n8910) );
  MOAI22 U17832 ( .A1(n27722), .A2(n1271), .B1(ram[4670]), .B2(n1272), 
        .ZN(n8911) );
  MOAI22 U17833 ( .A1(n27487), .A2(n1271), .B1(ram[4671]), .B2(n1272), 
        .ZN(n8912) );
  MOAI22 U17834 ( .A1(n29132), .A2(n1273), .B1(ram[4672]), .B2(n1274), 
        .ZN(n8913) );
  MOAI22 U17835 ( .A1(n28897), .A2(n1273), .B1(ram[4673]), .B2(n1274), 
        .ZN(n8914) );
  MOAI22 U17836 ( .A1(n28662), .A2(n1273), .B1(ram[4674]), .B2(n1274), 
        .ZN(n8915) );
  MOAI22 U17837 ( .A1(n28427), .A2(n1273), .B1(ram[4675]), .B2(n1274), 
        .ZN(n8916) );
  MOAI22 U17838 ( .A1(n28192), .A2(n1273), .B1(ram[4676]), .B2(n1274), 
        .ZN(n8917) );
  MOAI22 U17839 ( .A1(n27957), .A2(n1273), .B1(ram[4677]), .B2(n1274), 
        .ZN(n8918) );
  MOAI22 U17840 ( .A1(n27722), .A2(n1273), .B1(ram[4678]), .B2(n1274), 
        .ZN(n8919) );
  MOAI22 U17841 ( .A1(n27487), .A2(n1273), .B1(ram[4679]), .B2(n1274), 
        .ZN(n8920) );
  MOAI22 U17842 ( .A1(n29133), .A2(n1275), .B1(ram[4680]), .B2(n1276), 
        .ZN(n8921) );
  MOAI22 U17843 ( .A1(n28898), .A2(n1275), .B1(ram[4681]), .B2(n1276), 
        .ZN(n8922) );
  MOAI22 U17844 ( .A1(n28663), .A2(n1275), .B1(ram[4682]), .B2(n1276), 
        .ZN(n8923) );
  MOAI22 U17845 ( .A1(n28428), .A2(n1275), .B1(ram[4683]), .B2(n1276), 
        .ZN(n8924) );
  MOAI22 U17846 ( .A1(n28193), .A2(n1275), .B1(ram[4684]), .B2(n1276), 
        .ZN(n8925) );
  MOAI22 U17847 ( .A1(n27958), .A2(n1275), .B1(ram[4685]), .B2(n1276), 
        .ZN(n8926) );
  MOAI22 U17848 ( .A1(n27723), .A2(n1275), .B1(ram[4686]), .B2(n1276), 
        .ZN(n8927) );
  MOAI22 U17849 ( .A1(n27488), .A2(n1275), .B1(ram[4687]), .B2(n1276), 
        .ZN(n8928) );
  MOAI22 U17850 ( .A1(n29133), .A2(n1277), .B1(ram[4688]), .B2(n1278), 
        .ZN(n8929) );
  MOAI22 U17851 ( .A1(n28898), .A2(n1277), .B1(ram[4689]), .B2(n1278), 
        .ZN(n8930) );
  MOAI22 U17852 ( .A1(n28663), .A2(n1277), .B1(ram[4690]), .B2(n1278), 
        .ZN(n8931) );
  MOAI22 U17853 ( .A1(n28428), .A2(n1277), .B1(ram[4691]), .B2(n1278), 
        .ZN(n8932) );
  MOAI22 U17854 ( .A1(n28193), .A2(n1277), .B1(ram[4692]), .B2(n1278), 
        .ZN(n8933) );
  MOAI22 U17855 ( .A1(n27958), .A2(n1277), .B1(ram[4693]), .B2(n1278), 
        .ZN(n8934) );
  MOAI22 U17856 ( .A1(n27723), .A2(n1277), .B1(ram[4694]), .B2(n1278), 
        .ZN(n8935) );
  MOAI22 U17857 ( .A1(n27488), .A2(n1277), .B1(ram[4695]), .B2(n1278), 
        .ZN(n8936) );
  MOAI22 U17858 ( .A1(n29133), .A2(n1279), .B1(ram[4696]), .B2(n1280), 
        .ZN(n8937) );
  MOAI22 U17859 ( .A1(n28898), .A2(n1279), .B1(ram[4697]), .B2(n1280), 
        .ZN(n8938) );
  MOAI22 U17860 ( .A1(n28663), .A2(n1279), .B1(ram[4698]), .B2(n1280), 
        .ZN(n8939) );
  MOAI22 U17861 ( .A1(n28428), .A2(n1279), .B1(ram[4699]), .B2(n1280), 
        .ZN(n8940) );
  MOAI22 U17862 ( .A1(n28193), .A2(n1279), .B1(ram[4700]), .B2(n1280), 
        .ZN(n8941) );
  MOAI22 U17863 ( .A1(n27958), .A2(n1279), .B1(ram[4701]), .B2(n1280), 
        .ZN(n8942) );
  MOAI22 U17864 ( .A1(n27723), .A2(n1279), .B1(ram[4702]), .B2(n1280), 
        .ZN(n8943) );
  MOAI22 U17865 ( .A1(n27488), .A2(n1279), .B1(ram[4703]), .B2(n1280), 
        .ZN(n8944) );
  MOAI22 U17866 ( .A1(n29133), .A2(n1281), .B1(ram[4704]), .B2(n1282), 
        .ZN(n8945) );
  MOAI22 U17867 ( .A1(n28898), .A2(n1281), .B1(ram[4705]), .B2(n1282), 
        .ZN(n8946) );
  MOAI22 U17868 ( .A1(n28663), .A2(n1281), .B1(ram[4706]), .B2(n1282), 
        .ZN(n8947) );
  MOAI22 U17869 ( .A1(n28428), .A2(n1281), .B1(ram[4707]), .B2(n1282), 
        .ZN(n8948) );
  MOAI22 U17870 ( .A1(n28193), .A2(n1281), .B1(ram[4708]), .B2(n1282), 
        .ZN(n8949) );
  MOAI22 U17871 ( .A1(n27958), .A2(n1281), .B1(ram[4709]), .B2(n1282), 
        .ZN(n8950) );
  MOAI22 U17872 ( .A1(n27723), .A2(n1281), .B1(ram[4710]), .B2(n1282), 
        .ZN(n8951) );
  MOAI22 U17873 ( .A1(n27488), .A2(n1281), .B1(ram[4711]), .B2(n1282), 
        .ZN(n8952) );
  MOAI22 U17874 ( .A1(n29133), .A2(n1283), .B1(ram[4712]), .B2(n1284), 
        .ZN(n8953) );
  MOAI22 U17875 ( .A1(n28898), .A2(n1283), .B1(ram[4713]), .B2(n1284), 
        .ZN(n8954) );
  MOAI22 U17876 ( .A1(n28663), .A2(n1283), .B1(ram[4714]), .B2(n1284), 
        .ZN(n8955) );
  MOAI22 U17877 ( .A1(n28428), .A2(n1283), .B1(ram[4715]), .B2(n1284), 
        .ZN(n8956) );
  MOAI22 U17878 ( .A1(n28193), .A2(n1283), .B1(ram[4716]), .B2(n1284), 
        .ZN(n8957) );
  MOAI22 U17879 ( .A1(n27958), .A2(n1283), .B1(ram[4717]), .B2(n1284), 
        .ZN(n8958) );
  MOAI22 U17880 ( .A1(n27723), .A2(n1283), .B1(ram[4718]), .B2(n1284), 
        .ZN(n8959) );
  MOAI22 U17881 ( .A1(n27488), .A2(n1283), .B1(ram[4719]), .B2(n1284), 
        .ZN(n8960) );
  MOAI22 U17882 ( .A1(n29133), .A2(n1285), .B1(ram[4720]), .B2(n1286), 
        .ZN(n8961) );
  MOAI22 U17883 ( .A1(n28898), .A2(n1285), .B1(ram[4721]), .B2(n1286), 
        .ZN(n8962) );
  MOAI22 U17884 ( .A1(n28663), .A2(n1285), .B1(ram[4722]), .B2(n1286), 
        .ZN(n8963) );
  MOAI22 U17885 ( .A1(n28428), .A2(n1285), .B1(ram[4723]), .B2(n1286), 
        .ZN(n8964) );
  MOAI22 U17886 ( .A1(n28193), .A2(n1285), .B1(ram[4724]), .B2(n1286), 
        .ZN(n8965) );
  MOAI22 U17887 ( .A1(n27958), .A2(n1285), .B1(ram[4725]), .B2(n1286), 
        .ZN(n8966) );
  MOAI22 U17888 ( .A1(n27723), .A2(n1285), .B1(ram[4726]), .B2(n1286), 
        .ZN(n8967) );
  MOAI22 U17889 ( .A1(n27488), .A2(n1285), .B1(ram[4727]), .B2(n1286), 
        .ZN(n8968) );
  MOAI22 U17890 ( .A1(n29133), .A2(n1287), .B1(ram[4728]), .B2(n1288), 
        .ZN(n8969) );
  MOAI22 U17891 ( .A1(n28898), .A2(n1287), .B1(ram[4729]), .B2(n1288), 
        .ZN(n8970) );
  MOAI22 U17892 ( .A1(n28663), .A2(n1287), .B1(ram[4730]), .B2(n1288), 
        .ZN(n8971) );
  MOAI22 U17893 ( .A1(n28428), .A2(n1287), .B1(ram[4731]), .B2(n1288), 
        .ZN(n8972) );
  MOAI22 U17894 ( .A1(n28193), .A2(n1287), .B1(ram[4732]), .B2(n1288), 
        .ZN(n8973) );
  MOAI22 U17895 ( .A1(n27958), .A2(n1287), .B1(ram[4733]), .B2(n1288), 
        .ZN(n8974) );
  MOAI22 U17896 ( .A1(n27723), .A2(n1287), .B1(ram[4734]), .B2(n1288), 
        .ZN(n8975) );
  MOAI22 U17897 ( .A1(n27488), .A2(n1287), .B1(ram[4735]), .B2(n1288), 
        .ZN(n8976) );
  MOAI22 U17898 ( .A1(n29133), .A2(n1289), .B1(ram[4736]), .B2(n1290), 
        .ZN(n8977) );
  MOAI22 U17899 ( .A1(n28898), .A2(n1289), .B1(ram[4737]), .B2(n1290), 
        .ZN(n8978) );
  MOAI22 U17900 ( .A1(n28663), .A2(n1289), .B1(ram[4738]), .B2(n1290), 
        .ZN(n8979) );
  MOAI22 U17901 ( .A1(n28428), .A2(n1289), .B1(ram[4739]), .B2(n1290), 
        .ZN(n8980) );
  MOAI22 U17902 ( .A1(n28193), .A2(n1289), .B1(ram[4740]), .B2(n1290), 
        .ZN(n8981) );
  MOAI22 U17903 ( .A1(n27958), .A2(n1289), .B1(ram[4741]), .B2(n1290), 
        .ZN(n8982) );
  MOAI22 U17904 ( .A1(n27723), .A2(n1289), .B1(ram[4742]), .B2(n1290), 
        .ZN(n8983) );
  MOAI22 U17905 ( .A1(n27488), .A2(n1289), .B1(ram[4743]), .B2(n1290), 
        .ZN(n8984) );
  MOAI22 U17906 ( .A1(n29133), .A2(n1291), .B1(ram[4744]), .B2(n1292), 
        .ZN(n8985) );
  MOAI22 U17907 ( .A1(n28898), .A2(n1291), .B1(ram[4745]), .B2(n1292), 
        .ZN(n8986) );
  MOAI22 U17908 ( .A1(n28663), .A2(n1291), .B1(ram[4746]), .B2(n1292), 
        .ZN(n8987) );
  MOAI22 U17909 ( .A1(n28428), .A2(n1291), .B1(ram[4747]), .B2(n1292), 
        .ZN(n8988) );
  MOAI22 U17910 ( .A1(n28193), .A2(n1291), .B1(ram[4748]), .B2(n1292), 
        .ZN(n8989) );
  MOAI22 U17911 ( .A1(n27958), .A2(n1291), .B1(ram[4749]), .B2(n1292), 
        .ZN(n8990) );
  MOAI22 U17912 ( .A1(n27723), .A2(n1291), .B1(ram[4750]), .B2(n1292), 
        .ZN(n8991) );
  MOAI22 U17913 ( .A1(n27488), .A2(n1291), .B1(ram[4751]), .B2(n1292), 
        .ZN(n8992) );
  MOAI22 U17914 ( .A1(n29133), .A2(n1293), .B1(ram[4752]), .B2(n1294), 
        .ZN(n8993) );
  MOAI22 U17915 ( .A1(n28898), .A2(n1293), .B1(ram[4753]), .B2(n1294), 
        .ZN(n8994) );
  MOAI22 U17916 ( .A1(n28663), .A2(n1293), .B1(ram[4754]), .B2(n1294), 
        .ZN(n8995) );
  MOAI22 U17917 ( .A1(n28428), .A2(n1293), .B1(ram[4755]), .B2(n1294), 
        .ZN(n8996) );
  MOAI22 U17918 ( .A1(n28193), .A2(n1293), .B1(ram[4756]), .B2(n1294), 
        .ZN(n8997) );
  MOAI22 U17919 ( .A1(n27958), .A2(n1293), .B1(ram[4757]), .B2(n1294), 
        .ZN(n8998) );
  MOAI22 U17920 ( .A1(n27723), .A2(n1293), .B1(ram[4758]), .B2(n1294), 
        .ZN(n8999) );
  MOAI22 U17921 ( .A1(n27488), .A2(n1293), .B1(ram[4759]), .B2(n1294), 
        .ZN(n9000) );
  MOAI22 U17922 ( .A1(n29133), .A2(n1295), .B1(ram[4760]), .B2(n1296), 
        .ZN(n9001) );
  MOAI22 U17923 ( .A1(n28898), .A2(n1295), .B1(ram[4761]), .B2(n1296), 
        .ZN(n9002) );
  MOAI22 U17924 ( .A1(n28663), .A2(n1295), .B1(ram[4762]), .B2(n1296), 
        .ZN(n9003) );
  MOAI22 U17925 ( .A1(n28428), .A2(n1295), .B1(ram[4763]), .B2(n1296), 
        .ZN(n9004) );
  MOAI22 U17926 ( .A1(n28193), .A2(n1295), .B1(ram[4764]), .B2(n1296), 
        .ZN(n9005) );
  MOAI22 U17927 ( .A1(n27958), .A2(n1295), .B1(ram[4765]), .B2(n1296), 
        .ZN(n9006) );
  MOAI22 U17928 ( .A1(n27723), .A2(n1295), .B1(ram[4766]), .B2(n1296), 
        .ZN(n9007) );
  MOAI22 U17929 ( .A1(n27488), .A2(n1295), .B1(ram[4767]), .B2(n1296), 
        .ZN(n9008) );
  MOAI22 U17930 ( .A1(n29133), .A2(n1297), .B1(ram[4768]), .B2(n1298), 
        .ZN(n9009) );
  MOAI22 U17931 ( .A1(n28898), .A2(n1297), .B1(ram[4769]), .B2(n1298), 
        .ZN(n9010) );
  MOAI22 U17932 ( .A1(n28663), .A2(n1297), .B1(ram[4770]), .B2(n1298), 
        .ZN(n9011) );
  MOAI22 U17933 ( .A1(n28428), .A2(n1297), .B1(ram[4771]), .B2(n1298), 
        .ZN(n9012) );
  MOAI22 U17934 ( .A1(n28193), .A2(n1297), .B1(ram[4772]), .B2(n1298), 
        .ZN(n9013) );
  MOAI22 U17935 ( .A1(n27958), .A2(n1297), .B1(ram[4773]), .B2(n1298), 
        .ZN(n9014) );
  MOAI22 U17936 ( .A1(n27723), .A2(n1297), .B1(ram[4774]), .B2(n1298), 
        .ZN(n9015) );
  MOAI22 U17937 ( .A1(n27488), .A2(n1297), .B1(ram[4775]), .B2(n1298), 
        .ZN(n9016) );
  MOAI22 U17938 ( .A1(n29133), .A2(n1299), .B1(ram[4776]), .B2(n1300), 
        .ZN(n9017) );
  MOAI22 U17939 ( .A1(n28898), .A2(n1299), .B1(ram[4777]), .B2(n1300), 
        .ZN(n9018) );
  MOAI22 U17940 ( .A1(n28663), .A2(n1299), .B1(ram[4778]), .B2(n1300), 
        .ZN(n9019) );
  MOAI22 U17941 ( .A1(n28428), .A2(n1299), .B1(ram[4779]), .B2(n1300), 
        .ZN(n9020) );
  MOAI22 U17942 ( .A1(n28193), .A2(n1299), .B1(ram[4780]), .B2(n1300), 
        .ZN(n9021) );
  MOAI22 U17943 ( .A1(n27958), .A2(n1299), .B1(ram[4781]), .B2(n1300), 
        .ZN(n9022) );
  MOAI22 U17944 ( .A1(n27723), .A2(n1299), .B1(ram[4782]), .B2(n1300), 
        .ZN(n9023) );
  MOAI22 U17945 ( .A1(n27488), .A2(n1299), .B1(ram[4783]), .B2(n1300), 
        .ZN(n9024) );
  MOAI22 U17946 ( .A1(n29134), .A2(n1301), .B1(ram[4784]), .B2(n1302), 
        .ZN(n9025) );
  MOAI22 U17947 ( .A1(n28899), .A2(n1301), .B1(ram[4785]), .B2(n1302), 
        .ZN(n9026) );
  MOAI22 U17948 ( .A1(n28664), .A2(n1301), .B1(ram[4786]), .B2(n1302), 
        .ZN(n9027) );
  MOAI22 U17949 ( .A1(n28429), .A2(n1301), .B1(ram[4787]), .B2(n1302), 
        .ZN(n9028) );
  MOAI22 U17950 ( .A1(n28194), .A2(n1301), .B1(ram[4788]), .B2(n1302), 
        .ZN(n9029) );
  MOAI22 U17951 ( .A1(n27959), .A2(n1301), .B1(ram[4789]), .B2(n1302), 
        .ZN(n9030) );
  MOAI22 U17952 ( .A1(n27724), .A2(n1301), .B1(ram[4790]), .B2(n1302), 
        .ZN(n9031) );
  MOAI22 U17953 ( .A1(n27489), .A2(n1301), .B1(ram[4791]), .B2(n1302), 
        .ZN(n9032) );
  MOAI22 U17954 ( .A1(n29134), .A2(n1303), .B1(ram[4792]), .B2(n1304), 
        .ZN(n9033) );
  MOAI22 U17955 ( .A1(n28899), .A2(n1303), .B1(ram[4793]), .B2(n1304), 
        .ZN(n9034) );
  MOAI22 U17956 ( .A1(n28664), .A2(n1303), .B1(ram[4794]), .B2(n1304), 
        .ZN(n9035) );
  MOAI22 U17957 ( .A1(n28429), .A2(n1303), .B1(ram[4795]), .B2(n1304), 
        .ZN(n9036) );
  MOAI22 U17958 ( .A1(n28194), .A2(n1303), .B1(ram[4796]), .B2(n1304), 
        .ZN(n9037) );
  MOAI22 U17959 ( .A1(n27959), .A2(n1303), .B1(ram[4797]), .B2(n1304), 
        .ZN(n9038) );
  MOAI22 U17960 ( .A1(n27724), .A2(n1303), .B1(ram[4798]), .B2(n1304), 
        .ZN(n9039) );
  MOAI22 U17961 ( .A1(n27489), .A2(n1303), .B1(ram[4799]), .B2(n1304), 
        .ZN(n9040) );
  MOAI22 U17962 ( .A1(n29134), .A2(n1305), .B1(ram[4800]), .B2(n1306), 
        .ZN(n9041) );
  MOAI22 U17963 ( .A1(n28899), .A2(n1305), .B1(ram[4801]), .B2(n1306), 
        .ZN(n9042) );
  MOAI22 U17964 ( .A1(n28664), .A2(n1305), .B1(ram[4802]), .B2(n1306), 
        .ZN(n9043) );
  MOAI22 U17965 ( .A1(n28429), .A2(n1305), .B1(ram[4803]), .B2(n1306), 
        .ZN(n9044) );
  MOAI22 U17966 ( .A1(n28194), .A2(n1305), .B1(ram[4804]), .B2(n1306), 
        .ZN(n9045) );
  MOAI22 U17967 ( .A1(n27959), .A2(n1305), .B1(ram[4805]), .B2(n1306), 
        .ZN(n9046) );
  MOAI22 U17968 ( .A1(n27724), .A2(n1305), .B1(ram[4806]), .B2(n1306), 
        .ZN(n9047) );
  MOAI22 U17969 ( .A1(n27489), .A2(n1305), .B1(ram[4807]), .B2(n1306), 
        .ZN(n9048) );
  MOAI22 U17970 ( .A1(n29134), .A2(n1307), .B1(ram[4808]), .B2(n1308), 
        .ZN(n9049) );
  MOAI22 U17971 ( .A1(n28899), .A2(n1307), .B1(ram[4809]), .B2(n1308), 
        .ZN(n9050) );
  MOAI22 U17972 ( .A1(n28664), .A2(n1307), .B1(ram[4810]), .B2(n1308), 
        .ZN(n9051) );
  MOAI22 U17973 ( .A1(n28429), .A2(n1307), .B1(ram[4811]), .B2(n1308), 
        .ZN(n9052) );
  MOAI22 U17974 ( .A1(n28194), .A2(n1307), .B1(ram[4812]), .B2(n1308), 
        .ZN(n9053) );
  MOAI22 U17975 ( .A1(n27959), .A2(n1307), .B1(ram[4813]), .B2(n1308), 
        .ZN(n9054) );
  MOAI22 U17976 ( .A1(n27724), .A2(n1307), .B1(ram[4814]), .B2(n1308), 
        .ZN(n9055) );
  MOAI22 U17977 ( .A1(n27489), .A2(n1307), .B1(ram[4815]), .B2(n1308), 
        .ZN(n9056) );
  MOAI22 U17978 ( .A1(n29134), .A2(n1309), .B1(ram[4816]), .B2(n1310), 
        .ZN(n9057) );
  MOAI22 U17979 ( .A1(n28899), .A2(n1309), .B1(ram[4817]), .B2(n1310), 
        .ZN(n9058) );
  MOAI22 U17980 ( .A1(n28664), .A2(n1309), .B1(ram[4818]), .B2(n1310), 
        .ZN(n9059) );
  MOAI22 U17981 ( .A1(n28429), .A2(n1309), .B1(ram[4819]), .B2(n1310), 
        .ZN(n9060) );
  MOAI22 U17982 ( .A1(n28194), .A2(n1309), .B1(ram[4820]), .B2(n1310), 
        .ZN(n9061) );
  MOAI22 U17983 ( .A1(n27959), .A2(n1309), .B1(ram[4821]), .B2(n1310), 
        .ZN(n9062) );
  MOAI22 U17984 ( .A1(n27724), .A2(n1309), .B1(ram[4822]), .B2(n1310), 
        .ZN(n9063) );
  MOAI22 U17985 ( .A1(n27489), .A2(n1309), .B1(ram[4823]), .B2(n1310), 
        .ZN(n9064) );
  MOAI22 U17986 ( .A1(n29134), .A2(n1311), .B1(ram[4824]), .B2(n1312), 
        .ZN(n9065) );
  MOAI22 U17987 ( .A1(n28899), .A2(n1311), .B1(ram[4825]), .B2(n1312), 
        .ZN(n9066) );
  MOAI22 U17988 ( .A1(n28664), .A2(n1311), .B1(ram[4826]), .B2(n1312), 
        .ZN(n9067) );
  MOAI22 U17989 ( .A1(n28429), .A2(n1311), .B1(ram[4827]), .B2(n1312), 
        .ZN(n9068) );
  MOAI22 U17990 ( .A1(n28194), .A2(n1311), .B1(ram[4828]), .B2(n1312), 
        .ZN(n9069) );
  MOAI22 U17991 ( .A1(n27959), .A2(n1311), .B1(ram[4829]), .B2(n1312), 
        .ZN(n9070) );
  MOAI22 U17992 ( .A1(n27724), .A2(n1311), .B1(ram[4830]), .B2(n1312), 
        .ZN(n9071) );
  MOAI22 U17993 ( .A1(n27489), .A2(n1311), .B1(ram[4831]), .B2(n1312), 
        .ZN(n9072) );
  MOAI22 U17994 ( .A1(n29134), .A2(n1313), .B1(ram[4832]), .B2(n1314), 
        .ZN(n9073) );
  MOAI22 U17995 ( .A1(n28899), .A2(n1313), .B1(ram[4833]), .B2(n1314), 
        .ZN(n9074) );
  MOAI22 U17996 ( .A1(n28664), .A2(n1313), .B1(ram[4834]), .B2(n1314), 
        .ZN(n9075) );
  MOAI22 U17997 ( .A1(n28429), .A2(n1313), .B1(ram[4835]), .B2(n1314), 
        .ZN(n9076) );
  MOAI22 U17998 ( .A1(n28194), .A2(n1313), .B1(ram[4836]), .B2(n1314), 
        .ZN(n9077) );
  MOAI22 U17999 ( .A1(n27959), .A2(n1313), .B1(ram[4837]), .B2(n1314), 
        .ZN(n9078) );
  MOAI22 U18000 ( .A1(n27724), .A2(n1313), .B1(ram[4838]), .B2(n1314), 
        .ZN(n9079) );
  MOAI22 U18001 ( .A1(n27489), .A2(n1313), .B1(ram[4839]), .B2(n1314), 
        .ZN(n9080) );
  MOAI22 U18002 ( .A1(n29134), .A2(n1315), .B1(ram[4840]), .B2(n1316), 
        .ZN(n9081) );
  MOAI22 U18003 ( .A1(n28899), .A2(n1315), .B1(ram[4841]), .B2(n1316), 
        .ZN(n9082) );
  MOAI22 U18004 ( .A1(n28664), .A2(n1315), .B1(ram[4842]), .B2(n1316), 
        .ZN(n9083) );
  MOAI22 U18005 ( .A1(n28429), .A2(n1315), .B1(ram[4843]), .B2(n1316), 
        .ZN(n9084) );
  MOAI22 U18006 ( .A1(n28194), .A2(n1315), .B1(ram[4844]), .B2(n1316), 
        .ZN(n9085) );
  MOAI22 U18007 ( .A1(n27959), .A2(n1315), .B1(ram[4845]), .B2(n1316), 
        .ZN(n9086) );
  MOAI22 U18008 ( .A1(n27724), .A2(n1315), .B1(ram[4846]), .B2(n1316), 
        .ZN(n9087) );
  MOAI22 U18009 ( .A1(n27489), .A2(n1315), .B1(ram[4847]), .B2(n1316), 
        .ZN(n9088) );
  MOAI22 U18010 ( .A1(n29134), .A2(n1317), .B1(ram[4848]), .B2(n1318), 
        .ZN(n9089) );
  MOAI22 U18011 ( .A1(n28899), .A2(n1317), .B1(ram[4849]), .B2(n1318), 
        .ZN(n9090) );
  MOAI22 U18012 ( .A1(n28664), .A2(n1317), .B1(ram[4850]), .B2(n1318), 
        .ZN(n9091) );
  MOAI22 U18013 ( .A1(n28429), .A2(n1317), .B1(ram[4851]), .B2(n1318), 
        .ZN(n9092) );
  MOAI22 U18014 ( .A1(n28194), .A2(n1317), .B1(ram[4852]), .B2(n1318), 
        .ZN(n9093) );
  MOAI22 U18015 ( .A1(n27959), .A2(n1317), .B1(ram[4853]), .B2(n1318), 
        .ZN(n9094) );
  MOAI22 U18016 ( .A1(n27724), .A2(n1317), .B1(ram[4854]), .B2(n1318), 
        .ZN(n9095) );
  MOAI22 U18017 ( .A1(n27489), .A2(n1317), .B1(ram[4855]), .B2(n1318), 
        .ZN(n9096) );
  MOAI22 U18018 ( .A1(n29134), .A2(n1319), .B1(ram[4856]), .B2(n1320), 
        .ZN(n9097) );
  MOAI22 U18019 ( .A1(n28899), .A2(n1319), .B1(ram[4857]), .B2(n1320), 
        .ZN(n9098) );
  MOAI22 U18020 ( .A1(n28664), .A2(n1319), .B1(ram[4858]), .B2(n1320), 
        .ZN(n9099) );
  MOAI22 U18021 ( .A1(n28429), .A2(n1319), .B1(ram[4859]), .B2(n1320), 
        .ZN(n9100) );
  MOAI22 U18022 ( .A1(n28194), .A2(n1319), .B1(ram[4860]), .B2(n1320), 
        .ZN(n9101) );
  MOAI22 U18023 ( .A1(n27959), .A2(n1319), .B1(ram[4861]), .B2(n1320), 
        .ZN(n9102) );
  MOAI22 U18024 ( .A1(n27724), .A2(n1319), .B1(ram[4862]), .B2(n1320), 
        .ZN(n9103) );
  MOAI22 U18025 ( .A1(n27489), .A2(n1319), .B1(ram[4863]), .B2(n1320), 
        .ZN(n9104) );
  MOAI22 U18026 ( .A1(n29134), .A2(n1321), .B1(ram[4864]), .B2(n1322), 
        .ZN(n9105) );
  MOAI22 U18027 ( .A1(n28899), .A2(n1321), .B1(ram[4865]), .B2(n1322), 
        .ZN(n9106) );
  MOAI22 U18028 ( .A1(n28664), .A2(n1321), .B1(ram[4866]), .B2(n1322), 
        .ZN(n9107) );
  MOAI22 U18029 ( .A1(n28429), .A2(n1321), .B1(ram[4867]), .B2(n1322), 
        .ZN(n9108) );
  MOAI22 U18030 ( .A1(n28194), .A2(n1321), .B1(ram[4868]), .B2(n1322), 
        .ZN(n9109) );
  MOAI22 U18031 ( .A1(n27959), .A2(n1321), .B1(ram[4869]), .B2(n1322), 
        .ZN(n9110) );
  MOAI22 U18032 ( .A1(n27724), .A2(n1321), .B1(ram[4870]), .B2(n1322), 
        .ZN(n9111) );
  MOAI22 U18033 ( .A1(n27489), .A2(n1321), .B1(ram[4871]), .B2(n1322), 
        .ZN(n9112) );
  MOAI22 U18034 ( .A1(n29134), .A2(n1323), .B1(ram[4872]), .B2(n1324), 
        .ZN(n9113) );
  MOAI22 U18035 ( .A1(n28899), .A2(n1323), .B1(ram[4873]), .B2(n1324), 
        .ZN(n9114) );
  MOAI22 U18036 ( .A1(n28664), .A2(n1323), .B1(ram[4874]), .B2(n1324), 
        .ZN(n9115) );
  MOAI22 U18037 ( .A1(n28429), .A2(n1323), .B1(ram[4875]), .B2(n1324), 
        .ZN(n9116) );
  MOAI22 U18038 ( .A1(n28194), .A2(n1323), .B1(ram[4876]), .B2(n1324), 
        .ZN(n9117) );
  MOAI22 U18039 ( .A1(n27959), .A2(n1323), .B1(ram[4877]), .B2(n1324), 
        .ZN(n9118) );
  MOAI22 U18040 ( .A1(n27724), .A2(n1323), .B1(ram[4878]), .B2(n1324), 
        .ZN(n9119) );
  MOAI22 U18041 ( .A1(n27489), .A2(n1323), .B1(ram[4879]), .B2(n1324), 
        .ZN(n9120) );
  MOAI22 U18042 ( .A1(n29134), .A2(n1325), .B1(ram[4880]), .B2(n1326), 
        .ZN(n9121) );
  MOAI22 U18043 ( .A1(n28899), .A2(n1325), .B1(ram[4881]), .B2(n1326), 
        .ZN(n9122) );
  MOAI22 U18044 ( .A1(n28664), .A2(n1325), .B1(ram[4882]), .B2(n1326), 
        .ZN(n9123) );
  MOAI22 U18045 ( .A1(n28429), .A2(n1325), .B1(ram[4883]), .B2(n1326), 
        .ZN(n9124) );
  MOAI22 U18046 ( .A1(n28194), .A2(n1325), .B1(ram[4884]), .B2(n1326), 
        .ZN(n9125) );
  MOAI22 U18047 ( .A1(n27959), .A2(n1325), .B1(ram[4885]), .B2(n1326), 
        .ZN(n9126) );
  MOAI22 U18048 ( .A1(n27724), .A2(n1325), .B1(ram[4886]), .B2(n1326), 
        .ZN(n9127) );
  MOAI22 U18049 ( .A1(n27489), .A2(n1325), .B1(ram[4887]), .B2(n1326), 
        .ZN(n9128) );
  MOAI22 U18050 ( .A1(n29135), .A2(n1327), .B1(ram[4888]), .B2(n1328), 
        .ZN(n9129) );
  MOAI22 U18051 ( .A1(n28900), .A2(n1327), .B1(ram[4889]), .B2(n1328), 
        .ZN(n9130) );
  MOAI22 U18052 ( .A1(n28665), .A2(n1327), .B1(ram[4890]), .B2(n1328), 
        .ZN(n9131) );
  MOAI22 U18053 ( .A1(n28430), .A2(n1327), .B1(ram[4891]), .B2(n1328), 
        .ZN(n9132) );
  MOAI22 U18054 ( .A1(n28195), .A2(n1327), .B1(ram[4892]), .B2(n1328), 
        .ZN(n9133) );
  MOAI22 U18055 ( .A1(n27960), .A2(n1327), .B1(ram[4893]), .B2(n1328), 
        .ZN(n9134) );
  MOAI22 U18056 ( .A1(n27725), .A2(n1327), .B1(ram[4894]), .B2(n1328), 
        .ZN(n9135) );
  MOAI22 U18057 ( .A1(n27490), .A2(n1327), .B1(ram[4895]), .B2(n1328), 
        .ZN(n9136) );
  MOAI22 U18058 ( .A1(n29135), .A2(n1329), .B1(ram[4896]), .B2(n1330), 
        .ZN(n9137) );
  MOAI22 U18059 ( .A1(n28900), .A2(n1329), .B1(ram[4897]), .B2(n1330), 
        .ZN(n9138) );
  MOAI22 U18060 ( .A1(n28665), .A2(n1329), .B1(ram[4898]), .B2(n1330), 
        .ZN(n9139) );
  MOAI22 U18061 ( .A1(n28430), .A2(n1329), .B1(ram[4899]), .B2(n1330), 
        .ZN(n9140) );
  MOAI22 U18062 ( .A1(n28195), .A2(n1329), .B1(ram[4900]), .B2(n1330), 
        .ZN(n9141) );
  MOAI22 U18063 ( .A1(n27960), .A2(n1329), .B1(ram[4901]), .B2(n1330), 
        .ZN(n9142) );
  MOAI22 U18064 ( .A1(n27725), .A2(n1329), .B1(ram[4902]), .B2(n1330), 
        .ZN(n9143) );
  MOAI22 U18065 ( .A1(n27490), .A2(n1329), .B1(ram[4903]), .B2(n1330), 
        .ZN(n9144) );
  MOAI22 U18066 ( .A1(n29135), .A2(n1331), .B1(ram[4904]), .B2(n1332), 
        .ZN(n9145) );
  MOAI22 U18067 ( .A1(n28900), .A2(n1331), .B1(ram[4905]), .B2(n1332), 
        .ZN(n9146) );
  MOAI22 U18068 ( .A1(n28665), .A2(n1331), .B1(ram[4906]), .B2(n1332), 
        .ZN(n9147) );
  MOAI22 U18069 ( .A1(n28430), .A2(n1331), .B1(ram[4907]), .B2(n1332), 
        .ZN(n9148) );
  MOAI22 U18070 ( .A1(n28195), .A2(n1331), .B1(ram[4908]), .B2(n1332), 
        .ZN(n9149) );
  MOAI22 U18071 ( .A1(n27960), .A2(n1331), .B1(ram[4909]), .B2(n1332), 
        .ZN(n9150) );
  MOAI22 U18072 ( .A1(n27725), .A2(n1331), .B1(ram[4910]), .B2(n1332), 
        .ZN(n9151) );
  MOAI22 U18073 ( .A1(n27490), .A2(n1331), .B1(ram[4911]), .B2(n1332), 
        .ZN(n9152) );
  MOAI22 U18074 ( .A1(n29135), .A2(n1333), .B1(ram[4912]), .B2(n1334), 
        .ZN(n9153) );
  MOAI22 U18075 ( .A1(n28900), .A2(n1333), .B1(ram[4913]), .B2(n1334), 
        .ZN(n9154) );
  MOAI22 U18076 ( .A1(n28665), .A2(n1333), .B1(ram[4914]), .B2(n1334), 
        .ZN(n9155) );
  MOAI22 U18077 ( .A1(n28430), .A2(n1333), .B1(ram[4915]), .B2(n1334), 
        .ZN(n9156) );
  MOAI22 U18078 ( .A1(n28195), .A2(n1333), .B1(ram[4916]), .B2(n1334), 
        .ZN(n9157) );
  MOAI22 U18079 ( .A1(n27960), .A2(n1333), .B1(ram[4917]), .B2(n1334), 
        .ZN(n9158) );
  MOAI22 U18080 ( .A1(n27725), .A2(n1333), .B1(ram[4918]), .B2(n1334), 
        .ZN(n9159) );
  MOAI22 U18081 ( .A1(n27490), .A2(n1333), .B1(ram[4919]), .B2(n1334), 
        .ZN(n9160) );
  MOAI22 U18082 ( .A1(n29135), .A2(n1335), .B1(ram[4920]), .B2(n1336), 
        .ZN(n9161) );
  MOAI22 U18083 ( .A1(n28900), .A2(n1335), .B1(ram[4921]), .B2(n1336), 
        .ZN(n9162) );
  MOAI22 U18084 ( .A1(n28665), .A2(n1335), .B1(ram[4922]), .B2(n1336), 
        .ZN(n9163) );
  MOAI22 U18085 ( .A1(n28430), .A2(n1335), .B1(ram[4923]), .B2(n1336), 
        .ZN(n9164) );
  MOAI22 U18086 ( .A1(n28195), .A2(n1335), .B1(ram[4924]), .B2(n1336), 
        .ZN(n9165) );
  MOAI22 U18087 ( .A1(n27960), .A2(n1335), .B1(ram[4925]), .B2(n1336), 
        .ZN(n9166) );
  MOAI22 U18088 ( .A1(n27725), .A2(n1335), .B1(ram[4926]), .B2(n1336), 
        .ZN(n9167) );
  MOAI22 U18089 ( .A1(n27490), .A2(n1335), .B1(ram[4927]), .B2(n1336), 
        .ZN(n9168) );
  MOAI22 U18090 ( .A1(n29135), .A2(n1337), .B1(ram[4928]), .B2(n1338), 
        .ZN(n9169) );
  MOAI22 U18091 ( .A1(n28900), .A2(n1337), .B1(ram[4929]), .B2(n1338), 
        .ZN(n9170) );
  MOAI22 U18092 ( .A1(n28665), .A2(n1337), .B1(ram[4930]), .B2(n1338), 
        .ZN(n9171) );
  MOAI22 U18093 ( .A1(n28430), .A2(n1337), .B1(ram[4931]), .B2(n1338), 
        .ZN(n9172) );
  MOAI22 U18094 ( .A1(n28195), .A2(n1337), .B1(ram[4932]), .B2(n1338), 
        .ZN(n9173) );
  MOAI22 U18095 ( .A1(n27960), .A2(n1337), .B1(ram[4933]), .B2(n1338), 
        .ZN(n9174) );
  MOAI22 U18096 ( .A1(n27725), .A2(n1337), .B1(ram[4934]), .B2(n1338), 
        .ZN(n9175) );
  MOAI22 U18097 ( .A1(n27490), .A2(n1337), .B1(ram[4935]), .B2(n1338), 
        .ZN(n9176) );
  MOAI22 U18098 ( .A1(n29135), .A2(n1339), .B1(ram[4936]), .B2(n1340), 
        .ZN(n9177) );
  MOAI22 U18099 ( .A1(n28900), .A2(n1339), .B1(ram[4937]), .B2(n1340), 
        .ZN(n9178) );
  MOAI22 U18100 ( .A1(n28665), .A2(n1339), .B1(ram[4938]), .B2(n1340), 
        .ZN(n9179) );
  MOAI22 U18101 ( .A1(n28430), .A2(n1339), .B1(ram[4939]), .B2(n1340), 
        .ZN(n9180) );
  MOAI22 U18102 ( .A1(n28195), .A2(n1339), .B1(ram[4940]), .B2(n1340), 
        .ZN(n9181) );
  MOAI22 U18103 ( .A1(n27960), .A2(n1339), .B1(ram[4941]), .B2(n1340), 
        .ZN(n9182) );
  MOAI22 U18104 ( .A1(n27725), .A2(n1339), .B1(ram[4942]), .B2(n1340), 
        .ZN(n9183) );
  MOAI22 U18105 ( .A1(n27490), .A2(n1339), .B1(ram[4943]), .B2(n1340), 
        .ZN(n9184) );
  MOAI22 U18106 ( .A1(n29135), .A2(n1341), .B1(ram[4944]), .B2(n1342), 
        .ZN(n9185) );
  MOAI22 U18107 ( .A1(n28900), .A2(n1341), .B1(ram[4945]), .B2(n1342), 
        .ZN(n9186) );
  MOAI22 U18108 ( .A1(n28665), .A2(n1341), .B1(ram[4946]), .B2(n1342), 
        .ZN(n9187) );
  MOAI22 U18109 ( .A1(n28430), .A2(n1341), .B1(ram[4947]), .B2(n1342), 
        .ZN(n9188) );
  MOAI22 U18110 ( .A1(n28195), .A2(n1341), .B1(ram[4948]), .B2(n1342), 
        .ZN(n9189) );
  MOAI22 U18111 ( .A1(n27960), .A2(n1341), .B1(ram[4949]), .B2(n1342), 
        .ZN(n9190) );
  MOAI22 U18112 ( .A1(n27725), .A2(n1341), .B1(ram[4950]), .B2(n1342), 
        .ZN(n9191) );
  MOAI22 U18113 ( .A1(n27490), .A2(n1341), .B1(ram[4951]), .B2(n1342), 
        .ZN(n9192) );
  MOAI22 U18114 ( .A1(n29135), .A2(n1343), .B1(ram[4952]), .B2(n1344), 
        .ZN(n9193) );
  MOAI22 U18115 ( .A1(n28900), .A2(n1343), .B1(ram[4953]), .B2(n1344), 
        .ZN(n9194) );
  MOAI22 U18116 ( .A1(n28665), .A2(n1343), .B1(ram[4954]), .B2(n1344), 
        .ZN(n9195) );
  MOAI22 U18117 ( .A1(n28430), .A2(n1343), .B1(ram[4955]), .B2(n1344), 
        .ZN(n9196) );
  MOAI22 U18118 ( .A1(n28195), .A2(n1343), .B1(ram[4956]), .B2(n1344), 
        .ZN(n9197) );
  MOAI22 U18119 ( .A1(n27960), .A2(n1343), .B1(ram[4957]), .B2(n1344), 
        .ZN(n9198) );
  MOAI22 U18120 ( .A1(n27725), .A2(n1343), .B1(ram[4958]), .B2(n1344), 
        .ZN(n9199) );
  MOAI22 U18121 ( .A1(n27490), .A2(n1343), .B1(ram[4959]), .B2(n1344), 
        .ZN(n9200) );
  MOAI22 U18122 ( .A1(n29135), .A2(n1345), .B1(ram[4960]), .B2(n1346), 
        .ZN(n9201) );
  MOAI22 U18123 ( .A1(n28900), .A2(n1345), .B1(ram[4961]), .B2(n1346), 
        .ZN(n9202) );
  MOAI22 U18124 ( .A1(n28665), .A2(n1345), .B1(ram[4962]), .B2(n1346), 
        .ZN(n9203) );
  MOAI22 U18125 ( .A1(n28430), .A2(n1345), .B1(ram[4963]), .B2(n1346), 
        .ZN(n9204) );
  MOAI22 U18126 ( .A1(n28195), .A2(n1345), .B1(ram[4964]), .B2(n1346), 
        .ZN(n9205) );
  MOAI22 U18127 ( .A1(n27960), .A2(n1345), .B1(ram[4965]), .B2(n1346), 
        .ZN(n9206) );
  MOAI22 U18128 ( .A1(n27725), .A2(n1345), .B1(ram[4966]), .B2(n1346), 
        .ZN(n9207) );
  MOAI22 U18129 ( .A1(n27490), .A2(n1345), .B1(ram[4967]), .B2(n1346), 
        .ZN(n9208) );
  MOAI22 U18130 ( .A1(n29135), .A2(n1347), .B1(ram[4968]), .B2(n1348), 
        .ZN(n9209) );
  MOAI22 U18131 ( .A1(n28900), .A2(n1347), .B1(ram[4969]), .B2(n1348), 
        .ZN(n9210) );
  MOAI22 U18132 ( .A1(n28665), .A2(n1347), .B1(ram[4970]), .B2(n1348), 
        .ZN(n9211) );
  MOAI22 U18133 ( .A1(n28430), .A2(n1347), .B1(ram[4971]), .B2(n1348), 
        .ZN(n9212) );
  MOAI22 U18134 ( .A1(n28195), .A2(n1347), .B1(ram[4972]), .B2(n1348), 
        .ZN(n9213) );
  MOAI22 U18135 ( .A1(n27960), .A2(n1347), .B1(ram[4973]), .B2(n1348), 
        .ZN(n9214) );
  MOAI22 U18136 ( .A1(n27725), .A2(n1347), .B1(ram[4974]), .B2(n1348), 
        .ZN(n9215) );
  MOAI22 U18137 ( .A1(n27490), .A2(n1347), .B1(ram[4975]), .B2(n1348), 
        .ZN(n9216) );
  MOAI22 U18138 ( .A1(n29135), .A2(n1349), .B1(ram[4976]), .B2(n1350), 
        .ZN(n9217) );
  MOAI22 U18139 ( .A1(n28900), .A2(n1349), .B1(ram[4977]), .B2(n1350), 
        .ZN(n9218) );
  MOAI22 U18140 ( .A1(n28665), .A2(n1349), .B1(ram[4978]), .B2(n1350), 
        .ZN(n9219) );
  MOAI22 U18141 ( .A1(n28430), .A2(n1349), .B1(ram[4979]), .B2(n1350), 
        .ZN(n9220) );
  MOAI22 U18142 ( .A1(n28195), .A2(n1349), .B1(ram[4980]), .B2(n1350), 
        .ZN(n9221) );
  MOAI22 U18143 ( .A1(n27960), .A2(n1349), .B1(ram[4981]), .B2(n1350), 
        .ZN(n9222) );
  MOAI22 U18144 ( .A1(n27725), .A2(n1349), .B1(ram[4982]), .B2(n1350), 
        .ZN(n9223) );
  MOAI22 U18145 ( .A1(n27490), .A2(n1349), .B1(ram[4983]), .B2(n1350), 
        .ZN(n9224) );
  MOAI22 U18146 ( .A1(n29135), .A2(n1351), .B1(ram[4984]), .B2(n1352), 
        .ZN(n9225) );
  MOAI22 U18147 ( .A1(n28900), .A2(n1351), .B1(ram[4985]), .B2(n1352), 
        .ZN(n9226) );
  MOAI22 U18148 ( .A1(n28665), .A2(n1351), .B1(ram[4986]), .B2(n1352), 
        .ZN(n9227) );
  MOAI22 U18149 ( .A1(n28430), .A2(n1351), .B1(ram[4987]), .B2(n1352), 
        .ZN(n9228) );
  MOAI22 U18150 ( .A1(n28195), .A2(n1351), .B1(ram[4988]), .B2(n1352), 
        .ZN(n9229) );
  MOAI22 U18151 ( .A1(n27960), .A2(n1351), .B1(ram[4989]), .B2(n1352), 
        .ZN(n9230) );
  MOAI22 U18152 ( .A1(n27725), .A2(n1351), .B1(ram[4990]), .B2(n1352), 
        .ZN(n9231) );
  MOAI22 U18153 ( .A1(n27490), .A2(n1351), .B1(ram[4991]), .B2(n1352), 
        .ZN(n9232) );
  MOAI22 U18154 ( .A1(n29136), .A2(n1353), .B1(ram[4992]), .B2(n1354), 
        .ZN(n9233) );
  MOAI22 U18155 ( .A1(n28901), .A2(n1353), .B1(ram[4993]), .B2(n1354), 
        .ZN(n9234) );
  MOAI22 U18156 ( .A1(n28666), .A2(n1353), .B1(ram[4994]), .B2(n1354), 
        .ZN(n9235) );
  MOAI22 U18157 ( .A1(n28431), .A2(n1353), .B1(ram[4995]), .B2(n1354), 
        .ZN(n9236) );
  MOAI22 U18158 ( .A1(n28196), .A2(n1353), .B1(ram[4996]), .B2(n1354), 
        .ZN(n9237) );
  MOAI22 U18159 ( .A1(n27961), .A2(n1353), .B1(ram[4997]), .B2(n1354), 
        .ZN(n9238) );
  MOAI22 U18160 ( .A1(n27726), .A2(n1353), .B1(ram[4998]), .B2(n1354), 
        .ZN(n9239) );
  MOAI22 U18161 ( .A1(n27491), .A2(n1353), .B1(ram[4999]), .B2(n1354), 
        .ZN(n9240) );
  MOAI22 U18162 ( .A1(n29136), .A2(n1355), .B1(ram[5000]), .B2(n1356), 
        .ZN(n9241) );
  MOAI22 U18163 ( .A1(n28901), .A2(n1355), .B1(ram[5001]), .B2(n1356), 
        .ZN(n9242) );
  MOAI22 U18164 ( .A1(n28666), .A2(n1355), .B1(ram[5002]), .B2(n1356), 
        .ZN(n9243) );
  MOAI22 U18165 ( .A1(n28431), .A2(n1355), .B1(ram[5003]), .B2(n1356), 
        .ZN(n9244) );
  MOAI22 U18166 ( .A1(n28196), .A2(n1355), .B1(ram[5004]), .B2(n1356), 
        .ZN(n9245) );
  MOAI22 U18167 ( .A1(n27961), .A2(n1355), .B1(ram[5005]), .B2(n1356), 
        .ZN(n9246) );
  MOAI22 U18168 ( .A1(n27726), .A2(n1355), .B1(ram[5006]), .B2(n1356), 
        .ZN(n9247) );
  MOAI22 U18169 ( .A1(n27491), .A2(n1355), .B1(ram[5007]), .B2(n1356), 
        .ZN(n9248) );
  MOAI22 U18170 ( .A1(n29136), .A2(n1357), .B1(ram[5008]), .B2(n1358), 
        .ZN(n9249) );
  MOAI22 U18171 ( .A1(n28901), .A2(n1357), .B1(ram[5009]), .B2(n1358), 
        .ZN(n9250) );
  MOAI22 U18172 ( .A1(n28666), .A2(n1357), .B1(ram[5010]), .B2(n1358), 
        .ZN(n9251) );
  MOAI22 U18173 ( .A1(n28431), .A2(n1357), .B1(ram[5011]), .B2(n1358), 
        .ZN(n9252) );
  MOAI22 U18174 ( .A1(n28196), .A2(n1357), .B1(ram[5012]), .B2(n1358), 
        .ZN(n9253) );
  MOAI22 U18175 ( .A1(n27961), .A2(n1357), .B1(ram[5013]), .B2(n1358), 
        .ZN(n9254) );
  MOAI22 U18176 ( .A1(n27726), .A2(n1357), .B1(ram[5014]), .B2(n1358), 
        .ZN(n9255) );
  MOAI22 U18177 ( .A1(n27491), .A2(n1357), .B1(ram[5015]), .B2(n1358), 
        .ZN(n9256) );
  MOAI22 U18178 ( .A1(n29136), .A2(n1359), .B1(ram[5016]), .B2(n1360), 
        .ZN(n9257) );
  MOAI22 U18179 ( .A1(n28901), .A2(n1359), .B1(ram[5017]), .B2(n1360), 
        .ZN(n9258) );
  MOAI22 U18180 ( .A1(n28666), .A2(n1359), .B1(ram[5018]), .B2(n1360), 
        .ZN(n9259) );
  MOAI22 U18181 ( .A1(n28431), .A2(n1359), .B1(ram[5019]), .B2(n1360), 
        .ZN(n9260) );
  MOAI22 U18182 ( .A1(n28196), .A2(n1359), .B1(ram[5020]), .B2(n1360), 
        .ZN(n9261) );
  MOAI22 U18183 ( .A1(n27961), .A2(n1359), .B1(ram[5021]), .B2(n1360), 
        .ZN(n9262) );
  MOAI22 U18184 ( .A1(n27726), .A2(n1359), .B1(ram[5022]), .B2(n1360), 
        .ZN(n9263) );
  MOAI22 U18185 ( .A1(n27491), .A2(n1359), .B1(ram[5023]), .B2(n1360), 
        .ZN(n9264) );
  MOAI22 U18186 ( .A1(n29136), .A2(n1361), .B1(ram[5024]), .B2(n1362), 
        .ZN(n9265) );
  MOAI22 U18187 ( .A1(n28901), .A2(n1361), .B1(ram[5025]), .B2(n1362), 
        .ZN(n9266) );
  MOAI22 U18188 ( .A1(n28666), .A2(n1361), .B1(ram[5026]), .B2(n1362), 
        .ZN(n9267) );
  MOAI22 U18189 ( .A1(n28431), .A2(n1361), .B1(ram[5027]), .B2(n1362), 
        .ZN(n9268) );
  MOAI22 U18190 ( .A1(n28196), .A2(n1361), .B1(ram[5028]), .B2(n1362), 
        .ZN(n9269) );
  MOAI22 U18191 ( .A1(n27961), .A2(n1361), .B1(ram[5029]), .B2(n1362), 
        .ZN(n9270) );
  MOAI22 U18192 ( .A1(n27726), .A2(n1361), .B1(ram[5030]), .B2(n1362), 
        .ZN(n9271) );
  MOAI22 U18193 ( .A1(n27491), .A2(n1361), .B1(ram[5031]), .B2(n1362), 
        .ZN(n9272) );
  MOAI22 U18194 ( .A1(n29136), .A2(n1363), .B1(ram[5032]), .B2(n1364), 
        .ZN(n9273) );
  MOAI22 U18195 ( .A1(n28901), .A2(n1363), .B1(ram[5033]), .B2(n1364), 
        .ZN(n9274) );
  MOAI22 U18196 ( .A1(n28666), .A2(n1363), .B1(ram[5034]), .B2(n1364), 
        .ZN(n9275) );
  MOAI22 U18197 ( .A1(n28431), .A2(n1363), .B1(ram[5035]), .B2(n1364), 
        .ZN(n9276) );
  MOAI22 U18198 ( .A1(n28196), .A2(n1363), .B1(ram[5036]), .B2(n1364), 
        .ZN(n9277) );
  MOAI22 U18199 ( .A1(n27961), .A2(n1363), .B1(ram[5037]), .B2(n1364), 
        .ZN(n9278) );
  MOAI22 U18200 ( .A1(n27726), .A2(n1363), .B1(ram[5038]), .B2(n1364), 
        .ZN(n9279) );
  MOAI22 U18201 ( .A1(n27491), .A2(n1363), .B1(ram[5039]), .B2(n1364), 
        .ZN(n9280) );
  MOAI22 U18202 ( .A1(n29136), .A2(n1365), .B1(ram[5040]), .B2(n1366), 
        .ZN(n9281) );
  MOAI22 U18203 ( .A1(n28901), .A2(n1365), .B1(ram[5041]), .B2(n1366), 
        .ZN(n9282) );
  MOAI22 U18204 ( .A1(n28666), .A2(n1365), .B1(ram[5042]), .B2(n1366), 
        .ZN(n9283) );
  MOAI22 U18205 ( .A1(n28431), .A2(n1365), .B1(ram[5043]), .B2(n1366), 
        .ZN(n9284) );
  MOAI22 U18206 ( .A1(n28196), .A2(n1365), .B1(ram[5044]), .B2(n1366), 
        .ZN(n9285) );
  MOAI22 U18207 ( .A1(n27961), .A2(n1365), .B1(ram[5045]), .B2(n1366), 
        .ZN(n9286) );
  MOAI22 U18208 ( .A1(n27726), .A2(n1365), .B1(ram[5046]), .B2(n1366), 
        .ZN(n9287) );
  MOAI22 U18209 ( .A1(n27491), .A2(n1365), .B1(ram[5047]), .B2(n1366), 
        .ZN(n9288) );
  MOAI22 U18210 ( .A1(n29136), .A2(n1367), .B1(ram[5048]), .B2(n1368), 
        .ZN(n9289) );
  MOAI22 U18211 ( .A1(n28901), .A2(n1367), .B1(ram[5049]), .B2(n1368), 
        .ZN(n9290) );
  MOAI22 U18212 ( .A1(n28666), .A2(n1367), .B1(ram[5050]), .B2(n1368), 
        .ZN(n9291) );
  MOAI22 U18213 ( .A1(n28431), .A2(n1367), .B1(ram[5051]), .B2(n1368), 
        .ZN(n9292) );
  MOAI22 U18214 ( .A1(n28196), .A2(n1367), .B1(ram[5052]), .B2(n1368), 
        .ZN(n9293) );
  MOAI22 U18215 ( .A1(n27961), .A2(n1367), .B1(ram[5053]), .B2(n1368), 
        .ZN(n9294) );
  MOAI22 U18216 ( .A1(n27726), .A2(n1367), .B1(ram[5054]), .B2(n1368), 
        .ZN(n9295) );
  MOAI22 U18217 ( .A1(n27491), .A2(n1367), .B1(ram[5055]), .B2(n1368), 
        .ZN(n9296) );
  MOAI22 U18218 ( .A1(n29136), .A2(n1369), .B1(ram[5056]), .B2(n1370), 
        .ZN(n9297) );
  MOAI22 U18219 ( .A1(n28901), .A2(n1369), .B1(ram[5057]), .B2(n1370), 
        .ZN(n9298) );
  MOAI22 U18220 ( .A1(n28666), .A2(n1369), .B1(ram[5058]), .B2(n1370), 
        .ZN(n9299) );
  MOAI22 U18221 ( .A1(n28431), .A2(n1369), .B1(ram[5059]), .B2(n1370), 
        .ZN(n9300) );
  MOAI22 U18222 ( .A1(n28196), .A2(n1369), .B1(ram[5060]), .B2(n1370), 
        .ZN(n9301) );
  MOAI22 U18223 ( .A1(n27961), .A2(n1369), .B1(ram[5061]), .B2(n1370), 
        .ZN(n9302) );
  MOAI22 U18224 ( .A1(n27726), .A2(n1369), .B1(ram[5062]), .B2(n1370), 
        .ZN(n9303) );
  MOAI22 U18225 ( .A1(n27491), .A2(n1369), .B1(ram[5063]), .B2(n1370), 
        .ZN(n9304) );
  MOAI22 U18226 ( .A1(n29136), .A2(n1371), .B1(ram[5064]), .B2(n1372), 
        .ZN(n9305) );
  MOAI22 U18227 ( .A1(n28901), .A2(n1371), .B1(ram[5065]), .B2(n1372), 
        .ZN(n9306) );
  MOAI22 U18228 ( .A1(n28666), .A2(n1371), .B1(ram[5066]), .B2(n1372), 
        .ZN(n9307) );
  MOAI22 U18229 ( .A1(n28431), .A2(n1371), .B1(ram[5067]), .B2(n1372), 
        .ZN(n9308) );
  MOAI22 U18230 ( .A1(n28196), .A2(n1371), .B1(ram[5068]), .B2(n1372), 
        .ZN(n9309) );
  MOAI22 U18231 ( .A1(n27961), .A2(n1371), .B1(ram[5069]), .B2(n1372), 
        .ZN(n9310) );
  MOAI22 U18232 ( .A1(n27726), .A2(n1371), .B1(ram[5070]), .B2(n1372), 
        .ZN(n9311) );
  MOAI22 U18233 ( .A1(n27491), .A2(n1371), .B1(ram[5071]), .B2(n1372), 
        .ZN(n9312) );
  MOAI22 U18234 ( .A1(n29136), .A2(n1373), .B1(ram[5072]), .B2(n1374), 
        .ZN(n9313) );
  MOAI22 U18235 ( .A1(n28901), .A2(n1373), .B1(ram[5073]), .B2(n1374), 
        .ZN(n9314) );
  MOAI22 U18236 ( .A1(n28666), .A2(n1373), .B1(ram[5074]), .B2(n1374), 
        .ZN(n9315) );
  MOAI22 U18237 ( .A1(n28431), .A2(n1373), .B1(ram[5075]), .B2(n1374), 
        .ZN(n9316) );
  MOAI22 U18238 ( .A1(n28196), .A2(n1373), .B1(ram[5076]), .B2(n1374), 
        .ZN(n9317) );
  MOAI22 U18239 ( .A1(n27961), .A2(n1373), .B1(ram[5077]), .B2(n1374), 
        .ZN(n9318) );
  MOAI22 U18240 ( .A1(n27726), .A2(n1373), .B1(ram[5078]), .B2(n1374), 
        .ZN(n9319) );
  MOAI22 U18241 ( .A1(n27491), .A2(n1373), .B1(ram[5079]), .B2(n1374), 
        .ZN(n9320) );
  MOAI22 U18242 ( .A1(n29136), .A2(n1375), .B1(ram[5080]), .B2(n1376), 
        .ZN(n9321) );
  MOAI22 U18243 ( .A1(n28901), .A2(n1375), .B1(ram[5081]), .B2(n1376), 
        .ZN(n9322) );
  MOAI22 U18244 ( .A1(n28666), .A2(n1375), .B1(ram[5082]), .B2(n1376), 
        .ZN(n9323) );
  MOAI22 U18245 ( .A1(n28431), .A2(n1375), .B1(ram[5083]), .B2(n1376), 
        .ZN(n9324) );
  MOAI22 U18246 ( .A1(n28196), .A2(n1375), .B1(ram[5084]), .B2(n1376), 
        .ZN(n9325) );
  MOAI22 U18247 ( .A1(n27961), .A2(n1375), .B1(ram[5085]), .B2(n1376), 
        .ZN(n9326) );
  MOAI22 U18248 ( .A1(n27726), .A2(n1375), .B1(ram[5086]), .B2(n1376), 
        .ZN(n9327) );
  MOAI22 U18249 ( .A1(n27491), .A2(n1375), .B1(ram[5087]), .B2(n1376), 
        .ZN(n9328) );
  MOAI22 U18250 ( .A1(n29136), .A2(n1377), .B1(ram[5088]), .B2(n1378), 
        .ZN(n9329) );
  MOAI22 U18251 ( .A1(n28901), .A2(n1377), .B1(ram[5089]), .B2(n1378), 
        .ZN(n9330) );
  MOAI22 U18252 ( .A1(n28666), .A2(n1377), .B1(ram[5090]), .B2(n1378), 
        .ZN(n9331) );
  MOAI22 U18253 ( .A1(n28431), .A2(n1377), .B1(ram[5091]), .B2(n1378), 
        .ZN(n9332) );
  MOAI22 U18254 ( .A1(n28196), .A2(n1377), .B1(ram[5092]), .B2(n1378), 
        .ZN(n9333) );
  MOAI22 U18255 ( .A1(n27961), .A2(n1377), .B1(ram[5093]), .B2(n1378), 
        .ZN(n9334) );
  MOAI22 U18256 ( .A1(n27726), .A2(n1377), .B1(ram[5094]), .B2(n1378), 
        .ZN(n9335) );
  MOAI22 U18257 ( .A1(n27491), .A2(n1377), .B1(ram[5095]), .B2(n1378), 
        .ZN(n9336) );
  MOAI22 U18258 ( .A1(n29137), .A2(n1379), .B1(ram[5096]), .B2(n1380), 
        .ZN(n9337) );
  MOAI22 U18259 ( .A1(n28902), .A2(n1379), .B1(ram[5097]), .B2(n1380), 
        .ZN(n9338) );
  MOAI22 U18260 ( .A1(n28667), .A2(n1379), .B1(ram[5098]), .B2(n1380), 
        .ZN(n9339) );
  MOAI22 U18261 ( .A1(n28432), .A2(n1379), .B1(ram[5099]), .B2(n1380), 
        .ZN(n9340) );
  MOAI22 U18262 ( .A1(n28197), .A2(n1379), .B1(ram[5100]), .B2(n1380), 
        .ZN(n9341) );
  MOAI22 U18263 ( .A1(n27962), .A2(n1379), .B1(ram[5101]), .B2(n1380), 
        .ZN(n9342) );
  MOAI22 U18264 ( .A1(n27727), .A2(n1379), .B1(ram[5102]), .B2(n1380), 
        .ZN(n9343) );
  MOAI22 U18265 ( .A1(n27492), .A2(n1379), .B1(ram[5103]), .B2(n1380), 
        .ZN(n9344) );
  MOAI22 U18266 ( .A1(n29137), .A2(n1381), .B1(ram[5104]), .B2(n1382), 
        .ZN(n9345) );
  MOAI22 U18267 ( .A1(n28902), .A2(n1381), .B1(ram[5105]), .B2(n1382), 
        .ZN(n9346) );
  MOAI22 U18268 ( .A1(n28667), .A2(n1381), .B1(ram[5106]), .B2(n1382), 
        .ZN(n9347) );
  MOAI22 U18269 ( .A1(n28432), .A2(n1381), .B1(ram[5107]), .B2(n1382), 
        .ZN(n9348) );
  MOAI22 U18270 ( .A1(n28197), .A2(n1381), .B1(ram[5108]), .B2(n1382), 
        .ZN(n9349) );
  MOAI22 U18271 ( .A1(n27962), .A2(n1381), .B1(ram[5109]), .B2(n1382), 
        .ZN(n9350) );
  MOAI22 U18272 ( .A1(n27727), .A2(n1381), .B1(ram[5110]), .B2(n1382), 
        .ZN(n9351) );
  MOAI22 U18273 ( .A1(n27492), .A2(n1381), .B1(ram[5111]), .B2(n1382), 
        .ZN(n9352) );
  MOAI22 U18274 ( .A1(n29137), .A2(n1383), .B1(ram[5112]), .B2(n1384), 
        .ZN(n9353) );
  MOAI22 U18275 ( .A1(n28902), .A2(n1383), .B1(ram[5113]), .B2(n1384), 
        .ZN(n9354) );
  MOAI22 U18276 ( .A1(n28667), .A2(n1383), .B1(ram[5114]), .B2(n1384), 
        .ZN(n9355) );
  MOAI22 U18277 ( .A1(n28432), .A2(n1383), .B1(ram[5115]), .B2(n1384), 
        .ZN(n9356) );
  MOAI22 U18278 ( .A1(n28197), .A2(n1383), .B1(ram[5116]), .B2(n1384), 
        .ZN(n9357) );
  MOAI22 U18279 ( .A1(n27962), .A2(n1383), .B1(ram[5117]), .B2(n1384), 
        .ZN(n9358) );
  MOAI22 U18280 ( .A1(n27727), .A2(n1383), .B1(ram[5118]), .B2(n1384), 
        .ZN(n9359) );
  MOAI22 U18281 ( .A1(n27492), .A2(n1383), .B1(ram[5119]), .B2(n1384), 
        .ZN(n9360) );
  MOAI22 U18282 ( .A1(n29137), .A2(n1385), .B1(ram[5120]), .B2(n1386), 
        .ZN(n9361) );
  MOAI22 U18283 ( .A1(n28902), .A2(n1385), .B1(ram[5121]), .B2(n1386), 
        .ZN(n9362) );
  MOAI22 U18284 ( .A1(n28667), .A2(n1385), .B1(ram[5122]), .B2(n1386), 
        .ZN(n9363) );
  MOAI22 U18285 ( .A1(n28432), .A2(n1385), .B1(ram[5123]), .B2(n1386), 
        .ZN(n9364) );
  MOAI22 U18286 ( .A1(n28197), .A2(n1385), .B1(ram[5124]), .B2(n1386), 
        .ZN(n9365) );
  MOAI22 U18287 ( .A1(n27962), .A2(n1385), .B1(ram[5125]), .B2(n1386), 
        .ZN(n9366) );
  MOAI22 U18288 ( .A1(n27727), .A2(n1385), .B1(ram[5126]), .B2(n1386), 
        .ZN(n9367) );
  MOAI22 U18289 ( .A1(n27492), .A2(n1385), .B1(ram[5127]), .B2(n1386), 
        .ZN(n9368) );
  MOAI22 U18290 ( .A1(n29137), .A2(n1388), .B1(ram[5128]), .B2(n1389), 
        .ZN(n9369) );
  MOAI22 U18291 ( .A1(n28902), .A2(n1388), .B1(ram[5129]), .B2(n1389), 
        .ZN(n9370) );
  MOAI22 U18292 ( .A1(n28667), .A2(n1388), .B1(ram[5130]), .B2(n1389), 
        .ZN(n9371) );
  MOAI22 U18293 ( .A1(n28432), .A2(n1388), .B1(ram[5131]), .B2(n1389), 
        .ZN(n9372) );
  MOAI22 U18294 ( .A1(n28197), .A2(n1388), .B1(ram[5132]), .B2(n1389), 
        .ZN(n9373) );
  MOAI22 U18295 ( .A1(n27962), .A2(n1388), .B1(ram[5133]), .B2(n1389), 
        .ZN(n9374) );
  MOAI22 U18296 ( .A1(n27727), .A2(n1388), .B1(ram[5134]), .B2(n1389), 
        .ZN(n9375) );
  MOAI22 U18297 ( .A1(n27492), .A2(n1388), .B1(ram[5135]), .B2(n1389), 
        .ZN(n9376) );
  MOAI22 U18298 ( .A1(n29137), .A2(n1390), .B1(ram[5136]), .B2(n1391), 
        .ZN(n9377) );
  MOAI22 U18299 ( .A1(n28902), .A2(n1390), .B1(ram[5137]), .B2(n1391), 
        .ZN(n9378) );
  MOAI22 U18300 ( .A1(n28667), .A2(n1390), .B1(ram[5138]), .B2(n1391), 
        .ZN(n9379) );
  MOAI22 U18301 ( .A1(n28432), .A2(n1390), .B1(ram[5139]), .B2(n1391), 
        .ZN(n9380) );
  MOAI22 U18302 ( .A1(n28197), .A2(n1390), .B1(ram[5140]), .B2(n1391), 
        .ZN(n9381) );
  MOAI22 U18303 ( .A1(n27962), .A2(n1390), .B1(ram[5141]), .B2(n1391), 
        .ZN(n9382) );
  MOAI22 U18304 ( .A1(n27727), .A2(n1390), .B1(ram[5142]), .B2(n1391), 
        .ZN(n9383) );
  MOAI22 U18305 ( .A1(n27492), .A2(n1390), .B1(ram[5143]), .B2(n1391), 
        .ZN(n9384) );
  MOAI22 U18306 ( .A1(n29137), .A2(n1392), .B1(ram[5144]), .B2(n1393), 
        .ZN(n9385) );
  MOAI22 U18307 ( .A1(n28902), .A2(n1392), .B1(ram[5145]), .B2(n1393), 
        .ZN(n9386) );
  MOAI22 U18308 ( .A1(n28667), .A2(n1392), .B1(ram[5146]), .B2(n1393), 
        .ZN(n9387) );
  MOAI22 U18309 ( .A1(n28432), .A2(n1392), .B1(ram[5147]), .B2(n1393), 
        .ZN(n9388) );
  MOAI22 U18310 ( .A1(n28197), .A2(n1392), .B1(ram[5148]), .B2(n1393), 
        .ZN(n9389) );
  MOAI22 U18311 ( .A1(n27962), .A2(n1392), .B1(ram[5149]), .B2(n1393), 
        .ZN(n9390) );
  MOAI22 U18312 ( .A1(n27727), .A2(n1392), .B1(ram[5150]), .B2(n1393), 
        .ZN(n9391) );
  MOAI22 U18313 ( .A1(n27492), .A2(n1392), .B1(ram[5151]), .B2(n1393), 
        .ZN(n9392) );
  MOAI22 U18314 ( .A1(n29137), .A2(n1394), .B1(ram[5152]), .B2(n1395), 
        .ZN(n9393) );
  MOAI22 U18315 ( .A1(n28902), .A2(n1394), .B1(ram[5153]), .B2(n1395), 
        .ZN(n9394) );
  MOAI22 U18316 ( .A1(n28667), .A2(n1394), .B1(ram[5154]), .B2(n1395), 
        .ZN(n9395) );
  MOAI22 U18317 ( .A1(n28432), .A2(n1394), .B1(ram[5155]), .B2(n1395), 
        .ZN(n9396) );
  MOAI22 U18318 ( .A1(n28197), .A2(n1394), .B1(ram[5156]), .B2(n1395), 
        .ZN(n9397) );
  MOAI22 U18319 ( .A1(n27962), .A2(n1394), .B1(ram[5157]), .B2(n1395), 
        .ZN(n9398) );
  MOAI22 U18320 ( .A1(n27727), .A2(n1394), .B1(ram[5158]), .B2(n1395), 
        .ZN(n9399) );
  MOAI22 U18321 ( .A1(n27492), .A2(n1394), .B1(ram[5159]), .B2(n1395), 
        .ZN(n9400) );
  MOAI22 U18322 ( .A1(n29137), .A2(n1396), .B1(ram[5160]), .B2(n1397), 
        .ZN(n9401) );
  MOAI22 U18323 ( .A1(n28902), .A2(n1396), .B1(ram[5161]), .B2(n1397), 
        .ZN(n9402) );
  MOAI22 U18324 ( .A1(n28667), .A2(n1396), .B1(ram[5162]), .B2(n1397), 
        .ZN(n9403) );
  MOAI22 U18325 ( .A1(n28432), .A2(n1396), .B1(ram[5163]), .B2(n1397), 
        .ZN(n9404) );
  MOAI22 U18326 ( .A1(n28197), .A2(n1396), .B1(ram[5164]), .B2(n1397), 
        .ZN(n9405) );
  MOAI22 U18327 ( .A1(n27962), .A2(n1396), .B1(ram[5165]), .B2(n1397), 
        .ZN(n9406) );
  MOAI22 U18328 ( .A1(n27727), .A2(n1396), .B1(ram[5166]), .B2(n1397), 
        .ZN(n9407) );
  MOAI22 U18329 ( .A1(n27492), .A2(n1396), .B1(ram[5167]), .B2(n1397), 
        .ZN(n9408) );
  MOAI22 U18330 ( .A1(n29137), .A2(n1398), .B1(ram[5168]), .B2(n1399), 
        .ZN(n9409) );
  MOAI22 U18331 ( .A1(n28902), .A2(n1398), .B1(ram[5169]), .B2(n1399), 
        .ZN(n9410) );
  MOAI22 U18332 ( .A1(n28667), .A2(n1398), .B1(ram[5170]), .B2(n1399), 
        .ZN(n9411) );
  MOAI22 U18333 ( .A1(n28432), .A2(n1398), .B1(ram[5171]), .B2(n1399), 
        .ZN(n9412) );
  MOAI22 U18334 ( .A1(n28197), .A2(n1398), .B1(ram[5172]), .B2(n1399), 
        .ZN(n9413) );
  MOAI22 U18335 ( .A1(n27962), .A2(n1398), .B1(ram[5173]), .B2(n1399), 
        .ZN(n9414) );
  MOAI22 U18336 ( .A1(n27727), .A2(n1398), .B1(ram[5174]), .B2(n1399), 
        .ZN(n9415) );
  MOAI22 U18337 ( .A1(n27492), .A2(n1398), .B1(ram[5175]), .B2(n1399), 
        .ZN(n9416) );
  MOAI22 U18338 ( .A1(n29137), .A2(n1400), .B1(ram[5176]), .B2(n1401), 
        .ZN(n9417) );
  MOAI22 U18339 ( .A1(n28902), .A2(n1400), .B1(ram[5177]), .B2(n1401), 
        .ZN(n9418) );
  MOAI22 U18340 ( .A1(n28667), .A2(n1400), .B1(ram[5178]), .B2(n1401), 
        .ZN(n9419) );
  MOAI22 U18341 ( .A1(n28432), .A2(n1400), .B1(ram[5179]), .B2(n1401), 
        .ZN(n9420) );
  MOAI22 U18342 ( .A1(n28197), .A2(n1400), .B1(ram[5180]), .B2(n1401), 
        .ZN(n9421) );
  MOAI22 U18343 ( .A1(n27962), .A2(n1400), .B1(ram[5181]), .B2(n1401), 
        .ZN(n9422) );
  MOAI22 U18344 ( .A1(n27727), .A2(n1400), .B1(ram[5182]), .B2(n1401), 
        .ZN(n9423) );
  MOAI22 U18345 ( .A1(n27492), .A2(n1400), .B1(ram[5183]), .B2(n1401), 
        .ZN(n9424) );
  MOAI22 U18346 ( .A1(n29137), .A2(n1402), .B1(ram[5184]), .B2(n1403), 
        .ZN(n9425) );
  MOAI22 U18347 ( .A1(n28902), .A2(n1402), .B1(ram[5185]), .B2(n1403), 
        .ZN(n9426) );
  MOAI22 U18348 ( .A1(n28667), .A2(n1402), .B1(ram[5186]), .B2(n1403), 
        .ZN(n9427) );
  MOAI22 U18349 ( .A1(n28432), .A2(n1402), .B1(ram[5187]), .B2(n1403), 
        .ZN(n9428) );
  MOAI22 U18350 ( .A1(n28197), .A2(n1402), .B1(ram[5188]), .B2(n1403), 
        .ZN(n9429) );
  MOAI22 U18351 ( .A1(n27962), .A2(n1402), .B1(ram[5189]), .B2(n1403), 
        .ZN(n9430) );
  MOAI22 U18352 ( .A1(n27727), .A2(n1402), .B1(ram[5190]), .B2(n1403), 
        .ZN(n9431) );
  MOAI22 U18353 ( .A1(n27492), .A2(n1402), .B1(ram[5191]), .B2(n1403), 
        .ZN(n9432) );
  MOAI22 U18354 ( .A1(n29137), .A2(n1404), .B1(ram[5192]), .B2(n1405), 
        .ZN(n9433) );
  MOAI22 U18355 ( .A1(n28902), .A2(n1404), .B1(ram[5193]), .B2(n1405), 
        .ZN(n9434) );
  MOAI22 U18356 ( .A1(n28667), .A2(n1404), .B1(ram[5194]), .B2(n1405), 
        .ZN(n9435) );
  MOAI22 U18357 ( .A1(n28432), .A2(n1404), .B1(ram[5195]), .B2(n1405), 
        .ZN(n9436) );
  MOAI22 U18358 ( .A1(n28197), .A2(n1404), .B1(ram[5196]), .B2(n1405), 
        .ZN(n9437) );
  MOAI22 U18359 ( .A1(n27962), .A2(n1404), .B1(ram[5197]), .B2(n1405), 
        .ZN(n9438) );
  MOAI22 U18360 ( .A1(n27727), .A2(n1404), .B1(ram[5198]), .B2(n1405), 
        .ZN(n9439) );
  MOAI22 U18361 ( .A1(n27492), .A2(n1404), .B1(ram[5199]), .B2(n1405), 
        .ZN(n9440) );
  MOAI22 U18362 ( .A1(n29138), .A2(n1406), .B1(ram[5200]), .B2(n1407), 
        .ZN(n9441) );
  MOAI22 U18363 ( .A1(n28903), .A2(n1406), .B1(ram[5201]), .B2(n1407), 
        .ZN(n9442) );
  MOAI22 U18364 ( .A1(n28668), .A2(n1406), .B1(ram[5202]), .B2(n1407), 
        .ZN(n9443) );
  MOAI22 U18365 ( .A1(n28433), .A2(n1406), .B1(ram[5203]), .B2(n1407), 
        .ZN(n9444) );
  MOAI22 U18366 ( .A1(n28198), .A2(n1406), .B1(ram[5204]), .B2(n1407), 
        .ZN(n9445) );
  MOAI22 U18367 ( .A1(n27963), .A2(n1406), .B1(ram[5205]), .B2(n1407), 
        .ZN(n9446) );
  MOAI22 U18368 ( .A1(n27728), .A2(n1406), .B1(ram[5206]), .B2(n1407), 
        .ZN(n9447) );
  MOAI22 U18369 ( .A1(n27493), .A2(n1406), .B1(ram[5207]), .B2(n1407), 
        .ZN(n9448) );
  MOAI22 U18370 ( .A1(n29138), .A2(n1408), .B1(ram[5208]), .B2(n1409), 
        .ZN(n9449) );
  MOAI22 U18371 ( .A1(n28903), .A2(n1408), .B1(ram[5209]), .B2(n1409), 
        .ZN(n9450) );
  MOAI22 U18372 ( .A1(n28668), .A2(n1408), .B1(ram[5210]), .B2(n1409), 
        .ZN(n9451) );
  MOAI22 U18373 ( .A1(n28433), .A2(n1408), .B1(ram[5211]), .B2(n1409), 
        .ZN(n9452) );
  MOAI22 U18374 ( .A1(n28198), .A2(n1408), .B1(ram[5212]), .B2(n1409), 
        .ZN(n9453) );
  MOAI22 U18375 ( .A1(n27963), .A2(n1408), .B1(ram[5213]), .B2(n1409), 
        .ZN(n9454) );
  MOAI22 U18376 ( .A1(n27728), .A2(n1408), .B1(ram[5214]), .B2(n1409), 
        .ZN(n9455) );
  MOAI22 U18377 ( .A1(n27493), .A2(n1408), .B1(ram[5215]), .B2(n1409), 
        .ZN(n9456) );
  MOAI22 U18378 ( .A1(n29138), .A2(n1410), .B1(ram[5216]), .B2(n1411), 
        .ZN(n9457) );
  MOAI22 U18379 ( .A1(n28903), .A2(n1410), .B1(ram[5217]), .B2(n1411), 
        .ZN(n9458) );
  MOAI22 U18380 ( .A1(n28668), .A2(n1410), .B1(ram[5218]), .B2(n1411), 
        .ZN(n9459) );
  MOAI22 U18381 ( .A1(n28433), .A2(n1410), .B1(ram[5219]), .B2(n1411), 
        .ZN(n9460) );
  MOAI22 U18382 ( .A1(n28198), .A2(n1410), .B1(ram[5220]), .B2(n1411), 
        .ZN(n9461) );
  MOAI22 U18383 ( .A1(n27963), .A2(n1410), .B1(ram[5221]), .B2(n1411), 
        .ZN(n9462) );
  MOAI22 U18384 ( .A1(n27728), .A2(n1410), .B1(ram[5222]), .B2(n1411), 
        .ZN(n9463) );
  MOAI22 U18385 ( .A1(n27493), .A2(n1410), .B1(ram[5223]), .B2(n1411), 
        .ZN(n9464) );
  MOAI22 U18386 ( .A1(n29138), .A2(n1412), .B1(ram[5224]), .B2(n1413), 
        .ZN(n9465) );
  MOAI22 U18387 ( .A1(n28903), .A2(n1412), .B1(ram[5225]), .B2(n1413), 
        .ZN(n9466) );
  MOAI22 U18388 ( .A1(n28668), .A2(n1412), .B1(ram[5226]), .B2(n1413), 
        .ZN(n9467) );
  MOAI22 U18389 ( .A1(n28433), .A2(n1412), .B1(ram[5227]), .B2(n1413), 
        .ZN(n9468) );
  MOAI22 U18390 ( .A1(n28198), .A2(n1412), .B1(ram[5228]), .B2(n1413), 
        .ZN(n9469) );
  MOAI22 U18391 ( .A1(n27963), .A2(n1412), .B1(ram[5229]), .B2(n1413), 
        .ZN(n9470) );
  MOAI22 U18392 ( .A1(n27728), .A2(n1412), .B1(ram[5230]), .B2(n1413), 
        .ZN(n9471) );
  MOAI22 U18393 ( .A1(n27493), .A2(n1412), .B1(ram[5231]), .B2(n1413), 
        .ZN(n9472) );
  MOAI22 U18394 ( .A1(n29138), .A2(n1414), .B1(ram[5232]), .B2(n1415), 
        .ZN(n9473) );
  MOAI22 U18395 ( .A1(n28903), .A2(n1414), .B1(ram[5233]), .B2(n1415), 
        .ZN(n9474) );
  MOAI22 U18396 ( .A1(n28668), .A2(n1414), .B1(ram[5234]), .B2(n1415), 
        .ZN(n9475) );
  MOAI22 U18397 ( .A1(n28433), .A2(n1414), .B1(ram[5235]), .B2(n1415), 
        .ZN(n9476) );
  MOAI22 U18398 ( .A1(n28198), .A2(n1414), .B1(ram[5236]), .B2(n1415), 
        .ZN(n9477) );
  MOAI22 U18399 ( .A1(n27963), .A2(n1414), .B1(ram[5237]), .B2(n1415), 
        .ZN(n9478) );
  MOAI22 U18400 ( .A1(n27728), .A2(n1414), .B1(ram[5238]), .B2(n1415), 
        .ZN(n9479) );
  MOAI22 U18401 ( .A1(n27493), .A2(n1414), .B1(ram[5239]), .B2(n1415), 
        .ZN(n9480) );
  MOAI22 U18402 ( .A1(n29138), .A2(n1416), .B1(ram[5240]), .B2(n1417), 
        .ZN(n9481) );
  MOAI22 U18403 ( .A1(n28903), .A2(n1416), .B1(ram[5241]), .B2(n1417), 
        .ZN(n9482) );
  MOAI22 U18404 ( .A1(n28668), .A2(n1416), .B1(ram[5242]), .B2(n1417), 
        .ZN(n9483) );
  MOAI22 U18405 ( .A1(n28433), .A2(n1416), .B1(ram[5243]), .B2(n1417), 
        .ZN(n9484) );
  MOAI22 U18406 ( .A1(n28198), .A2(n1416), .B1(ram[5244]), .B2(n1417), 
        .ZN(n9485) );
  MOAI22 U18407 ( .A1(n27963), .A2(n1416), .B1(ram[5245]), .B2(n1417), 
        .ZN(n9486) );
  MOAI22 U18408 ( .A1(n27728), .A2(n1416), .B1(ram[5246]), .B2(n1417), 
        .ZN(n9487) );
  MOAI22 U18409 ( .A1(n27493), .A2(n1416), .B1(ram[5247]), .B2(n1417), 
        .ZN(n9488) );
  MOAI22 U18410 ( .A1(n29138), .A2(n1418), .B1(ram[5248]), .B2(n1419), 
        .ZN(n9489) );
  MOAI22 U18411 ( .A1(n28903), .A2(n1418), .B1(ram[5249]), .B2(n1419), 
        .ZN(n9490) );
  MOAI22 U18412 ( .A1(n28668), .A2(n1418), .B1(ram[5250]), .B2(n1419), 
        .ZN(n9491) );
  MOAI22 U18413 ( .A1(n28433), .A2(n1418), .B1(ram[5251]), .B2(n1419), 
        .ZN(n9492) );
  MOAI22 U18414 ( .A1(n28198), .A2(n1418), .B1(ram[5252]), .B2(n1419), 
        .ZN(n9493) );
  MOAI22 U18415 ( .A1(n27963), .A2(n1418), .B1(ram[5253]), .B2(n1419), 
        .ZN(n9494) );
  MOAI22 U18416 ( .A1(n27728), .A2(n1418), .B1(ram[5254]), .B2(n1419), 
        .ZN(n9495) );
  MOAI22 U18417 ( .A1(n27493), .A2(n1418), .B1(ram[5255]), .B2(n1419), 
        .ZN(n9496) );
  MOAI22 U18418 ( .A1(n29138), .A2(n1420), .B1(ram[5256]), .B2(n1421), 
        .ZN(n9497) );
  MOAI22 U18419 ( .A1(n28903), .A2(n1420), .B1(ram[5257]), .B2(n1421), 
        .ZN(n9498) );
  MOAI22 U18420 ( .A1(n28668), .A2(n1420), .B1(ram[5258]), .B2(n1421), 
        .ZN(n9499) );
  MOAI22 U18421 ( .A1(n28433), .A2(n1420), .B1(ram[5259]), .B2(n1421), 
        .ZN(n9500) );
  MOAI22 U18422 ( .A1(n28198), .A2(n1420), .B1(ram[5260]), .B2(n1421), 
        .ZN(n9501) );
  MOAI22 U18423 ( .A1(n27963), .A2(n1420), .B1(ram[5261]), .B2(n1421), 
        .ZN(n9502) );
  MOAI22 U18424 ( .A1(n27728), .A2(n1420), .B1(ram[5262]), .B2(n1421), 
        .ZN(n9503) );
  MOAI22 U18425 ( .A1(n27493), .A2(n1420), .B1(ram[5263]), .B2(n1421), 
        .ZN(n9504) );
  MOAI22 U18426 ( .A1(n29138), .A2(n1422), .B1(ram[5264]), .B2(n1423), 
        .ZN(n9505) );
  MOAI22 U18427 ( .A1(n28903), .A2(n1422), .B1(ram[5265]), .B2(n1423), 
        .ZN(n9506) );
  MOAI22 U18428 ( .A1(n28668), .A2(n1422), .B1(ram[5266]), .B2(n1423), 
        .ZN(n9507) );
  MOAI22 U18429 ( .A1(n28433), .A2(n1422), .B1(ram[5267]), .B2(n1423), 
        .ZN(n9508) );
  MOAI22 U18430 ( .A1(n28198), .A2(n1422), .B1(ram[5268]), .B2(n1423), 
        .ZN(n9509) );
  MOAI22 U18431 ( .A1(n27963), .A2(n1422), .B1(ram[5269]), .B2(n1423), 
        .ZN(n9510) );
  MOAI22 U18432 ( .A1(n27728), .A2(n1422), .B1(ram[5270]), .B2(n1423), 
        .ZN(n9511) );
  MOAI22 U18433 ( .A1(n27493), .A2(n1422), .B1(ram[5271]), .B2(n1423), 
        .ZN(n9512) );
  MOAI22 U18434 ( .A1(n29138), .A2(n1424), .B1(ram[5272]), .B2(n1425), 
        .ZN(n9513) );
  MOAI22 U18435 ( .A1(n28903), .A2(n1424), .B1(ram[5273]), .B2(n1425), 
        .ZN(n9514) );
  MOAI22 U18436 ( .A1(n28668), .A2(n1424), .B1(ram[5274]), .B2(n1425), 
        .ZN(n9515) );
  MOAI22 U18437 ( .A1(n28433), .A2(n1424), .B1(ram[5275]), .B2(n1425), 
        .ZN(n9516) );
  MOAI22 U18438 ( .A1(n28198), .A2(n1424), .B1(ram[5276]), .B2(n1425), 
        .ZN(n9517) );
  MOAI22 U18439 ( .A1(n27963), .A2(n1424), .B1(ram[5277]), .B2(n1425), 
        .ZN(n9518) );
  MOAI22 U18440 ( .A1(n27728), .A2(n1424), .B1(ram[5278]), .B2(n1425), 
        .ZN(n9519) );
  MOAI22 U18441 ( .A1(n27493), .A2(n1424), .B1(ram[5279]), .B2(n1425), 
        .ZN(n9520) );
  MOAI22 U18442 ( .A1(n29138), .A2(n1426), .B1(ram[5280]), .B2(n1427), 
        .ZN(n9521) );
  MOAI22 U18443 ( .A1(n28903), .A2(n1426), .B1(ram[5281]), .B2(n1427), 
        .ZN(n9522) );
  MOAI22 U18444 ( .A1(n28668), .A2(n1426), .B1(ram[5282]), .B2(n1427), 
        .ZN(n9523) );
  MOAI22 U18445 ( .A1(n28433), .A2(n1426), .B1(ram[5283]), .B2(n1427), 
        .ZN(n9524) );
  MOAI22 U18446 ( .A1(n28198), .A2(n1426), .B1(ram[5284]), .B2(n1427), 
        .ZN(n9525) );
  MOAI22 U18447 ( .A1(n27963), .A2(n1426), .B1(ram[5285]), .B2(n1427), 
        .ZN(n9526) );
  MOAI22 U18448 ( .A1(n27728), .A2(n1426), .B1(ram[5286]), .B2(n1427), 
        .ZN(n9527) );
  MOAI22 U18449 ( .A1(n27493), .A2(n1426), .B1(ram[5287]), .B2(n1427), 
        .ZN(n9528) );
  MOAI22 U18450 ( .A1(n29138), .A2(n1428), .B1(ram[5288]), .B2(n1429), 
        .ZN(n9529) );
  MOAI22 U18451 ( .A1(n28903), .A2(n1428), .B1(ram[5289]), .B2(n1429), 
        .ZN(n9530) );
  MOAI22 U18452 ( .A1(n28668), .A2(n1428), .B1(ram[5290]), .B2(n1429), 
        .ZN(n9531) );
  MOAI22 U18453 ( .A1(n28433), .A2(n1428), .B1(ram[5291]), .B2(n1429), 
        .ZN(n9532) );
  MOAI22 U18454 ( .A1(n28198), .A2(n1428), .B1(ram[5292]), .B2(n1429), 
        .ZN(n9533) );
  MOAI22 U18455 ( .A1(n27963), .A2(n1428), .B1(ram[5293]), .B2(n1429), 
        .ZN(n9534) );
  MOAI22 U18456 ( .A1(n27728), .A2(n1428), .B1(ram[5294]), .B2(n1429), 
        .ZN(n9535) );
  MOAI22 U18457 ( .A1(n27493), .A2(n1428), .B1(ram[5295]), .B2(n1429), 
        .ZN(n9536) );
  MOAI22 U18458 ( .A1(n29138), .A2(n1430), .B1(ram[5296]), .B2(n1431), 
        .ZN(n9537) );
  MOAI22 U18459 ( .A1(n28903), .A2(n1430), .B1(ram[5297]), .B2(n1431), 
        .ZN(n9538) );
  MOAI22 U18460 ( .A1(n28668), .A2(n1430), .B1(ram[5298]), .B2(n1431), 
        .ZN(n9539) );
  MOAI22 U18461 ( .A1(n28433), .A2(n1430), .B1(ram[5299]), .B2(n1431), 
        .ZN(n9540) );
  MOAI22 U18462 ( .A1(n28198), .A2(n1430), .B1(ram[5300]), .B2(n1431), 
        .ZN(n9541) );
  MOAI22 U18463 ( .A1(n27963), .A2(n1430), .B1(ram[5301]), .B2(n1431), 
        .ZN(n9542) );
  MOAI22 U18464 ( .A1(n27728), .A2(n1430), .B1(ram[5302]), .B2(n1431), 
        .ZN(n9543) );
  MOAI22 U18465 ( .A1(n27493), .A2(n1430), .B1(ram[5303]), .B2(n1431), 
        .ZN(n9544) );
  MOAI22 U18466 ( .A1(n29139), .A2(n1432), .B1(ram[5304]), .B2(n1433), 
        .ZN(n9545) );
  MOAI22 U18467 ( .A1(n28904), .A2(n1432), .B1(ram[5305]), .B2(n1433), 
        .ZN(n9546) );
  MOAI22 U18468 ( .A1(n28669), .A2(n1432), .B1(ram[5306]), .B2(n1433), 
        .ZN(n9547) );
  MOAI22 U18469 ( .A1(n28434), .A2(n1432), .B1(ram[5307]), .B2(n1433), 
        .ZN(n9548) );
  MOAI22 U18470 ( .A1(n28199), .A2(n1432), .B1(ram[5308]), .B2(n1433), 
        .ZN(n9549) );
  MOAI22 U18471 ( .A1(n27964), .A2(n1432), .B1(ram[5309]), .B2(n1433), 
        .ZN(n9550) );
  MOAI22 U18472 ( .A1(n27729), .A2(n1432), .B1(ram[5310]), .B2(n1433), 
        .ZN(n9551) );
  MOAI22 U18473 ( .A1(n27494), .A2(n1432), .B1(ram[5311]), .B2(n1433), 
        .ZN(n9552) );
  MOAI22 U18474 ( .A1(n29139), .A2(n1434), .B1(ram[5312]), .B2(n1435), 
        .ZN(n9553) );
  MOAI22 U18475 ( .A1(n28904), .A2(n1434), .B1(ram[5313]), .B2(n1435), 
        .ZN(n9554) );
  MOAI22 U18476 ( .A1(n28669), .A2(n1434), .B1(ram[5314]), .B2(n1435), 
        .ZN(n9555) );
  MOAI22 U18477 ( .A1(n28434), .A2(n1434), .B1(ram[5315]), .B2(n1435), 
        .ZN(n9556) );
  MOAI22 U18478 ( .A1(n28199), .A2(n1434), .B1(ram[5316]), .B2(n1435), 
        .ZN(n9557) );
  MOAI22 U18479 ( .A1(n27964), .A2(n1434), .B1(ram[5317]), .B2(n1435), 
        .ZN(n9558) );
  MOAI22 U18480 ( .A1(n27729), .A2(n1434), .B1(ram[5318]), .B2(n1435), 
        .ZN(n9559) );
  MOAI22 U18481 ( .A1(n27494), .A2(n1434), .B1(ram[5319]), .B2(n1435), 
        .ZN(n9560) );
  MOAI22 U18482 ( .A1(n29139), .A2(n1436), .B1(ram[5320]), .B2(n1437), 
        .ZN(n9561) );
  MOAI22 U18483 ( .A1(n28904), .A2(n1436), .B1(ram[5321]), .B2(n1437), 
        .ZN(n9562) );
  MOAI22 U18484 ( .A1(n28669), .A2(n1436), .B1(ram[5322]), .B2(n1437), 
        .ZN(n9563) );
  MOAI22 U18485 ( .A1(n28434), .A2(n1436), .B1(ram[5323]), .B2(n1437), 
        .ZN(n9564) );
  MOAI22 U18486 ( .A1(n28199), .A2(n1436), .B1(ram[5324]), .B2(n1437), 
        .ZN(n9565) );
  MOAI22 U18487 ( .A1(n27964), .A2(n1436), .B1(ram[5325]), .B2(n1437), 
        .ZN(n9566) );
  MOAI22 U18488 ( .A1(n27729), .A2(n1436), .B1(ram[5326]), .B2(n1437), 
        .ZN(n9567) );
  MOAI22 U18489 ( .A1(n27494), .A2(n1436), .B1(ram[5327]), .B2(n1437), 
        .ZN(n9568) );
  MOAI22 U18490 ( .A1(n29139), .A2(n1438), .B1(ram[5328]), .B2(n1439), 
        .ZN(n9569) );
  MOAI22 U18491 ( .A1(n28904), .A2(n1438), .B1(ram[5329]), .B2(n1439), 
        .ZN(n9570) );
  MOAI22 U18492 ( .A1(n28669), .A2(n1438), .B1(ram[5330]), .B2(n1439), 
        .ZN(n9571) );
  MOAI22 U18493 ( .A1(n28434), .A2(n1438), .B1(ram[5331]), .B2(n1439), 
        .ZN(n9572) );
  MOAI22 U18494 ( .A1(n28199), .A2(n1438), .B1(ram[5332]), .B2(n1439), 
        .ZN(n9573) );
  MOAI22 U18495 ( .A1(n27964), .A2(n1438), .B1(ram[5333]), .B2(n1439), 
        .ZN(n9574) );
  MOAI22 U18496 ( .A1(n27729), .A2(n1438), .B1(ram[5334]), .B2(n1439), 
        .ZN(n9575) );
  MOAI22 U18497 ( .A1(n27494), .A2(n1438), .B1(ram[5335]), .B2(n1439), 
        .ZN(n9576) );
  MOAI22 U18498 ( .A1(n29139), .A2(n1440), .B1(ram[5336]), .B2(n1441), 
        .ZN(n9577) );
  MOAI22 U18499 ( .A1(n28904), .A2(n1440), .B1(ram[5337]), .B2(n1441), 
        .ZN(n9578) );
  MOAI22 U18500 ( .A1(n28669), .A2(n1440), .B1(ram[5338]), .B2(n1441), 
        .ZN(n9579) );
  MOAI22 U18501 ( .A1(n28434), .A2(n1440), .B1(ram[5339]), .B2(n1441), 
        .ZN(n9580) );
  MOAI22 U18502 ( .A1(n28199), .A2(n1440), .B1(ram[5340]), .B2(n1441), 
        .ZN(n9581) );
  MOAI22 U18503 ( .A1(n27964), .A2(n1440), .B1(ram[5341]), .B2(n1441), 
        .ZN(n9582) );
  MOAI22 U18504 ( .A1(n27729), .A2(n1440), .B1(ram[5342]), .B2(n1441), 
        .ZN(n9583) );
  MOAI22 U18505 ( .A1(n27494), .A2(n1440), .B1(ram[5343]), .B2(n1441), 
        .ZN(n9584) );
  MOAI22 U18506 ( .A1(n29139), .A2(n1442), .B1(ram[5344]), .B2(n1443), 
        .ZN(n9585) );
  MOAI22 U18507 ( .A1(n28904), .A2(n1442), .B1(ram[5345]), .B2(n1443), 
        .ZN(n9586) );
  MOAI22 U18508 ( .A1(n28669), .A2(n1442), .B1(ram[5346]), .B2(n1443), 
        .ZN(n9587) );
  MOAI22 U18509 ( .A1(n28434), .A2(n1442), .B1(ram[5347]), .B2(n1443), 
        .ZN(n9588) );
  MOAI22 U18510 ( .A1(n28199), .A2(n1442), .B1(ram[5348]), .B2(n1443), 
        .ZN(n9589) );
  MOAI22 U18511 ( .A1(n27964), .A2(n1442), .B1(ram[5349]), .B2(n1443), 
        .ZN(n9590) );
  MOAI22 U18512 ( .A1(n27729), .A2(n1442), .B1(ram[5350]), .B2(n1443), 
        .ZN(n9591) );
  MOAI22 U18513 ( .A1(n27494), .A2(n1442), .B1(ram[5351]), .B2(n1443), 
        .ZN(n9592) );
  MOAI22 U18514 ( .A1(n29139), .A2(n1444), .B1(ram[5352]), .B2(n1445), 
        .ZN(n9593) );
  MOAI22 U18515 ( .A1(n28904), .A2(n1444), .B1(ram[5353]), .B2(n1445), 
        .ZN(n9594) );
  MOAI22 U18516 ( .A1(n28669), .A2(n1444), .B1(ram[5354]), .B2(n1445), 
        .ZN(n9595) );
  MOAI22 U18517 ( .A1(n28434), .A2(n1444), .B1(ram[5355]), .B2(n1445), 
        .ZN(n9596) );
  MOAI22 U18518 ( .A1(n28199), .A2(n1444), .B1(ram[5356]), .B2(n1445), 
        .ZN(n9597) );
  MOAI22 U18519 ( .A1(n27964), .A2(n1444), .B1(ram[5357]), .B2(n1445), 
        .ZN(n9598) );
  MOAI22 U18520 ( .A1(n27729), .A2(n1444), .B1(ram[5358]), .B2(n1445), 
        .ZN(n9599) );
  MOAI22 U18521 ( .A1(n27494), .A2(n1444), .B1(ram[5359]), .B2(n1445), 
        .ZN(n9600) );
  MOAI22 U18522 ( .A1(n29139), .A2(n1446), .B1(ram[5360]), .B2(n1447), 
        .ZN(n9601) );
  MOAI22 U18523 ( .A1(n28904), .A2(n1446), .B1(ram[5361]), .B2(n1447), 
        .ZN(n9602) );
  MOAI22 U18524 ( .A1(n28669), .A2(n1446), .B1(ram[5362]), .B2(n1447), 
        .ZN(n9603) );
  MOAI22 U18525 ( .A1(n28434), .A2(n1446), .B1(ram[5363]), .B2(n1447), 
        .ZN(n9604) );
  MOAI22 U18526 ( .A1(n28199), .A2(n1446), .B1(ram[5364]), .B2(n1447), 
        .ZN(n9605) );
  MOAI22 U18527 ( .A1(n27964), .A2(n1446), .B1(ram[5365]), .B2(n1447), 
        .ZN(n9606) );
  MOAI22 U18528 ( .A1(n27729), .A2(n1446), .B1(ram[5366]), .B2(n1447), 
        .ZN(n9607) );
  MOAI22 U18529 ( .A1(n27494), .A2(n1446), .B1(ram[5367]), .B2(n1447), 
        .ZN(n9608) );
  MOAI22 U18530 ( .A1(n29139), .A2(n1448), .B1(ram[5368]), .B2(n1449), 
        .ZN(n9609) );
  MOAI22 U18531 ( .A1(n28904), .A2(n1448), .B1(ram[5369]), .B2(n1449), 
        .ZN(n9610) );
  MOAI22 U18532 ( .A1(n28669), .A2(n1448), .B1(ram[5370]), .B2(n1449), 
        .ZN(n9611) );
  MOAI22 U18533 ( .A1(n28434), .A2(n1448), .B1(ram[5371]), .B2(n1449), 
        .ZN(n9612) );
  MOAI22 U18534 ( .A1(n28199), .A2(n1448), .B1(ram[5372]), .B2(n1449), 
        .ZN(n9613) );
  MOAI22 U18535 ( .A1(n27964), .A2(n1448), .B1(ram[5373]), .B2(n1449), 
        .ZN(n9614) );
  MOAI22 U18536 ( .A1(n27729), .A2(n1448), .B1(ram[5374]), .B2(n1449), 
        .ZN(n9615) );
  MOAI22 U18537 ( .A1(n27494), .A2(n1448), .B1(ram[5375]), .B2(n1449), 
        .ZN(n9616) );
  MOAI22 U18538 ( .A1(n29139), .A2(n1450), .B1(ram[5376]), .B2(n1451), 
        .ZN(n9617) );
  MOAI22 U18539 ( .A1(n28904), .A2(n1450), .B1(ram[5377]), .B2(n1451), 
        .ZN(n9618) );
  MOAI22 U18540 ( .A1(n28669), .A2(n1450), .B1(ram[5378]), .B2(n1451), 
        .ZN(n9619) );
  MOAI22 U18541 ( .A1(n28434), .A2(n1450), .B1(ram[5379]), .B2(n1451), 
        .ZN(n9620) );
  MOAI22 U18542 ( .A1(n28199), .A2(n1450), .B1(ram[5380]), .B2(n1451), 
        .ZN(n9621) );
  MOAI22 U18543 ( .A1(n27964), .A2(n1450), .B1(ram[5381]), .B2(n1451), 
        .ZN(n9622) );
  MOAI22 U18544 ( .A1(n27729), .A2(n1450), .B1(ram[5382]), .B2(n1451), 
        .ZN(n9623) );
  MOAI22 U18545 ( .A1(n27494), .A2(n1450), .B1(ram[5383]), .B2(n1451), 
        .ZN(n9624) );
  MOAI22 U18546 ( .A1(n29139), .A2(n1452), .B1(ram[5384]), .B2(n1453), 
        .ZN(n9625) );
  MOAI22 U18547 ( .A1(n28904), .A2(n1452), .B1(ram[5385]), .B2(n1453), 
        .ZN(n9626) );
  MOAI22 U18548 ( .A1(n28669), .A2(n1452), .B1(ram[5386]), .B2(n1453), 
        .ZN(n9627) );
  MOAI22 U18549 ( .A1(n28434), .A2(n1452), .B1(ram[5387]), .B2(n1453), 
        .ZN(n9628) );
  MOAI22 U18550 ( .A1(n28199), .A2(n1452), .B1(ram[5388]), .B2(n1453), 
        .ZN(n9629) );
  MOAI22 U18551 ( .A1(n27964), .A2(n1452), .B1(ram[5389]), .B2(n1453), 
        .ZN(n9630) );
  MOAI22 U18552 ( .A1(n27729), .A2(n1452), .B1(ram[5390]), .B2(n1453), 
        .ZN(n9631) );
  MOAI22 U18553 ( .A1(n27494), .A2(n1452), .B1(ram[5391]), .B2(n1453), 
        .ZN(n9632) );
  MOAI22 U18554 ( .A1(n29139), .A2(n1454), .B1(ram[5392]), .B2(n1455), 
        .ZN(n9633) );
  MOAI22 U18555 ( .A1(n28904), .A2(n1454), .B1(ram[5393]), .B2(n1455), 
        .ZN(n9634) );
  MOAI22 U18556 ( .A1(n28669), .A2(n1454), .B1(ram[5394]), .B2(n1455), 
        .ZN(n9635) );
  MOAI22 U18557 ( .A1(n28434), .A2(n1454), .B1(ram[5395]), .B2(n1455), 
        .ZN(n9636) );
  MOAI22 U18558 ( .A1(n28199), .A2(n1454), .B1(ram[5396]), .B2(n1455), 
        .ZN(n9637) );
  MOAI22 U18559 ( .A1(n27964), .A2(n1454), .B1(ram[5397]), .B2(n1455), 
        .ZN(n9638) );
  MOAI22 U18560 ( .A1(n27729), .A2(n1454), .B1(ram[5398]), .B2(n1455), 
        .ZN(n9639) );
  MOAI22 U18561 ( .A1(n27494), .A2(n1454), .B1(ram[5399]), .B2(n1455), 
        .ZN(n9640) );
  MOAI22 U18562 ( .A1(n29139), .A2(n1456), .B1(ram[5400]), .B2(n1457), 
        .ZN(n9641) );
  MOAI22 U18563 ( .A1(n28904), .A2(n1456), .B1(ram[5401]), .B2(n1457), 
        .ZN(n9642) );
  MOAI22 U18564 ( .A1(n28669), .A2(n1456), .B1(ram[5402]), .B2(n1457), 
        .ZN(n9643) );
  MOAI22 U18565 ( .A1(n28434), .A2(n1456), .B1(ram[5403]), .B2(n1457), 
        .ZN(n9644) );
  MOAI22 U18566 ( .A1(n28199), .A2(n1456), .B1(ram[5404]), .B2(n1457), 
        .ZN(n9645) );
  MOAI22 U18567 ( .A1(n27964), .A2(n1456), .B1(ram[5405]), .B2(n1457), 
        .ZN(n9646) );
  MOAI22 U18568 ( .A1(n27729), .A2(n1456), .B1(ram[5406]), .B2(n1457), 
        .ZN(n9647) );
  MOAI22 U18569 ( .A1(n27494), .A2(n1456), .B1(ram[5407]), .B2(n1457), 
        .ZN(n9648) );
  MOAI22 U18570 ( .A1(n29140), .A2(n1458), .B1(ram[5408]), .B2(n1459), 
        .ZN(n9649) );
  MOAI22 U18571 ( .A1(n28905), .A2(n1458), .B1(ram[5409]), .B2(n1459), 
        .ZN(n9650) );
  MOAI22 U18572 ( .A1(n28670), .A2(n1458), .B1(ram[5410]), .B2(n1459), 
        .ZN(n9651) );
  MOAI22 U18573 ( .A1(n28435), .A2(n1458), .B1(ram[5411]), .B2(n1459), 
        .ZN(n9652) );
  MOAI22 U18574 ( .A1(n28200), .A2(n1458), .B1(ram[5412]), .B2(n1459), 
        .ZN(n9653) );
  MOAI22 U18575 ( .A1(n27965), .A2(n1458), .B1(ram[5413]), .B2(n1459), 
        .ZN(n9654) );
  MOAI22 U18576 ( .A1(n27730), .A2(n1458), .B1(ram[5414]), .B2(n1459), 
        .ZN(n9655) );
  MOAI22 U18577 ( .A1(n27495), .A2(n1458), .B1(ram[5415]), .B2(n1459), 
        .ZN(n9656) );
  MOAI22 U18578 ( .A1(n29140), .A2(n1460), .B1(ram[5416]), .B2(n1461), 
        .ZN(n9657) );
  MOAI22 U18579 ( .A1(n28905), .A2(n1460), .B1(ram[5417]), .B2(n1461), 
        .ZN(n9658) );
  MOAI22 U18580 ( .A1(n28670), .A2(n1460), .B1(ram[5418]), .B2(n1461), 
        .ZN(n9659) );
  MOAI22 U18581 ( .A1(n28435), .A2(n1460), .B1(ram[5419]), .B2(n1461), 
        .ZN(n9660) );
  MOAI22 U18582 ( .A1(n28200), .A2(n1460), .B1(ram[5420]), .B2(n1461), 
        .ZN(n9661) );
  MOAI22 U18583 ( .A1(n27965), .A2(n1460), .B1(ram[5421]), .B2(n1461), 
        .ZN(n9662) );
  MOAI22 U18584 ( .A1(n27730), .A2(n1460), .B1(ram[5422]), .B2(n1461), 
        .ZN(n9663) );
  MOAI22 U18585 ( .A1(n27495), .A2(n1460), .B1(ram[5423]), .B2(n1461), 
        .ZN(n9664) );
  MOAI22 U18586 ( .A1(n29140), .A2(n1462), .B1(ram[5424]), .B2(n1463), 
        .ZN(n9665) );
  MOAI22 U18587 ( .A1(n28905), .A2(n1462), .B1(ram[5425]), .B2(n1463), 
        .ZN(n9666) );
  MOAI22 U18588 ( .A1(n28670), .A2(n1462), .B1(ram[5426]), .B2(n1463), 
        .ZN(n9667) );
  MOAI22 U18589 ( .A1(n28435), .A2(n1462), .B1(ram[5427]), .B2(n1463), 
        .ZN(n9668) );
  MOAI22 U18590 ( .A1(n28200), .A2(n1462), .B1(ram[5428]), .B2(n1463), 
        .ZN(n9669) );
  MOAI22 U18591 ( .A1(n27965), .A2(n1462), .B1(ram[5429]), .B2(n1463), 
        .ZN(n9670) );
  MOAI22 U18592 ( .A1(n27730), .A2(n1462), .B1(ram[5430]), .B2(n1463), 
        .ZN(n9671) );
  MOAI22 U18593 ( .A1(n27495), .A2(n1462), .B1(ram[5431]), .B2(n1463), 
        .ZN(n9672) );
  MOAI22 U18594 ( .A1(n29140), .A2(n1464), .B1(ram[5432]), .B2(n1465), 
        .ZN(n9673) );
  MOAI22 U18595 ( .A1(n28905), .A2(n1464), .B1(ram[5433]), .B2(n1465), 
        .ZN(n9674) );
  MOAI22 U18596 ( .A1(n28670), .A2(n1464), .B1(ram[5434]), .B2(n1465), 
        .ZN(n9675) );
  MOAI22 U18597 ( .A1(n28435), .A2(n1464), .B1(ram[5435]), .B2(n1465), 
        .ZN(n9676) );
  MOAI22 U18598 ( .A1(n28200), .A2(n1464), .B1(ram[5436]), .B2(n1465), 
        .ZN(n9677) );
  MOAI22 U18599 ( .A1(n27965), .A2(n1464), .B1(ram[5437]), .B2(n1465), 
        .ZN(n9678) );
  MOAI22 U18600 ( .A1(n27730), .A2(n1464), .B1(ram[5438]), .B2(n1465), 
        .ZN(n9679) );
  MOAI22 U18601 ( .A1(n27495), .A2(n1464), .B1(ram[5439]), .B2(n1465), 
        .ZN(n9680) );
  MOAI22 U18602 ( .A1(n29140), .A2(n1466), .B1(ram[5440]), .B2(n1467), 
        .ZN(n9681) );
  MOAI22 U18603 ( .A1(n28905), .A2(n1466), .B1(ram[5441]), .B2(n1467), 
        .ZN(n9682) );
  MOAI22 U18604 ( .A1(n28670), .A2(n1466), .B1(ram[5442]), .B2(n1467), 
        .ZN(n9683) );
  MOAI22 U18605 ( .A1(n28435), .A2(n1466), .B1(ram[5443]), .B2(n1467), 
        .ZN(n9684) );
  MOAI22 U18606 ( .A1(n28200), .A2(n1466), .B1(ram[5444]), .B2(n1467), 
        .ZN(n9685) );
  MOAI22 U18607 ( .A1(n27965), .A2(n1466), .B1(ram[5445]), .B2(n1467), 
        .ZN(n9686) );
  MOAI22 U18608 ( .A1(n27730), .A2(n1466), .B1(ram[5446]), .B2(n1467), 
        .ZN(n9687) );
  MOAI22 U18609 ( .A1(n27495), .A2(n1466), .B1(ram[5447]), .B2(n1467), 
        .ZN(n9688) );
  MOAI22 U18610 ( .A1(n29140), .A2(n1468), .B1(ram[5448]), .B2(n1469), 
        .ZN(n9689) );
  MOAI22 U18611 ( .A1(n28905), .A2(n1468), .B1(ram[5449]), .B2(n1469), 
        .ZN(n9690) );
  MOAI22 U18612 ( .A1(n28670), .A2(n1468), .B1(ram[5450]), .B2(n1469), 
        .ZN(n9691) );
  MOAI22 U18613 ( .A1(n28435), .A2(n1468), .B1(ram[5451]), .B2(n1469), 
        .ZN(n9692) );
  MOAI22 U18614 ( .A1(n28200), .A2(n1468), .B1(ram[5452]), .B2(n1469), 
        .ZN(n9693) );
  MOAI22 U18615 ( .A1(n27965), .A2(n1468), .B1(ram[5453]), .B2(n1469), 
        .ZN(n9694) );
  MOAI22 U18616 ( .A1(n27730), .A2(n1468), .B1(ram[5454]), .B2(n1469), 
        .ZN(n9695) );
  MOAI22 U18617 ( .A1(n27495), .A2(n1468), .B1(ram[5455]), .B2(n1469), 
        .ZN(n9696) );
  MOAI22 U18618 ( .A1(n29140), .A2(n1470), .B1(ram[5456]), .B2(n1471), 
        .ZN(n9697) );
  MOAI22 U18619 ( .A1(n28905), .A2(n1470), .B1(ram[5457]), .B2(n1471), 
        .ZN(n9698) );
  MOAI22 U18620 ( .A1(n28670), .A2(n1470), .B1(ram[5458]), .B2(n1471), 
        .ZN(n9699) );
  MOAI22 U18621 ( .A1(n28435), .A2(n1470), .B1(ram[5459]), .B2(n1471), 
        .ZN(n9700) );
  MOAI22 U18622 ( .A1(n28200), .A2(n1470), .B1(ram[5460]), .B2(n1471), 
        .ZN(n9701) );
  MOAI22 U18623 ( .A1(n27965), .A2(n1470), .B1(ram[5461]), .B2(n1471), 
        .ZN(n9702) );
  MOAI22 U18624 ( .A1(n27730), .A2(n1470), .B1(ram[5462]), .B2(n1471), 
        .ZN(n9703) );
  MOAI22 U18625 ( .A1(n27495), .A2(n1470), .B1(ram[5463]), .B2(n1471), 
        .ZN(n9704) );
  MOAI22 U18626 ( .A1(n29140), .A2(n1472), .B1(ram[5464]), .B2(n1473), 
        .ZN(n9705) );
  MOAI22 U18627 ( .A1(n28905), .A2(n1472), .B1(ram[5465]), .B2(n1473), 
        .ZN(n9706) );
  MOAI22 U18628 ( .A1(n28670), .A2(n1472), .B1(ram[5466]), .B2(n1473), 
        .ZN(n9707) );
  MOAI22 U18629 ( .A1(n28435), .A2(n1472), .B1(ram[5467]), .B2(n1473), 
        .ZN(n9708) );
  MOAI22 U18630 ( .A1(n28200), .A2(n1472), .B1(ram[5468]), .B2(n1473), 
        .ZN(n9709) );
  MOAI22 U18631 ( .A1(n27965), .A2(n1472), .B1(ram[5469]), .B2(n1473), 
        .ZN(n9710) );
  MOAI22 U18632 ( .A1(n27730), .A2(n1472), .B1(ram[5470]), .B2(n1473), 
        .ZN(n9711) );
  MOAI22 U18633 ( .A1(n27495), .A2(n1472), .B1(ram[5471]), .B2(n1473), 
        .ZN(n9712) );
  MOAI22 U18634 ( .A1(n29140), .A2(n1474), .B1(ram[5472]), .B2(n1475), 
        .ZN(n9713) );
  MOAI22 U18635 ( .A1(n28905), .A2(n1474), .B1(ram[5473]), .B2(n1475), 
        .ZN(n9714) );
  MOAI22 U18636 ( .A1(n28670), .A2(n1474), .B1(ram[5474]), .B2(n1475), 
        .ZN(n9715) );
  MOAI22 U18637 ( .A1(n28435), .A2(n1474), .B1(ram[5475]), .B2(n1475), 
        .ZN(n9716) );
  MOAI22 U18638 ( .A1(n28200), .A2(n1474), .B1(ram[5476]), .B2(n1475), 
        .ZN(n9717) );
  MOAI22 U18639 ( .A1(n27965), .A2(n1474), .B1(ram[5477]), .B2(n1475), 
        .ZN(n9718) );
  MOAI22 U18640 ( .A1(n27730), .A2(n1474), .B1(ram[5478]), .B2(n1475), 
        .ZN(n9719) );
  MOAI22 U18641 ( .A1(n27495), .A2(n1474), .B1(ram[5479]), .B2(n1475), 
        .ZN(n9720) );
  MOAI22 U18642 ( .A1(n29140), .A2(n1476), .B1(ram[5480]), .B2(n1477), 
        .ZN(n9721) );
  MOAI22 U18643 ( .A1(n28905), .A2(n1476), .B1(ram[5481]), .B2(n1477), 
        .ZN(n9722) );
  MOAI22 U18644 ( .A1(n28670), .A2(n1476), .B1(ram[5482]), .B2(n1477), 
        .ZN(n9723) );
  MOAI22 U18645 ( .A1(n28435), .A2(n1476), .B1(ram[5483]), .B2(n1477), 
        .ZN(n9724) );
  MOAI22 U18646 ( .A1(n28200), .A2(n1476), .B1(ram[5484]), .B2(n1477), 
        .ZN(n9725) );
  MOAI22 U18647 ( .A1(n27965), .A2(n1476), .B1(ram[5485]), .B2(n1477), 
        .ZN(n9726) );
  MOAI22 U18648 ( .A1(n27730), .A2(n1476), .B1(ram[5486]), .B2(n1477), 
        .ZN(n9727) );
  MOAI22 U18649 ( .A1(n27495), .A2(n1476), .B1(ram[5487]), .B2(n1477), 
        .ZN(n9728) );
  MOAI22 U18650 ( .A1(n29140), .A2(n1478), .B1(ram[5488]), .B2(n1479), 
        .ZN(n9729) );
  MOAI22 U18651 ( .A1(n28905), .A2(n1478), .B1(ram[5489]), .B2(n1479), 
        .ZN(n9730) );
  MOAI22 U18652 ( .A1(n28670), .A2(n1478), .B1(ram[5490]), .B2(n1479), 
        .ZN(n9731) );
  MOAI22 U18653 ( .A1(n28435), .A2(n1478), .B1(ram[5491]), .B2(n1479), 
        .ZN(n9732) );
  MOAI22 U18654 ( .A1(n28200), .A2(n1478), .B1(ram[5492]), .B2(n1479), 
        .ZN(n9733) );
  MOAI22 U18655 ( .A1(n27965), .A2(n1478), .B1(ram[5493]), .B2(n1479), 
        .ZN(n9734) );
  MOAI22 U18656 ( .A1(n27730), .A2(n1478), .B1(ram[5494]), .B2(n1479), 
        .ZN(n9735) );
  MOAI22 U18657 ( .A1(n27495), .A2(n1478), .B1(ram[5495]), .B2(n1479), 
        .ZN(n9736) );
  MOAI22 U18658 ( .A1(n29140), .A2(n1480), .B1(ram[5496]), .B2(n1481), 
        .ZN(n9737) );
  MOAI22 U18659 ( .A1(n28905), .A2(n1480), .B1(ram[5497]), .B2(n1481), 
        .ZN(n9738) );
  MOAI22 U18660 ( .A1(n28670), .A2(n1480), .B1(ram[5498]), .B2(n1481), 
        .ZN(n9739) );
  MOAI22 U18661 ( .A1(n28435), .A2(n1480), .B1(ram[5499]), .B2(n1481), 
        .ZN(n9740) );
  MOAI22 U18662 ( .A1(n28200), .A2(n1480), .B1(ram[5500]), .B2(n1481), 
        .ZN(n9741) );
  MOAI22 U18663 ( .A1(n27965), .A2(n1480), .B1(ram[5501]), .B2(n1481), 
        .ZN(n9742) );
  MOAI22 U18664 ( .A1(n27730), .A2(n1480), .B1(ram[5502]), .B2(n1481), 
        .ZN(n9743) );
  MOAI22 U18665 ( .A1(n27495), .A2(n1480), .B1(ram[5503]), .B2(n1481), 
        .ZN(n9744) );
  MOAI22 U18666 ( .A1(n29140), .A2(n1482), .B1(ram[5504]), .B2(n1483), 
        .ZN(n9745) );
  MOAI22 U18667 ( .A1(n28905), .A2(n1482), .B1(ram[5505]), .B2(n1483), 
        .ZN(n9746) );
  MOAI22 U18668 ( .A1(n28670), .A2(n1482), .B1(ram[5506]), .B2(n1483), 
        .ZN(n9747) );
  MOAI22 U18669 ( .A1(n28435), .A2(n1482), .B1(ram[5507]), .B2(n1483), 
        .ZN(n9748) );
  MOAI22 U18670 ( .A1(n28200), .A2(n1482), .B1(ram[5508]), .B2(n1483), 
        .ZN(n9749) );
  MOAI22 U18671 ( .A1(n27965), .A2(n1482), .B1(ram[5509]), .B2(n1483), 
        .ZN(n9750) );
  MOAI22 U18672 ( .A1(n27730), .A2(n1482), .B1(ram[5510]), .B2(n1483), 
        .ZN(n9751) );
  MOAI22 U18673 ( .A1(n27495), .A2(n1482), .B1(ram[5511]), .B2(n1483), 
        .ZN(n9752) );
  MOAI22 U18674 ( .A1(n29141), .A2(n1484), .B1(ram[5512]), .B2(n1485), 
        .ZN(n9753) );
  MOAI22 U18675 ( .A1(n28906), .A2(n1484), .B1(ram[5513]), .B2(n1485), 
        .ZN(n9754) );
  MOAI22 U18676 ( .A1(n28671), .A2(n1484), .B1(ram[5514]), .B2(n1485), 
        .ZN(n9755) );
  MOAI22 U18677 ( .A1(n28436), .A2(n1484), .B1(ram[5515]), .B2(n1485), 
        .ZN(n9756) );
  MOAI22 U18678 ( .A1(n28201), .A2(n1484), .B1(ram[5516]), .B2(n1485), 
        .ZN(n9757) );
  MOAI22 U18679 ( .A1(n27966), .A2(n1484), .B1(ram[5517]), .B2(n1485), 
        .ZN(n9758) );
  MOAI22 U18680 ( .A1(n27731), .A2(n1484), .B1(ram[5518]), .B2(n1485), 
        .ZN(n9759) );
  MOAI22 U18681 ( .A1(n27496), .A2(n1484), .B1(ram[5519]), .B2(n1485), 
        .ZN(n9760) );
  MOAI22 U18682 ( .A1(n29141), .A2(n1486), .B1(ram[5520]), .B2(n1487), 
        .ZN(n9761) );
  MOAI22 U18683 ( .A1(n28906), .A2(n1486), .B1(ram[5521]), .B2(n1487), 
        .ZN(n9762) );
  MOAI22 U18684 ( .A1(n28671), .A2(n1486), .B1(ram[5522]), .B2(n1487), 
        .ZN(n9763) );
  MOAI22 U18685 ( .A1(n28436), .A2(n1486), .B1(ram[5523]), .B2(n1487), 
        .ZN(n9764) );
  MOAI22 U18686 ( .A1(n28201), .A2(n1486), .B1(ram[5524]), .B2(n1487), 
        .ZN(n9765) );
  MOAI22 U18687 ( .A1(n27966), .A2(n1486), .B1(ram[5525]), .B2(n1487), 
        .ZN(n9766) );
  MOAI22 U18688 ( .A1(n27731), .A2(n1486), .B1(ram[5526]), .B2(n1487), 
        .ZN(n9767) );
  MOAI22 U18689 ( .A1(n27496), .A2(n1486), .B1(ram[5527]), .B2(n1487), 
        .ZN(n9768) );
  MOAI22 U18690 ( .A1(n29141), .A2(n1488), .B1(ram[5528]), .B2(n1489), 
        .ZN(n9769) );
  MOAI22 U18691 ( .A1(n28906), .A2(n1488), .B1(ram[5529]), .B2(n1489), 
        .ZN(n9770) );
  MOAI22 U18692 ( .A1(n28671), .A2(n1488), .B1(ram[5530]), .B2(n1489), 
        .ZN(n9771) );
  MOAI22 U18693 ( .A1(n28436), .A2(n1488), .B1(ram[5531]), .B2(n1489), 
        .ZN(n9772) );
  MOAI22 U18694 ( .A1(n28201), .A2(n1488), .B1(ram[5532]), .B2(n1489), 
        .ZN(n9773) );
  MOAI22 U18695 ( .A1(n27966), .A2(n1488), .B1(ram[5533]), .B2(n1489), 
        .ZN(n9774) );
  MOAI22 U18696 ( .A1(n27731), .A2(n1488), .B1(ram[5534]), .B2(n1489), 
        .ZN(n9775) );
  MOAI22 U18697 ( .A1(n27496), .A2(n1488), .B1(ram[5535]), .B2(n1489), 
        .ZN(n9776) );
  MOAI22 U18698 ( .A1(n29141), .A2(n1490), .B1(ram[5536]), .B2(n1491), 
        .ZN(n9777) );
  MOAI22 U18699 ( .A1(n28906), .A2(n1490), .B1(ram[5537]), .B2(n1491), 
        .ZN(n9778) );
  MOAI22 U18700 ( .A1(n28671), .A2(n1490), .B1(ram[5538]), .B2(n1491), 
        .ZN(n9779) );
  MOAI22 U18701 ( .A1(n28436), .A2(n1490), .B1(ram[5539]), .B2(n1491), 
        .ZN(n9780) );
  MOAI22 U18702 ( .A1(n28201), .A2(n1490), .B1(ram[5540]), .B2(n1491), 
        .ZN(n9781) );
  MOAI22 U18703 ( .A1(n27966), .A2(n1490), .B1(ram[5541]), .B2(n1491), 
        .ZN(n9782) );
  MOAI22 U18704 ( .A1(n27731), .A2(n1490), .B1(ram[5542]), .B2(n1491), 
        .ZN(n9783) );
  MOAI22 U18705 ( .A1(n27496), .A2(n1490), .B1(ram[5543]), .B2(n1491), 
        .ZN(n9784) );
  MOAI22 U18706 ( .A1(n29141), .A2(n1492), .B1(ram[5544]), .B2(n1493), 
        .ZN(n9785) );
  MOAI22 U18707 ( .A1(n28906), .A2(n1492), .B1(ram[5545]), .B2(n1493), 
        .ZN(n9786) );
  MOAI22 U18708 ( .A1(n28671), .A2(n1492), .B1(ram[5546]), .B2(n1493), 
        .ZN(n9787) );
  MOAI22 U18709 ( .A1(n28436), .A2(n1492), .B1(ram[5547]), .B2(n1493), 
        .ZN(n9788) );
  MOAI22 U18710 ( .A1(n28201), .A2(n1492), .B1(ram[5548]), .B2(n1493), 
        .ZN(n9789) );
  MOAI22 U18711 ( .A1(n27966), .A2(n1492), .B1(ram[5549]), .B2(n1493), 
        .ZN(n9790) );
  MOAI22 U18712 ( .A1(n27731), .A2(n1492), .B1(ram[5550]), .B2(n1493), 
        .ZN(n9791) );
  MOAI22 U18713 ( .A1(n27496), .A2(n1492), .B1(ram[5551]), .B2(n1493), 
        .ZN(n9792) );
  MOAI22 U18714 ( .A1(n29141), .A2(n1494), .B1(ram[5552]), .B2(n1495), 
        .ZN(n9793) );
  MOAI22 U18715 ( .A1(n28906), .A2(n1494), .B1(ram[5553]), .B2(n1495), 
        .ZN(n9794) );
  MOAI22 U18716 ( .A1(n28671), .A2(n1494), .B1(ram[5554]), .B2(n1495), 
        .ZN(n9795) );
  MOAI22 U18717 ( .A1(n28436), .A2(n1494), .B1(ram[5555]), .B2(n1495), 
        .ZN(n9796) );
  MOAI22 U18718 ( .A1(n28201), .A2(n1494), .B1(ram[5556]), .B2(n1495), 
        .ZN(n9797) );
  MOAI22 U18719 ( .A1(n27966), .A2(n1494), .B1(ram[5557]), .B2(n1495), 
        .ZN(n9798) );
  MOAI22 U18720 ( .A1(n27731), .A2(n1494), .B1(ram[5558]), .B2(n1495), 
        .ZN(n9799) );
  MOAI22 U18721 ( .A1(n27496), .A2(n1494), .B1(ram[5559]), .B2(n1495), 
        .ZN(n9800) );
  MOAI22 U18722 ( .A1(n29141), .A2(n1496), .B1(ram[5560]), .B2(n1497), 
        .ZN(n9801) );
  MOAI22 U18723 ( .A1(n28906), .A2(n1496), .B1(ram[5561]), .B2(n1497), 
        .ZN(n9802) );
  MOAI22 U18724 ( .A1(n28671), .A2(n1496), .B1(ram[5562]), .B2(n1497), 
        .ZN(n9803) );
  MOAI22 U18725 ( .A1(n28436), .A2(n1496), .B1(ram[5563]), .B2(n1497), 
        .ZN(n9804) );
  MOAI22 U18726 ( .A1(n28201), .A2(n1496), .B1(ram[5564]), .B2(n1497), 
        .ZN(n9805) );
  MOAI22 U18727 ( .A1(n27966), .A2(n1496), .B1(ram[5565]), .B2(n1497), 
        .ZN(n9806) );
  MOAI22 U18728 ( .A1(n27731), .A2(n1496), .B1(ram[5566]), .B2(n1497), 
        .ZN(n9807) );
  MOAI22 U18729 ( .A1(n27496), .A2(n1496), .B1(ram[5567]), .B2(n1497), 
        .ZN(n9808) );
  MOAI22 U18730 ( .A1(n29141), .A2(n1498), .B1(ram[5568]), .B2(n1499), 
        .ZN(n9809) );
  MOAI22 U18731 ( .A1(n28906), .A2(n1498), .B1(ram[5569]), .B2(n1499), 
        .ZN(n9810) );
  MOAI22 U18732 ( .A1(n28671), .A2(n1498), .B1(ram[5570]), .B2(n1499), 
        .ZN(n9811) );
  MOAI22 U18733 ( .A1(n28436), .A2(n1498), .B1(ram[5571]), .B2(n1499), 
        .ZN(n9812) );
  MOAI22 U18734 ( .A1(n28201), .A2(n1498), .B1(ram[5572]), .B2(n1499), 
        .ZN(n9813) );
  MOAI22 U18735 ( .A1(n27966), .A2(n1498), .B1(ram[5573]), .B2(n1499), 
        .ZN(n9814) );
  MOAI22 U18736 ( .A1(n27731), .A2(n1498), .B1(ram[5574]), .B2(n1499), 
        .ZN(n9815) );
  MOAI22 U18737 ( .A1(n27496), .A2(n1498), .B1(ram[5575]), .B2(n1499), 
        .ZN(n9816) );
  MOAI22 U18738 ( .A1(n29141), .A2(n1500), .B1(ram[5576]), .B2(n1501), 
        .ZN(n9817) );
  MOAI22 U18739 ( .A1(n28906), .A2(n1500), .B1(ram[5577]), .B2(n1501), 
        .ZN(n9818) );
  MOAI22 U18740 ( .A1(n28671), .A2(n1500), .B1(ram[5578]), .B2(n1501), 
        .ZN(n9819) );
  MOAI22 U18741 ( .A1(n28436), .A2(n1500), .B1(ram[5579]), .B2(n1501), 
        .ZN(n9820) );
  MOAI22 U18742 ( .A1(n28201), .A2(n1500), .B1(ram[5580]), .B2(n1501), 
        .ZN(n9821) );
  MOAI22 U18743 ( .A1(n27966), .A2(n1500), .B1(ram[5581]), .B2(n1501), 
        .ZN(n9822) );
  MOAI22 U18744 ( .A1(n27731), .A2(n1500), .B1(ram[5582]), .B2(n1501), 
        .ZN(n9823) );
  MOAI22 U18745 ( .A1(n27496), .A2(n1500), .B1(ram[5583]), .B2(n1501), 
        .ZN(n9824) );
  MOAI22 U18746 ( .A1(n29141), .A2(n1502), .B1(ram[5584]), .B2(n1503), 
        .ZN(n9825) );
  MOAI22 U18747 ( .A1(n28906), .A2(n1502), .B1(ram[5585]), .B2(n1503), 
        .ZN(n9826) );
  MOAI22 U18748 ( .A1(n28671), .A2(n1502), .B1(ram[5586]), .B2(n1503), 
        .ZN(n9827) );
  MOAI22 U18749 ( .A1(n28436), .A2(n1502), .B1(ram[5587]), .B2(n1503), 
        .ZN(n9828) );
  MOAI22 U18750 ( .A1(n28201), .A2(n1502), .B1(ram[5588]), .B2(n1503), 
        .ZN(n9829) );
  MOAI22 U18751 ( .A1(n27966), .A2(n1502), .B1(ram[5589]), .B2(n1503), 
        .ZN(n9830) );
  MOAI22 U18752 ( .A1(n27731), .A2(n1502), .B1(ram[5590]), .B2(n1503), 
        .ZN(n9831) );
  MOAI22 U18753 ( .A1(n27496), .A2(n1502), .B1(ram[5591]), .B2(n1503), 
        .ZN(n9832) );
  MOAI22 U18754 ( .A1(n29141), .A2(n1504), .B1(ram[5592]), .B2(n1505), 
        .ZN(n9833) );
  MOAI22 U18755 ( .A1(n28906), .A2(n1504), .B1(ram[5593]), .B2(n1505), 
        .ZN(n9834) );
  MOAI22 U18756 ( .A1(n28671), .A2(n1504), .B1(ram[5594]), .B2(n1505), 
        .ZN(n9835) );
  MOAI22 U18757 ( .A1(n28436), .A2(n1504), .B1(ram[5595]), .B2(n1505), 
        .ZN(n9836) );
  MOAI22 U18758 ( .A1(n28201), .A2(n1504), .B1(ram[5596]), .B2(n1505), 
        .ZN(n9837) );
  MOAI22 U18759 ( .A1(n27966), .A2(n1504), .B1(ram[5597]), .B2(n1505), 
        .ZN(n9838) );
  MOAI22 U18760 ( .A1(n27731), .A2(n1504), .B1(ram[5598]), .B2(n1505), 
        .ZN(n9839) );
  MOAI22 U18761 ( .A1(n27496), .A2(n1504), .B1(ram[5599]), .B2(n1505), 
        .ZN(n9840) );
  MOAI22 U18762 ( .A1(n29141), .A2(n1506), .B1(ram[5600]), .B2(n1507), 
        .ZN(n9841) );
  MOAI22 U18763 ( .A1(n28906), .A2(n1506), .B1(ram[5601]), .B2(n1507), 
        .ZN(n9842) );
  MOAI22 U18764 ( .A1(n28671), .A2(n1506), .B1(ram[5602]), .B2(n1507), 
        .ZN(n9843) );
  MOAI22 U18765 ( .A1(n28436), .A2(n1506), .B1(ram[5603]), .B2(n1507), 
        .ZN(n9844) );
  MOAI22 U18766 ( .A1(n28201), .A2(n1506), .B1(ram[5604]), .B2(n1507), 
        .ZN(n9845) );
  MOAI22 U18767 ( .A1(n27966), .A2(n1506), .B1(ram[5605]), .B2(n1507), 
        .ZN(n9846) );
  MOAI22 U18768 ( .A1(n27731), .A2(n1506), .B1(ram[5606]), .B2(n1507), 
        .ZN(n9847) );
  MOAI22 U18769 ( .A1(n27496), .A2(n1506), .B1(ram[5607]), .B2(n1507), 
        .ZN(n9848) );
  MOAI22 U18770 ( .A1(n29141), .A2(n1508), .B1(ram[5608]), .B2(n1509), 
        .ZN(n9849) );
  MOAI22 U18771 ( .A1(n28906), .A2(n1508), .B1(ram[5609]), .B2(n1509), 
        .ZN(n9850) );
  MOAI22 U18772 ( .A1(n28671), .A2(n1508), .B1(ram[5610]), .B2(n1509), 
        .ZN(n9851) );
  MOAI22 U18773 ( .A1(n28436), .A2(n1508), .B1(ram[5611]), .B2(n1509), 
        .ZN(n9852) );
  MOAI22 U18774 ( .A1(n28201), .A2(n1508), .B1(ram[5612]), .B2(n1509), 
        .ZN(n9853) );
  MOAI22 U18775 ( .A1(n27966), .A2(n1508), .B1(ram[5613]), .B2(n1509), 
        .ZN(n9854) );
  MOAI22 U18776 ( .A1(n27731), .A2(n1508), .B1(ram[5614]), .B2(n1509), 
        .ZN(n9855) );
  MOAI22 U18777 ( .A1(n27496), .A2(n1508), .B1(ram[5615]), .B2(n1509), 
        .ZN(n9856) );
  MOAI22 U18778 ( .A1(n29142), .A2(n1510), .B1(ram[5616]), .B2(n1511), 
        .ZN(n9857) );
  MOAI22 U18779 ( .A1(n28907), .A2(n1510), .B1(ram[5617]), .B2(n1511), 
        .ZN(n9858) );
  MOAI22 U18780 ( .A1(n28672), .A2(n1510), .B1(ram[5618]), .B2(n1511), 
        .ZN(n9859) );
  MOAI22 U18781 ( .A1(n28437), .A2(n1510), .B1(ram[5619]), .B2(n1511), 
        .ZN(n9860) );
  MOAI22 U18782 ( .A1(n28202), .A2(n1510), .B1(ram[5620]), .B2(n1511), 
        .ZN(n9861) );
  MOAI22 U18783 ( .A1(n27967), .A2(n1510), .B1(ram[5621]), .B2(n1511), 
        .ZN(n9862) );
  MOAI22 U18784 ( .A1(n27732), .A2(n1510), .B1(ram[5622]), .B2(n1511), 
        .ZN(n9863) );
  MOAI22 U18785 ( .A1(n27497), .A2(n1510), .B1(ram[5623]), .B2(n1511), 
        .ZN(n9864) );
  MOAI22 U18786 ( .A1(n29142), .A2(n1512), .B1(ram[5624]), .B2(n1513), 
        .ZN(n9865) );
  MOAI22 U18787 ( .A1(n28907), .A2(n1512), .B1(ram[5625]), .B2(n1513), 
        .ZN(n9866) );
  MOAI22 U18788 ( .A1(n28672), .A2(n1512), .B1(ram[5626]), .B2(n1513), 
        .ZN(n9867) );
  MOAI22 U18789 ( .A1(n28437), .A2(n1512), .B1(ram[5627]), .B2(n1513), 
        .ZN(n9868) );
  MOAI22 U18790 ( .A1(n28202), .A2(n1512), .B1(ram[5628]), .B2(n1513), 
        .ZN(n9869) );
  MOAI22 U18791 ( .A1(n27967), .A2(n1512), .B1(ram[5629]), .B2(n1513), 
        .ZN(n9870) );
  MOAI22 U18792 ( .A1(n27732), .A2(n1512), .B1(ram[5630]), .B2(n1513), 
        .ZN(n9871) );
  MOAI22 U18793 ( .A1(n27497), .A2(n1512), .B1(ram[5631]), .B2(n1513), 
        .ZN(n9872) );
  MOAI22 U18794 ( .A1(n29142), .A2(n1514), .B1(ram[5632]), .B2(n1515), 
        .ZN(n9873) );
  MOAI22 U18795 ( .A1(n28907), .A2(n1514), .B1(ram[5633]), .B2(n1515), 
        .ZN(n9874) );
  MOAI22 U18796 ( .A1(n28672), .A2(n1514), .B1(ram[5634]), .B2(n1515), 
        .ZN(n9875) );
  MOAI22 U18797 ( .A1(n28437), .A2(n1514), .B1(ram[5635]), .B2(n1515), 
        .ZN(n9876) );
  MOAI22 U18798 ( .A1(n28202), .A2(n1514), .B1(ram[5636]), .B2(n1515), 
        .ZN(n9877) );
  MOAI22 U18799 ( .A1(n27967), .A2(n1514), .B1(ram[5637]), .B2(n1515), 
        .ZN(n9878) );
  MOAI22 U18800 ( .A1(n27732), .A2(n1514), .B1(ram[5638]), .B2(n1515), 
        .ZN(n9879) );
  MOAI22 U18801 ( .A1(n27497), .A2(n1514), .B1(ram[5639]), .B2(n1515), 
        .ZN(n9880) );
  MOAI22 U18802 ( .A1(n29142), .A2(n1517), .B1(ram[5640]), .B2(n1518), 
        .ZN(n9881) );
  MOAI22 U18803 ( .A1(n28907), .A2(n1517), .B1(ram[5641]), .B2(n1518), 
        .ZN(n9882) );
  MOAI22 U18804 ( .A1(n28672), .A2(n1517), .B1(ram[5642]), .B2(n1518), 
        .ZN(n9883) );
  MOAI22 U18805 ( .A1(n28437), .A2(n1517), .B1(ram[5643]), .B2(n1518), 
        .ZN(n9884) );
  MOAI22 U18806 ( .A1(n28202), .A2(n1517), .B1(ram[5644]), .B2(n1518), 
        .ZN(n9885) );
  MOAI22 U18807 ( .A1(n27967), .A2(n1517), .B1(ram[5645]), .B2(n1518), 
        .ZN(n9886) );
  MOAI22 U18808 ( .A1(n27732), .A2(n1517), .B1(ram[5646]), .B2(n1518), 
        .ZN(n9887) );
  MOAI22 U18809 ( .A1(n27497), .A2(n1517), .B1(ram[5647]), .B2(n1518), 
        .ZN(n9888) );
  MOAI22 U18810 ( .A1(n29142), .A2(n1519), .B1(ram[5648]), .B2(n1520), 
        .ZN(n9889) );
  MOAI22 U18811 ( .A1(n28907), .A2(n1519), .B1(ram[5649]), .B2(n1520), 
        .ZN(n9890) );
  MOAI22 U18812 ( .A1(n28672), .A2(n1519), .B1(ram[5650]), .B2(n1520), 
        .ZN(n9891) );
  MOAI22 U18813 ( .A1(n28437), .A2(n1519), .B1(ram[5651]), .B2(n1520), 
        .ZN(n9892) );
  MOAI22 U18814 ( .A1(n28202), .A2(n1519), .B1(ram[5652]), .B2(n1520), 
        .ZN(n9893) );
  MOAI22 U18815 ( .A1(n27967), .A2(n1519), .B1(ram[5653]), .B2(n1520), 
        .ZN(n9894) );
  MOAI22 U18816 ( .A1(n27732), .A2(n1519), .B1(ram[5654]), .B2(n1520), 
        .ZN(n9895) );
  MOAI22 U18817 ( .A1(n27497), .A2(n1519), .B1(ram[5655]), .B2(n1520), 
        .ZN(n9896) );
  MOAI22 U18818 ( .A1(n29142), .A2(n1521), .B1(ram[5656]), .B2(n1522), 
        .ZN(n9897) );
  MOAI22 U18819 ( .A1(n28907), .A2(n1521), .B1(ram[5657]), .B2(n1522), 
        .ZN(n9898) );
  MOAI22 U18820 ( .A1(n28672), .A2(n1521), .B1(ram[5658]), .B2(n1522), 
        .ZN(n9899) );
  MOAI22 U18821 ( .A1(n28437), .A2(n1521), .B1(ram[5659]), .B2(n1522), 
        .ZN(n9900) );
  MOAI22 U18822 ( .A1(n28202), .A2(n1521), .B1(ram[5660]), .B2(n1522), 
        .ZN(n9901) );
  MOAI22 U18823 ( .A1(n27967), .A2(n1521), .B1(ram[5661]), .B2(n1522), 
        .ZN(n9902) );
  MOAI22 U18824 ( .A1(n27732), .A2(n1521), .B1(ram[5662]), .B2(n1522), 
        .ZN(n9903) );
  MOAI22 U18825 ( .A1(n27497), .A2(n1521), .B1(ram[5663]), .B2(n1522), 
        .ZN(n9904) );
  MOAI22 U18826 ( .A1(n29142), .A2(n1523), .B1(ram[5664]), .B2(n1524), 
        .ZN(n9905) );
  MOAI22 U18827 ( .A1(n28907), .A2(n1523), .B1(ram[5665]), .B2(n1524), 
        .ZN(n9906) );
  MOAI22 U18828 ( .A1(n28672), .A2(n1523), .B1(ram[5666]), .B2(n1524), 
        .ZN(n9907) );
  MOAI22 U18829 ( .A1(n28437), .A2(n1523), .B1(ram[5667]), .B2(n1524), 
        .ZN(n9908) );
  MOAI22 U18830 ( .A1(n28202), .A2(n1523), .B1(ram[5668]), .B2(n1524), 
        .ZN(n9909) );
  MOAI22 U18831 ( .A1(n27967), .A2(n1523), .B1(ram[5669]), .B2(n1524), 
        .ZN(n9910) );
  MOAI22 U18832 ( .A1(n27732), .A2(n1523), .B1(ram[5670]), .B2(n1524), 
        .ZN(n9911) );
  MOAI22 U18833 ( .A1(n27497), .A2(n1523), .B1(ram[5671]), .B2(n1524), 
        .ZN(n9912) );
  MOAI22 U18834 ( .A1(n29142), .A2(n1525), .B1(ram[5672]), .B2(n1526), 
        .ZN(n9913) );
  MOAI22 U18835 ( .A1(n28907), .A2(n1525), .B1(ram[5673]), .B2(n1526), 
        .ZN(n9914) );
  MOAI22 U18836 ( .A1(n28672), .A2(n1525), .B1(ram[5674]), .B2(n1526), 
        .ZN(n9915) );
  MOAI22 U18837 ( .A1(n28437), .A2(n1525), .B1(ram[5675]), .B2(n1526), 
        .ZN(n9916) );
  MOAI22 U18838 ( .A1(n28202), .A2(n1525), .B1(ram[5676]), .B2(n1526), 
        .ZN(n9917) );
  MOAI22 U18839 ( .A1(n27967), .A2(n1525), .B1(ram[5677]), .B2(n1526), 
        .ZN(n9918) );
  MOAI22 U18840 ( .A1(n27732), .A2(n1525), .B1(ram[5678]), .B2(n1526), 
        .ZN(n9919) );
  MOAI22 U18841 ( .A1(n27497), .A2(n1525), .B1(ram[5679]), .B2(n1526), 
        .ZN(n9920) );
  MOAI22 U18842 ( .A1(n29142), .A2(n1527), .B1(ram[5680]), .B2(n1528), 
        .ZN(n9921) );
  MOAI22 U18843 ( .A1(n28907), .A2(n1527), .B1(ram[5681]), .B2(n1528), 
        .ZN(n9922) );
  MOAI22 U18844 ( .A1(n28672), .A2(n1527), .B1(ram[5682]), .B2(n1528), 
        .ZN(n9923) );
  MOAI22 U18845 ( .A1(n28437), .A2(n1527), .B1(ram[5683]), .B2(n1528), 
        .ZN(n9924) );
  MOAI22 U18846 ( .A1(n28202), .A2(n1527), .B1(ram[5684]), .B2(n1528), 
        .ZN(n9925) );
  MOAI22 U18847 ( .A1(n27967), .A2(n1527), .B1(ram[5685]), .B2(n1528), 
        .ZN(n9926) );
  MOAI22 U18848 ( .A1(n27732), .A2(n1527), .B1(ram[5686]), .B2(n1528), 
        .ZN(n9927) );
  MOAI22 U18849 ( .A1(n27497), .A2(n1527), .B1(ram[5687]), .B2(n1528), 
        .ZN(n9928) );
  MOAI22 U18850 ( .A1(n29142), .A2(n1529), .B1(ram[5688]), .B2(n1530), 
        .ZN(n9929) );
  MOAI22 U18851 ( .A1(n28907), .A2(n1529), .B1(ram[5689]), .B2(n1530), 
        .ZN(n9930) );
  MOAI22 U18852 ( .A1(n28672), .A2(n1529), .B1(ram[5690]), .B2(n1530), 
        .ZN(n9931) );
  MOAI22 U18853 ( .A1(n28437), .A2(n1529), .B1(ram[5691]), .B2(n1530), 
        .ZN(n9932) );
  MOAI22 U18854 ( .A1(n28202), .A2(n1529), .B1(ram[5692]), .B2(n1530), 
        .ZN(n9933) );
  MOAI22 U18855 ( .A1(n27967), .A2(n1529), .B1(ram[5693]), .B2(n1530), 
        .ZN(n9934) );
  MOAI22 U18856 ( .A1(n27732), .A2(n1529), .B1(ram[5694]), .B2(n1530), 
        .ZN(n9935) );
  MOAI22 U18857 ( .A1(n27497), .A2(n1529), .B1(ram[5695]), .B2(n1530), 
        .ZN(n9936) );
  MOAI22 U18858 ( .A1(n29142), .A2(n1531), .B1(ram[5696]), .B2(n1532), 
        .ZN(n9937) );
  MOAI22 U18859 ( .A1(n28907), .A2(n1531), .B1(ram[5697]), .B2(n1532), 
        .ZN(n9938) );
  MOAI22 U18860 ( .A1(n28672), .A2(n1531), .B1(ram[5698]), .B2(n1532), 
        .ZN(n9939) );
  MOAI22 U18861 ( .A1(n28437), .A2(n1531), .B1(ram[5699]), .B2(n1532), 
        .ZN(n9940) );
  MOAI22 U18862 ( .A1(n28202), .A2(n1531), .B1(ram[5700]), .B2(n1532), 
        .ZN(n9941) );
  MOAI22 U18863 ( .A1(n27967), .A2(n1531), .B1(ram[5701]), .B2(n1532), 
        .ZN(n9942) );
  MOAI22 U18864 ( .A1(n27732), .A2(n1531), .B1(ram[5702]), .B2(n1532), 
        .ZN(n9943) );
  MOAI22 U18865 ( .A1(n27497), .A2(n1531), .B1(ram[5703]), .B2(n1532), 
        .ZN(n9944) );
  MOAI22 U18866 ( .A1(n29142), .A2(n1533), .B1(ram[5704]), .B2(n1534), 
        .ZN(n9945) );
  MOAI22 U18867 ( .A1(n28907), .A2(n1533), .B1(ram[5705]), .B2(n1534), 
        .ZN(n9946) );
  MOAI22 U18868 ( .A1(n28672), .A2(n1533), .B1(ram[5706]), .B2(n1534), 
        .ZN(n9947) );
  MOAI22 U18869 ( .A1(n28437), .A2(n1533), .B1(ram[5707]), .B2(n1534), 
        .ZN(n9948) );
  MOAI22 U18870 ( .A1(n28202), .A2(n1533), .B1(ram[5708]), .B2(n1534), 
        .ZN(n9949) );
  MOAI22 U18871 ( .A1(n27967), .A2(n1533), .B1(ram[5709]), .B2(n1534), 
        .ZN(n9950) );
  MOAI22 U18872 ( .A1(n27732), .A2(n1533), .B1(ram[5710]), .B2(n1534), 
        .ZN(n9951) );
  MOAI22 U18873 ( .A1(n27497), .A2(n1533), .B1(ram[5711]), .B2(n1534), 
        .ZN(n9952) );
  MOAI22 U18874 ( .A1(n29142), .A2(n1535), .B1(ram[5712]), .B2(n1536), 
        .ZN(n9953) );
  MOAI22 U18875 ( .A1(n28907), .A2(n1535), .B1(ram[5713]), .B2(n1536), 
        .ZN(n9954) );
  MOAI22 U18876 ( .A1(n28672), .A2(n1535), .B1(ram[5714]), .B2(n1536), 
        .ZN(n9955) );
  MOAI22 U18877 ( .A1(n28437), .A2(n1535), .B1(ram[5715]), .B2(n1536), 
        .ZN(n9956) );
  MOAI22 U18878 ( .A1(n28202), .A2(n1535), .B1(ram[5716]), .B2(n1536), 
        .ZN(n9957) );
  MOAI22 U18879 ( .A1(n27967), .A2(n1535), .B1(ram[5717]), .B2(n1536), 
        .ZN(n9958) );
  MOAI22 U18880 ( .A1(n27732), .A2(n1535), .B1(ram[5718]), .B2(n1536), 
        .ZN(n9959) );
  MOAI22 U18881 ( .A1(n27497), .A2(n1535), .B1(ram[5719]), .B2(n1536), 
        .ZN(n9960) );
  MOAI22 U18882 ( .A1(n29143), .A2(n1537), .B1(ram[5720]), .B2(n1538), 
        .ZN(n9961) );
  MOAI22 U18883 ( .A1(n28908), .A2(n1537), .B1(ram[5721]), .B2(n1538), 
        .ZN(n9962) );
  MOAI22 U18884 ( .A1(n28673), .A2(n1537), .B1(ram[5722]), .B2(n1538), 
        .ZN(n9963) );
  MOAI22 U18885 ( .A1(n28438), .A2(n1537), .B1(ram[5723]), .B2(n1538), 
        .ZN(n9964) );
  MOAI22 U18886 ( .A1(n28203), .A2(n1537), .B1(ram[5724]), .B2(n1538), 
        .ZN(n9965) );
  MOAI22 U18887 ( .A1(n27968), .A2(n1537), .B1(ram[5725]), .B2(n1538), 
        .ZN(n9966) );
  MOAI22 U18888 ( .A1(n27733), .A2(n1537), .B1(ram[5726]), .B2(n1538), 
        .ZN(n9967) );
  MOAI22 U18889 ( .A1(n27498), .A2(n1537), .B1(ram[5727]), .B2(n1538), 
        .ZN(n9968) );
  MOAI22 U18890 ( .A1(n29143), .A2(n1539), .B1(ram[5728]), .B2(n1540), 
        .ZN(n9969) );
  MOAI22 U18891 ( .A1(n28908), .A2(n1539), .B1(ram[5729]), .B2(n1540), 
        .ZN(n9970) );
  MOAI22 U18892 ( .A1(n28673), .A2(n1539), .B1(ram[5730]), .B2(n1540), 
        .ZN(n9971) );
  MOAI22 U18893 ( .A1(n28438), .A2(n1539), .B1(ram[5731]), .B2(n1540), 
        .ZN(n9972) );
  MOAI22 U18894 ( .A1(n28203), .A2(n1539), .B1(ram[5732]), .B2(n1540), 
        .ZN(n9973) );
  MOAI22 U18895 ( .A1(n27968), .A2(n1539), .B1(ram[5733]), .B2(n1540), 
        .ZN(n9974) );
  MOAI22 U18896 ( .A1(n27733), .A2(n1539), .B1(ram[5734]), .B2(n1540), 
        .ZN(n9975) );
  MOAI22 U18897 ( .A1(n27498), .A2(n1539), .B1(ram[5735]), .B2(n1540), 
        .ZN(n9976) );
  MOAI22 U18898 ( .A1(n29143), .A2(n1541), .B1(ram[5736]), .B2(n1542), 
        .ZN(n9977) );
  MOAI22 U18899 ( .A1(n28908), .A2(n1541), .B1(ram[5737]), .B2(n1542), 
        .ZN(n9978) );
  MOAI22 U18900 ( .A1(n28673), .A2(n1541), .B1(ram[5738]), .B2(n1542), 
        .ZN(n9979) );
  MOAI22 U18901 ( .A1(n28438), .A2(n1541), .B1(ram[5739]), .B2(n1542), 
        .ZN(n9980) );
  MOAI22 U18902 ( .A1(n28203), .A2(n1541), .B1(ram[5740]), .B2(n1542), 
        .ZN(n9981) );
  MOAI22 U18903 ( .A1(n27968), .A2(n1541), .B1(ram[5741]), .B2(n1542), 
        .ZN(n9982) );
  MOAI22 U18904 ( .A1(n27733), .A2(n1541), .B1(ram[5742]), .B2(n1542), 
        .ZN(n9983) );
  MOAI22 U18905 ( .A1(n27498), .A2(n1541), .B1(ram[5743]), .B2(n1542), 
        .ZN(n9984) );
  MOAI22 U18906 ( .A1(n29143), .A2(n1543), .B1(ram[5744]), .B2(n1544), 
        .ZN(n9985) );
  MOAI22 U18907 ( .A1(n28908), .A2(n1543), .B1(ram[5745]), .B2(n1544), 
        .ZN(n9986) );
  MOAI22 U18908 ( .A1(n28673), .A2(n1543), .B1(ram[5746]), .B2(n1544), 
        .ZN(n9987) );
  MOAI22 U18909 ( .A1(n28438), .A2(n1543), .B1(ram[5747]), .B2(n1544), 
        .ZN(n9988) );
  MOAI22 U18910 ( .A1(n28203), .A2(n1543), .B1(ram[5748]), .B2(n1544), 
        .ZN(n9989) );
  MOAI22 U18911 ( .A1(n27968), .A2(n1543), .B1(ram[5749]), .B2(n1544), 
        .ZN(n9990) );
  MOAI22 U18912 ( .A1(n27733), .A2(n1543), .B1(ram[5750]), .B2(n1544), 
        .ZN(n9991) );
  MOAI22 U18913 ( .A1(n27498), .A2(n1543), .B1(ram[5751]), .B2(n1544), 
        .ZN(n9992) );
  MOAI22 U18914 ( .A1(n29143), .A2(n1545), .B1(ram[5752]), .B2(n1546), 
        .ZN(n9993) );
  MOAI22 U18915 ( .A1(n28908), .A2(n1545), .B1(ram[5753]), .B2(n1546), 
        .ZN(n9994) );
  MOAI22 U18916 ( .A1(n28673), .A2(n1545), .B1(ram[5754]), .B2(n1546), 
        .ZN(n9995) );
  MOAI22 U18917 ( .A1(n28438), .A2(n1545), .B1(ram[5755]), .B2(n1546), 
        .ZN(n9996) );
  MOAI22 U18918 ( .A1(n28203), .A2(n1545), .B1(ram[5756]), .B2(n1546), 
        .ZN(n9997) );
  MOAI22 U18919 ( .A1(n27968), .A2(n1545), .B1(ram[5757]), .B2(n1546), 
        .ZN(n9998) );
  MOAI22 U18920 ( .A1(n27733), .A2(n1545), .B1(ram[5758]), .B2(n1546), 
        .ZN(n9999) );
  MOAI22 U18921 ( .A1(n27498), .A2(n1545), .B1(ram[5759]), .B2(n1546), 
        .ZN(n10000) );
  MOAI22 U18922 ( .A1(n29143), .A2(n1547), .B1(ram[5760]), .B2(n1548), 
        .ZN(n10001) );
  MOAI22 U18923 ( .A1(n28908), .A2(n1547), .B1(ram[5761]), .B2(n1548), 
        .ZN(n10002) );
  MOAI22 U18924 ( .A1(n28673), .A2(n1547), .B1(ram[5762]), .B2(n1548), 
        .ZN(n10003) );
  MOAI22 U18925 ( .A1(n28438), .A2(n1547), .B1(ram[5763]), .B2(n1548), 
        .ZN(n10004) );
  MOAI22 U18926 ( .A1(n28203), .A2(n1547), .B1(ram[5764]), .B2(n1548), 
        .ZN(n10005) );
  MOAI22 U18927 ( .A1(n27968), .A2(n1547), .B1(ram[5765]), .B2(n1548), 
        .ZN(n10006) );
  MOAI22 U18928 ( .A1(n27733), .A2(n1547), .B1(ram[5766]), .B2(n1548), 
        .ZN(n10007) );
  MOAI22 U18929 ( .A1(n27498), .A2(n1547), .B1(ram[5767]), .B2(n1548), 
        .ZN(n10008) );
  MOAI22 U18930 ( .A1(n29143), .A2(n1549), .B1(ram[5768]), .B2(n1550), 
        .ZN(n10009) );
  MOAI22 U18931 ( .A1(n28908), .A2(n1549), .B1(ram[5769]), .B2(n1550), 
        .ZN(n10010) );
  MOAI22 U18932 ( .A1(n28673), .A2(n1549), .B1(ram[5770]), .B2(n1550), 
        .ZN(n10011) );
  MOAI22 U18933 ( .A1(n28438), .A2(n1549), .B1(ram[5771]), .B2(n1550), 
        .ZN(n10012) );
  MOAI22 U18934 ( .A1(n28203), .A2(n1549), .B1(ram[5772]), .B2(n1550), 
        .ZN(n10013) );
  MOAI22 U18935 ( .A1(n27968), .A2(n1549), .B1(ram[5773]), .B2(n1550), 
        .ZN(n10014) );
  MOAI22 U18936 ( .A1(n27733), .A2(n1549), .B1(ram[5774]), .B2(n1550), 
        .ZN(n10015) );
  MOAI22 U18937 ( .A1(n27498), .A2(n1549), .B1(ram[5775]), .B2(n1550), 
        .ZN(n10016) );
  MOAI22 U18938 ( .A1(n29143), .A2(n1551), .B1(ram[5776]), .B2(n1552), 
        .ZN(n10017) );
  MOAI22 U18939 ( .A1(n28908), .A2(n1551), .B1(ram[5777]), .B2(n1552), 
        .ZN(n10018) );
  MOAI22 U18940 ( .A1(n28673), .A2(n1551), .B1(ram[5778]), .B2(n1552), 
        .ZN(n10019) );
  MOAI22 U18941 ( .A1(n28438), .A2(n1551), .B1(ram[5779]), .B2(n1552), 
        .ZN(n10020) );
  MOAI22 U18942 ( .A1(n28203), .A2(n1551), .B1(ram[5780]), .B2(n1552), 
        .ZN(n10021) );
  MOAI22 U18943 ( .A1(n27968), .A2(n1551), .B1(ram[5781]), .B2(n1552), 
        .ZN(n10022) );
  MOAI22 U18944 ( .A1(n27733), .A2(n1551), .B1(ram[5782]), .B2(n1552), 
        .ZN(n10023) );
  MOAI22 U18945 ( .A1(n27498), .A2(n1551), .B1(ram[5783]), .B2(n1552), 
        .ZN(n10024) );
  MOAI22 U18946 ( .A1(n29143), .A2(n1553), .B1(ram[5784]), .B2(n1554), 
        .ZN(n10025) );
  MOAI22 U18947 ( .A1(n28908), .A2(n1553), .B1(ram[5785]), .B2(n1554), 
        .ZN(n10026) );
  MOAI22 U18948 ( .A1(n28673), .A2(n1553), .B1(ram[5786]), .B2(n1554), 
        .ZN(n10027) );
  MOAI22 U18949 ( .A1(n28438), .A2(n1553), .B1(ram[5787]), .B2(n1554), 
        .ZN(n10028) );
  MOAI22 U18950 ( .A1(n28203), .A2(n1553), .B1(ram[5788]), .B2(n1554), 
        .ZN(n10029) );
  MOAI22 U18951 ( .A1(n27968), .A2(n1553), .B1(ram[5789]), .B2(n1554), 
        .ZN(n10030) );
  MOAI22 U18952 ( .A1(n27733), .A2(n1553), .B1(ram[5790]), .B2(n1554), 
        .ZN(n10031) );
  MOAI22 U18953 ( .A1(n27498), .A2(n1553), .B1(ram[5791]), .B2(n1554), 
        .ZN(n10032) );
  MOAI22 U18954 ( .A1(n29143), .A2(n1555), .B1(ram[5792]), .B2(n1556), 
        .ZN(n10033) );
  MOAI22 U18955 ( .A1(n28908), .A2(n1555), .B1(ram[5793]), .B2(n1556), 
        .ZN(n10034) );
  MOAI22 U18956 ( .A1(n28673), .A2(n1555), .B1(ram[5794]), .B2(n1556), 
        .ZN(n10035) );
  MOAI22 U18957 ( .A1(n28438), .A2(n1555), .B1(ram[5795]), .B2(n1556), 
        .ZN(n10036) );
  MOAI22 U18958 ( .A1(n28203), .A2(n1555), .B1(ram[5796]), .B2(n1556), 
        .ZN(n10037) );
  MOAI22 U18959 ( .A1(n27968), .A2(n1555), .B1(ram[5797]), .B2(n1556), 
        .ZN(n10038) );
  MOAI22 U18960 ( .A1(n27733), .A2(n1555), .B1(ram[5798]), .B2(n1556), 
        .ZN(n10039) );
  MOAI22 U18961 ( .A1(n27498), .A2(n1555), .B1(ram[5799]), .B2(n1556), 
        .ZN(n10040) );
  MOAI22 U18962 ( .A1(n29143), .A2(n1557), .B1(ram[5800]), .B2(n1558), 
        .ZN(n10041) );
  MOAI22 U18963 ( .A1(n28908), .A2(n1557), .B1(ram[5801]), .B2(n1558), 
        .ZN(n10042) );
  MOAI22 U18964 ( .A1(n28673), .A2(n1557), .B1(ram[5802]), .B2(n1558), 
        .ZN(n10043) );
  MOAI22 U18965 ( .A1(n28438), .A2(n1557), .B1(ram[5803]), .B2(n1558), 
        .ZN(n10044) );
  MOAI22 U18966 ( .A1(n28203), .A2(n1557), .B1(ram[5804]), .B2(n1558), 
        .ZN(n10045) );
  MOAI22 U18967 ( .A1(n27968), .A2(n1557), .B1(ram[5805]), .B2(n1558), 
        .ZN(n10046) );
  MOAI22 U18968 ( .A1(n27733), .A2(n1557), .B1(ram[5806]), .B2(n1558), 
        .ZN(n10047) );
  MOAI22 U18969 ( .A1(n27498), .A2(n1557), .B1(ram[5807]), .B2(n1558), 
        .ZN(n10048) );
  MOAI22 U18970 ( .A1(n29143), .A2(n1559), .B1(ram[5808]), .B2(n1560), 
        .ZN(n10049) );
  MOAI22 U18971 ( .A1(n28908), .A2(n1559), .B1(ram[5809]), .B2(n1560), 
        .ZN(n10050) );
  MOAI22 U18972 ( .A1(n28673), .A2(n1559), .B1(ram[5810]), .B2(n1560), 
        .ZN(n10051) );
  MOAI22 U18973 ( .A1(n28438), .A2(n1559), .B1(ram[5811]), .B2(n1560), 
        .ZN(n10052) );
  MOAI22 U18974 ( .A1(n28203), .A2(n1559), .B1(ram[5812]), .B2(n1560), 
        .ZN(n10053) );
  MOAI22 U18975 ( .A1(n27968), .A2(n1559), .B1(ram[5813]), .B2(n1560), 
        .ZN(n10054) );
  MOAI22 U18976 ( .A1(n27733), .A2(n1559), .B1(ram[5814]), .B2(n1560), 
        .ZN(n10055) );
  MOAI22 U18977 ( .A1(n27498), .A2(n1559), .B1(ram[5815]), .B2(n1560), 
        .ZN(n10056) );
  MOAI22 U18978 ( .A1(n29143), .A2(n1561), .B1(ram[5816]), .B2(n1562), 
        .ZN(n10057) );
  MOAI22 U18979 ( .A1(n28908), .A2(n1561), .B1(ram[5817]), .B2(n1562), 
        .ZN(n10058) );
  MOAI22 U18980 ( .A1(n28673), .A2(n1561), .B1(ram[5818]), .B2(n1562), 
        .ZN(n10059) );
  MOAI22 U18981 ( .A1(n28438), .A2(n1561), .B1(ram[5819]), .B2(n1562), 
        .ZN(n10060) );
  MOAI22 U18982 ( .A1(n28203), .A2(n1561), .B1(ram[5820]), .B2(n1562), 
        .ZN(n10061) );
  MOAI22 U18983 ( .A1(n27968), .A2(n1561), .B1(ram[5821]), .B2(n1562), 
        .ZN(n10062) );
  MOAI22 U18984 ( .A1(n27733), .A2(n1561), .B1(ram[5822]), .B2(n1562), 
        .ZN(n10063) );
  MOAI22 U18985 ( .A1(n27498), .A2(n1561), .B1(ram[5823]), .B2(n1562), 
        .ZN(n10064) );
  MOAI22 U18986 ( .A1(n29144), .A2(n1563), .B1(ram[5824]), .B2(n1564), 
        .ZN(n10065) );
  MOAI22 U18987 ( .A1(n28909), .A2(n1563), .B1(ram[5825]), .B2(n1564), 
        .ZN(n10066) );
  MOAI22 U18988 ( .A1(n28674), .A2(n1563), .B1(ram[5826]), .B2(n1564), 
        .ZN(n10067) );
  MOAI22 U18989 ( .A1(n28439), .A2(n1563), .B1(ram[5827]), .B2(n1564), 
        .ZN(n10068) );
  MOAI22 U18990 ( .A1(n28204), .A2(n1563), .B1(ram[5828]), .B2(n1564), 
        .ZN(n10069) );
  MOAI22 U18991 ( .A1(n27969), .A2(n1563), .B1(ram[5829]), .B2(n1564), 
        .ZN(n10070) );
  MOAI22 U18992 ( .A1(n27734), .A2(n1563), .B1(ram[5830]), .B2(n1564), 
        .ZN(n10071) );
  MOAI22 U18993 ( .A1(n27499), .A2(n1563), .B1(ram[5831]), .B2(n1564), 
        .ZN(n10072) );
  MOAI22 U18994 ( .A1(n29144), .A2(n1565), .B1(ram[5832]), .B2(n1566), 
        .ZN(n10073) );
  MOAI22 U18995 ( .A1(n28909), .A2(n1565), .B1(ram[5833]), .B2(n1566), 
        .ZN(n10074) );
  MOAI22 U18996 ( .A1(n28674), .A2(n1565), .B1(ram[5834]), .B2(n1566), 
        .ZN(n10075) );
  MOAI22 U18997 ( .A1(n28439), .A2(n1565), .B1(ram[5835]), .B2(n1566), 
        .ZN(n10076) );
  MOAI22 U18998 ( .A1(n28204), .A2(n1565), .B1(ram[5836]), .B2(n1566), 
        .ZN(n10077) );
  MOAI22 U18999 ( .A1(n27969), .A2(n1565), .B1(ram[5837]), .B2(n1566), 
        .ZN(n10078) );
  MOAI22 U19000 ( .A1(n27734), .A2(n1565), .B1(ram[5838]), .B2(n1566), 
        .ZN(n10079) );
  MOAI22 U19001 ( .A1(n27499), .A2(n1565), .B1(ram[5839]), .B2(n1566), 
        .ZN(n10080) );
  MOAI22 U19002 ( .A1(n29144), .A2(n1567), .B1(ram[5840]), .B2(n1568), 
        .ZN(n10081) );
  MOAI22 U19003 ( .A1(n28909), .A2(n1567), .B1(ram[5841]), .B2(n1568), 
        .ZN(n10082) );
  MOAI22 U19004 ( .A1(n28674), .A2(n1567), .B1(ram[5842]), .B2(n1568), 
        .ZN(n10083) );
  MOAI22 U19005 ( .A1(n28439), .A2(n1567), .B1(ram[5843]), .B2(n1568), 
        .ZN(n10084) );
  MOAI22 U19006 ( .A1(n28204), .A2(n1567), .B1(ram[5844]), .B2(n1568), 
        .ZN(n10085) );
  MOAI22 U19007 ( .A1(n27969), .A2(n1567), .B1(ram[5845]), .B2(n1568), 
        .ZN(n10086) );
  MOAI22 U19008 ( .A1(n27734), .A2(n1567), .B1(ram[5846]), .B2(n1568), 
        .ZN(n10087) );
  MOAI22 U19009 ( .A1(n27499), .A2(n1567), .B1(ram[5847]), .B2(n1568), 
        .ZN(n10088) );
  MOAI22 U19010 ( .A1(n29144), .A2(n1569), .B1(ram[5848]), .B2(n1570), 
        .ZN(n10089) );
  MOAI22 U19011 ( .A1(n28909), .A2(n1569), .B1(ram[5849]), .B2(n1570), 
        .ZN(n10090) );
  MOAI22 U19012 ( .A1(n28674), .A2(n1569), .B1(ram[5850]), .B2(n1570), 
        .ZN(n10091) );
  MOAI22 U19013 ( .A1(n28439), .A2(n1569), .B1(ram[5851]), .B2(n1570), 
        .ZN(n10092) );
  MOAI22 U19014 ( .A1(n28204), .A2(n1569), .B1(ram[5852]), .B2(n1570), 
        .ZN(n10093) );
  MOAI22 U19015 ( .A1(n27969), .A2(n1569), .B1(ram[5853]), .B2(n1570), 
        .ZN(n10094) );
  MOAI22 U19016 ( .A1(n27734), .A2(n1569), .B1(ram[5854]), .B2(n1570), 
        .ZN(n10095) );
  MOAI22 U19017 ( .A1(n27499), .A2(n1569), .B1(ram[5855]), .B2(n1570), 
        .ZN(n10096) );
  MOAI22 U19018 ( .A1(n29144), .A2(n1571), .B1(ram[5856]), .B2(n1572), 
        .ZN(n10097) );
  MOAI22 U19019 ( .A1(n28909), .A2(n1571), .B1(ram[5857]), .B2(n1572), 
        .ZN(n10098) );
  MOAI22 U19020 ( .A1(n28674), .A2(n1571), .B1(ram[5858]), .B2(n1572), 
        .ZN(n10099) );
  MOAI22 U19021 ( .A1(n28439), .A2(n1571), .B1(ram[5859]), .B2(n1572), 
        .ZN(n10100) );
  MOAI22 U19022 ( .A1(n28204), .A2(n1571), .B1(ram[5860]), .B2(n1572), 
        .ZN(n10101) );
  MOAI22 U19023 ( .A1(n27969), .A2(n1571), .B1(ram[5861]), .B2(n1572), 
        .ZN(n10102) );
  MOAI22 U19024 ( .A1(n27734), .A2(n1571), .B1(ram[5862]), .B2(n1572), 
        .ZN(n10103) );
  MOAI22 U19025 ( .A1(n27499), .A2(n1571), .B1(ram[5863]), .B2(n1572), 
        .ZN(n10104) );
  MOAI22 U19026 ( .A1(n29144), .A2(n1573), .B1(ram[5864]), .B2(n1574), 
        .ZN(n10105) );
  MOAI22 U19027 ( .A1(n28909), .A2(n1573), .B1(ram[5865]), .B2(n1574), 
        .ZN(n10106) );
  MOAI22 U19028 ( .A1(n28674), .A2(n1573), .B1(ram[5866]), .B2(n1574), 
        .ZN(n10107) );
  MOAI22 U19029 ( .A1(n28439), .A2(n1573), .B1(ram[5867]), .B2(n1574), 
        .ZN(n10108) );
  MOAI22 U19030 ( .A1(n28204), .A2(n1573), .B1(ram[5868]), .B2(n1574), 
        .ZN(n10109) );
  MOAI22 U19031 ( .A1(n27969), .A2(n1573), .B1(ram[5869]), .B2(n1574), 
        .ZN(n10110) );
  MOAI22 U19032 ( .A1(n27734), .A2(n1573), .B1(ram[5870]), .B2(n1574), 
        .ZN(n10111) );
  MOAI22 U19033 ( .A1(n27499), .A2(n1573), .B1(ram[5871]), .B2(n1574), 
        .ZN(n10112) );
  MOAI22 U19034 ( .A1(n29144), .A2(n1575), .B1(ram[5872]), .B2(n1576), 
        .ZN(n10113) );
  MOAI22 U19035 ( .A1(n28909), .A2(n1575), .B1(ram[5873]), .B2(n1576), 
        .ZN(n10114) );
  MOAI22 U19036 ( .A1(n28674), .A2(n1575), .B1(ram[5874]), .B2(n1576), 
        .ZN(n10115) );
  MOAI22 U19037 ( .A1(n28439), .A2(n1575), .B1(ram[5875]), .B2(n1576), 
        .ZN(n10116) );
  MOAI22 U19038 ( .A1(n28204), .A2(n1575), .B1(ram[5876]), .B2(n1576), 
        .ZN(n10117) );
  MOAI22 U19039 ( .A1(n27969), .A2(n1575), .B1(ram[5877]), .B2(n1576), 
        .ZN(n10118) );
  MOAI22 U19040 ( .A1(n27734), .A2(n1575), .B1(ram[5878]), .B2(n1576), 
        .ZN(n10119) );
  MOAI22 U19041 ( .A1(n27499), .A2(n1575), .B1(ram[5879]), .B2(n1576), 
        .ZN(n10120) );
  MOAI22 U19042 ( .A1(n29144), .A2(n1577), .B1(ram[5880]), .B2(n1578), 
        .ZN(n10121) );
  MOAI22 U19043 ( .A1(n28909), .A2(n1577), .B1(ram[5881]), .B2(n1578), 
        .ZN(n10122) );
  MOAI22 U19044 ( .A1(n28674), .A2(n1577), .B1(ram[5882]), .B2(n1578), 
        .ZN(n10123) );
  MOAI22 U19045 ( .A1(n28439), .A2(n1577), .B1(ram[5883]), .B2(n1578), 
        .ZN(n10124) );
  MOAI22 U19046 ( .A1(n28204), .A2(n1577), .B1(ram[5884]), .B2(n1578), 
        .ZN(n10125) );
  MOAI22 U19047 ( .A1(n27969), .A2(n1577), .B1(ram[5885]), .B2(n1578), 
        .ZN(n10126) );
  MOAI22 U19048 ( .A1(n27734), .A2(n1577), .B1(ram[5886]), .B2(n1578), 
        .ZN(n10127) );
  MOAI22 U19049 ( .A1(n27499), .A2(n1577), .B1(ram[5887]), .B2(n1578), 
        .ZN(n10128) );
  MOAI22 U19050 ( .A1(n29144), .A2(n1579), .B1(ram[5888]), .B2(n1580), 
        .ZN(n10129) );
  MOAI22 U19051 ( .A1(n28909), .A2(n1579), .B1(ram[5889]), .B2(n1580), 
        .ZN(n10130) );
  MOAI22 U19052 ( .A1(n28674), .A2(n1579), .B1(ram[5890]), .B2(n1580), 
        .ZN(n10131) );
  MOAI22 U19053 ( .A1(n28439), .A2(n1579), .B1(ram[5891]), .B2(n1580), 
        .ZN(n10132) );
  MOAI22 U19054 ( .A1(n28204), .A2(n1579), .B1(ram[5892]), .B2(n1580), 
        .ZN(n10133) );
  MOAI22 U19055 ( .A1(n27969), .A2(n1579), .B1(ram[5893]), .B2(n1580), 
        .ZN(n10134) );
  MOAI22 U19056 ( .A1(n27734), .A2(n1579), .B1(ram[5894]), .B2(n1580), 
        .ZN(n10135) );
  MOAI22 U19057 ( .A1(n27499), .A2(n1579), .B1(ram[5895]), .B2(n1580), 
        .ZN(n10136) );
  MOAI22 U19058 ( .A1(n29144), .A2(n1581), .B1(ram[5896]), .B2(n1582), 
        .ZN(n10137) );
  MOAI22 U19059 ( .A1(n28909), .A2(n1581), .B1(ram[5897]), .B2(n1582), 
        .ZN(n10138) );
  MOAI22 U19060 ( .A1(n28674), .A2(n1581), .B1(ram[5898]), .B2(n1582), 
        .ZN(n10139) );
  MOAI22 U19061 ( .A1(n28439), .A2(n1581), .B1(ram[5899]), .B2(n1582), 
        .ZN(n10140) );
  MOAI22 U19062 ( .A1(n28204), .A2(n1581), .B1(ram[5900]), .B2(n1582), 
        .ZN(n10141) );
  MOAI22 U19063 ( .A1(n27969), .A2(n1581), .B1(ram[5901]), .B2(n1582), 
        .ZN(n10142) );
  MOAI22 U19064 ( .A1(n27734), .A2(n1581), .B1(ram[5902]), .B2(n1582), 
        .ZN(n10143) );
  MOAI22 U19065 ( .A1(n27499), .A2(n1581), .B1(ram[5903]), .B2(n1582), 
        .ZN(n10144) );
  MOAI22 U19066 ( .A1(n29144), .A2(n1583), .B1(ram[5904]), .B2(n1584), 
        .ZN(n10145) );
  MOAI22 U19067 ( .A1(n28909), .A2(n1583), .B1(ram[5905]), .B2(n1584), 
        .ZN(n10146) );
  MOAI22 U19068 ( .A1(n28674), .A2(n1583), .B1(ram[5906]), .B2(n1584), 
        .ZN(n10147) );
  MOAI22 U19069 ( .A1(n28439), .A2(n1583), .B1(ram[5907]), .B2(n1584), 
        .ZN(n10148) );
  MOAI22 U19070 ( .A1(n28204), .A2(n1583), .B1(ram[5908]), .B2(n1584), 
        .ZN(n10149) );
  MOAI22 U19071 ( .A1(n27969), .A2(n1583), .B1(ram[5909]), .B2(n1584), 
        .ZN(n10150) );
  MOAI22 U19072 ( .A1(n27734), .A2(n1583), .B1(ram[5910]), .B2(n1584), 
        .ZN(n10151) );
  MOAI22 U19073 ( .A1(n27499), .A2(n1583), .B1(ram[5911]), .B2(n1584), 
        .ZN(n10152) );
  MOAI22 U19074 ( .A1(n29144), .A2(n1585), .B1(ram[5912]), .B2(n1586), 
        .ZN(n10153) );
  MOAI22 U19075 ( .A1(n28909), .A2(n1585), .B1(ram[5913]), .B2(n1586), 
        .ZN(n10154) );
  MOAI22 U19076 ( .A1(n28674), .A2(n1585), .B1(ram[5914]), .B2(n1586), 
        .ZN(n10155) );
  MOAI22 U19077 ( .A1(n28439), .A2(n1585), .B1(ram[5915]), .B2(n1586), 
        .ZN(n10156) );
  MOAI22 U19078 ( .A1(n28204), .A2(n1585), .B1(ram[5916]), .B2(n1586), 
        .ZN(n10157) );
  MOAI22 U19079 ( .A1(n27969), .A2(n1585), .B1(ram[5917]), .B2(n1586), 
        .ZN(n10158) );
  MOAI22 U19080 ( .A1(n27734), .A2(n1585), .B1(ram[5918]), .B2(n1586), 
        .ZN(n10159) );
  MOAI22 U19081 ( .A1(n27499), .A2(n1585), .B1(ram[5919]), .B2(n1586), 
        .ZN(n10160) );
  MOAI22 U19082 ( .A1(n29144), .A2(n1587), .B1(ram[5920]), .B2(n1588), 
        .ZN(n10161) );
  MOAI22 U19083 ( .A1(n28909), .A2(n1587), .B1(ram[5921]), .B2(n1588), 
        .ZN(n10162) );
  MOAI22 U19084 ( .A1(n28674), .A2(n1587), .B1(ram[5922]), .B2(n1588), 
        .ZN(n10163) );
  MOAI22 U19085 ( .A1(n28439), .A2(n1587), .B1(ram[5923]), .B2(n1588), 
        .ZN(n10164) );
  MOAI22 U19086 ( .A1(n28204), .A2(n1587), .B1(ram[5924]), .B2(n1588), 
        .ZN(n10165) );
  MOAI22 U19087 ( .A1(n27969), .A2(n1587), .B1(ram[5925]), .B2(n1588), 
        .ZN(n10166) );
  MOAI22 U19088 ( .A1(n27734), .A2(n1587), .B1(ram[5926]), .B2(n1588), 
        .ZN(n10167) );
  MOAI22 U19089 ( .A1(n27499), .A2(n1587), .B1(ram[5927]), .B2(n1588), 
        .ZN(n10168) );
  MOAI22 U19090 ( .A1(n29145), .A2(n1589), .B1(ram[5928]), .B2(n1590), 
        .ZN(n10169) );
  MOAI22 U19091 ( .A1(n28910), .A2(n1589), .B1(ram[5929]), .B2(n1590), 
        .ZN(n10170) );
  MOAI22 U19092 ( .A1(n28675), .A2(n1589), .B1(ram[5930]), .B2(n1590), 
        .ZN(n10171) );
  MOAI22 U19093 ( .A1(n28440), .A2(n1589), .B1(ram[5931]), .B2(n1590), 
        .ZN(n10172) );
  MOAI22 U19094 ( .A1(n28205), .A2(n1589), .B1(ram[5932]), .B2(n1590), 
        .ZN(n10173) );
  MOAI22 U19095 ( .A1(n27970), .A2(n1589), .B1(ram[5933]), .B2(n1590), 
        .ZN(n10174) );
  MOAI22 U19096 ( .A1(n27735), .A2(n1589), .B1(ram[5934]), .B2(n1590), 
        .ZN(n10175) );
  MOAI22 U19097 ( .A1(n27500), .A2(n1589), .B1(ram[5935]), .B2(n1590), 
        .ZN(n10176) );
  MOAI22 U19098 ( .A1(n29145), .A2(n1591), .B1(ram[5936]), .B2(n1592), 
        .ZN(n10177) );
  MOAI22 U19099 ( .A1(n28910), .A2(n1591), .B1(ram[5937]), .B2(n1592), 
        .ZN(n10178) );
  MOAI22 U19100 ( .A1(n28675), .A2(n1591), .B1(ram[5938]), .B2(n1592), 
        .ZN(n10179) );
  MOAI22 U19101 ( .A1(n28440), .A2(n1591), .B1(ram[5939]), .B2(n1592), 
        .ZN(n10180) );
  MOAI22 U19102 ( .A1(n28205), .A2(n1591), .B1(ram[5940]), .B2(n1592), 
        .ZN(n10181) );
  MOAI22 U19103 ( .A1(n27970), .A2(n1591), .B1(ram[5941]), .B2(n1592), 
        .ZN(n10182) );
  MOAI22 U19104 ( .A1(n27735), .A2(n1591), .B1(ram[5942]), .B2(n1592), 
        .ZN(n10183) );
  MOAI22 U19105 ( .A1(n27500), .A2(n1591), .B1(ram[5943]), .B2(n1592), 
        .ZN(n10184) );
  MOAI22 U19106 ( .A1(n29145), .A2(n1593), .B1(ram[5944]), .B2(n1594), 
        .ZN(n10185) );
  MOAI22 U19107 ( .A1(n28910), .A2(n1593), .B1(ram[5945]), .B2(n1594), 
        .ZN(n10186) );
  MOAI22 U19108 ( .A1(n28675), .A2(n1593), .B1(ram[5946]), .B2(n1594), 
        .ZN(n10187) );
  MOAI22 U19109 ( .A1(n28440), .A2(n1593), .B1(ram[5947]), .B2(n1594), 
        .ZN(n10188) );
  MOAI22 U19110 ( .A1(n28205), .A2(n1593), .B1(ram[5948]), .B2(n1594), 
        .ZN(n10189) );
  MOAI22 U19111 ( .A1(n27970), .A2(n1593), .B1(ram[5949]), .B2(n1594), 
        .ZN(n10190) );
  MOAI22 U19112 ( .A1(n27735), .A2(n1593), .B1(ram[5950]), .B2(n1594), 
        .ZN(n10191) );
  MOAI22 U19113 ( .A1(n27500), .A2(n1593), .B1(ram[5951]), .B2(n1594), 
        .ZN(n10192) );
  MOAI22 U19114 ( .A1(n29145), .A2(n1595), .B1(ram[5952]), .B2(n1596), 
        .ZN(n10193) );
  MOAI22 U19115 ( .A1(n28910), .A2(n1595), .B1(ram[5953]), .B2(n1596), 
        .ZN(n10194) );
  MOAI22 U19116 ( .A1(n28675), .A2(n1595), .B1(ram[5954]), .B2(n1596), 
        .ZN(n10195) );
  MOAI22 U19117 ( .A1(n28440), .A2(n1595), .B1(ram[5955]), .B2(n1596), 
        .ZN(n10196) );
  MOAI22 U19118 ( .A1(n28205), .A2(n1595), .B1(ram[5956]), .B2(n1596), 
        .ZN(n10197) );
  MOAI22 U19119 ( .A1(n27970), .A2(n1595), .B1(ram[5957]), .B2(n1596), 
        .ZN(n10198) );
  MOAI22 U19120 ( .A1(n27735), .A2(n1595), .B1(ram[5958]), .B2(n1596), 
        .ZN(n10199) );
  MOAI22 U19121 ( .A1(n27500), .A2(n1595), .B1(ram[5959]), .B2(n1596), 
        .ZN(n10200) );
  MOAI22 U19122 ( .A1(n29145), .A2(n1597), .B1(ram[5960]), .B2(n1598), 
        .ZN(n10201) );
  MOAI22 U19123 ( .A1(n28910), .A2(n1597), .B1(ram[5961]), .B2(n1598), 
        .ZN(n10202) );
  MOAI22 U19124 ( .A1(n28675), .A2(n1597), .B1(ram[5962]), .B2(n1598), 
        .ZN(n10203) );
  MOAI22 U19125 ( .A1(n28440), .A2(n1597), .B1(ram[5963]), .B2(n1598), 
        .ZN(n10204) );
  MOAI22 U19126 ( .A1(n28205), .A2(n1597), .B1(ram[5964]), .B2(n1598), 
        .ZN(n10205) );
  MOAI22 U19127 ( .A1(n27970), .A2(n1597), .B1(ram[5965]), .B2(n1598), 
        .ZN(n10206) );
  MOAI22 U19128 ( .A1(n27735), .A2(n1597), .B1(ram[5966]), .B2(n1598), 
        .ZN(n10207) );
  MOAI22 U19129 ( .A1(n27500), .A2(n1597), .B1(ram[5967]), .B2(n1598), 
        .ZN(n10208) );
  MOAI22 U19130 ( .A1(n29145), .A2(n1599), .B1(ram[5968]), .B2(n1600), 
        .ZN(n10209) );
  MOAI22 U19131 ( .A1(n28910), .A2(n1599), .B1(ram[5969]), .B2(n1600), 
        .ZN(n10210) );
  MOAI22 U19132 ( .A1(n28675), .A2(n1599), .B1(ram[5970]), .B2(n1600), 
        .ZN(n10211) );
  MOAI22 U19133 ( .A1(n28440), .A2(n1599), .B1(ram[5971]), .B2(n1600), 
        .ZN(n10212) );
  MOAI22 U19134 ( .A1(n28205), .A2(n1599), .B1(ram[5972]), .B2(n1600), 
        .ZN(n10213) );
  MOAI22 U19135 ( .A1(n27970), .A2(n1599), .B1(ram[5973]), .B2(n1600), 
        .ZN(n10214) );
  MOAI22 U19136 ( .A1(n27735), .A2(n1599), .B1(ram[5974]), .B2(n1600), 
        .ZN(n10215) );
  MOAI22 U19137 ( .A1(n27500), .A2(n1599), .B1(ram[5975]), .B2(n1600), 
        .ZN(n10216) );
  MOAI22 U19138 ( .A1(n29145), .A2(n1601), .B1(ram[5976]), .B2(n1602), 
        .ZN(n10217) );
  MOAI22 U19139 ( .A1(n28910), .A2(n1601), .B1(ram[5977]), .B2(n1602), 
        .ZN(n10218) );
  MOAI22 U19140 ( .A1(n28675), .A2(n1601), .B1(ram[5978]), .B2(n1602), 
        .ZN(n10219) );
  MOAI22 U19141 ( .A1(n28440), .A2(n1601), .B1(ram[5979]), .B2(n1602), 
        .ZN(n10220) );
  MOAI22 U19142 ( .A1(n28205), .A2(n1601), .B1(ram[5980]), .B2(n1602), 
        .ZN(n10221) );
  MOAI22 U19143 ( .A1(n27970), .A2(n1601), .B1(ram[5981]), .B2(n1602), 
        .ZN(n10222) );
  MOAI22 U19144 ( .A1(n27735), .A2(n1601), .B1(ram[5982]), .B2(n1602), 
        .ZN(n10223) );
  MOAI22 U19145 ( .A1(n27500), .A2(n1601), .B1(ram[5983]), .B2(n1602), 
        .ZN(n10224) );
  MOAI22 U19146 ( .A1(n29145), .A2(n1603), .B1(ram[5984]), .B2(n1604), 
        .ZN(n10225) );
  MOAI22 U19147 ( .A1(n28910), .A2(n1603), .B1(ram[5985]), .B2(n1604), 
        .ZN(n10226) );
  MOAI22 U19148 ( .A1(n28675), .A2(n1603), .B1(ram[5986]), .B2(n1604), 
        .ZN(n10227) );
  MOAI22 U19149 ( .A1(n28440), .A2(n1603), .B1(ram[5987]), .B2(n1604), 
        .ZN(n10228) );
  MOAI22 U19150 ( .A1(n28205), .A2(n1603), .B1(ram[5988]), .B2(n1604), 
        .ZN(n10229) );
  MOAI22 U19151 ( .A1(n27970), .A2(n1603), .B1(ram[5989]), .B2(n1604), 
        .ZN(n10230) );
  MOAI22 U19152 ( .A1(n27735), .A2(n1603), .B1(ram[5990]), .B2(n1604), 
        .ZN(n10231) );
  MOAI22 U19153 ( .A1(n27500), .A2(n1603), .B1(ram[5991]), .B2(n1604), 
        .ZN(n10232) );
  MOAI22 U19154 ( .A1(n29145), .A2(n1605), .B1(ram[5992]), .B2(n1606), 
        .ZN(n10233) );
  MOAI22 U19155 ( .A1(n28910), .A2(n1605), .B1(ram[5993]), .B2(n1606), 
        .ZN(n10234) );
  MOAI22 U19156 ( .A1(n28675), .A2(n1605), .B1(ram[5994]), .B2(n1606), 
        .ZN(n10235) );
  MOAI22 U19157 ( .A1(n28440), .A2(n1605), .B1(ram[5995]), .B2(n1606), 
        .ZN(n10236) );
  MOAI22 U19158 ( .A1(n28205), .A2(n1605), .B1(ram[5996]), .B2(n1606), 
        .ZN(n10237) );
  MOAI22 U19159 ( .A1(n27970), .A2(n1605), .B1(ram[5997]), .B2(n1606), 
        .ZN(n10238) );
  MOAI22 U19160 ( .A1(n27735), .A2(n1605), .B1(ram[5998]), .B2(n1606), 
        .ZN(n10239) );
  MOAI22 U19161 ( .A1(n27500), .A2(n1605), .B1(ram[5999]), .B2(n1606), 
        .ZN(n10240) );
  MOAI22 U19162 ( .A1(n29145), .A2(n1607), .B1(ram[6000]), .B2(n1608), 
        .ZN(n10241) );
  MOAI22 U19163 ( .A1(n28910), .A2(n1607), .B1(ram[6001]), .B2(n1608), 
        .ZN(n10242) );
  MOAI22 U19164 ( .A1(n28675), .A2(n1607), .B1(ram[6002]), .B2(n1608), 
        .ZN(n10243) );
  MOAI22 U19165 ( .A1(n28440), .A2(n1607), .B1(ram[6003]), .B2(n1608), 
        .ZN(n10244) );
  MOAI22 U19166 ( .A1(n28205), .A2(n1607), .B1(ram[6004]), .B2(n1608), 
        .ZN(n10245) );
  MOAI22 U19167 ( .A1(n27970), .A2(n1607), .B1(ram[6005]), .B2(n1608), 
        .ZN(n10246) );
  MOAI22 U19168 ( .A1(n27735), .A2(n1607), .B1(ram[6006]), .B2(n1608), 
        .ZN(n10247) );
  MOAI22 U19169 ( .A1(n27500), .A2(n1607), .B1(ram[6007]), .B2(n1608), 
        .ZN(n10248) );
  MOAI22 U19170 ( .A1(n29145), .A2(n1609), .B1(ram[6008]), .B2(n1610), 
        .ZN(n10249) );
  MOAI22 U19171 ( .A1(n28910), .A2(n1609), .B1(ram[6009]), .B2(n1610), 
        .ZN(n10250) );
  MOAI22 U19172 ( .A1(n28675), .A2(n1609), .B1(ram[6010]), .B2(n1610), 
        .ZN(n10251) );
  MOAI22 U19173 ( .A1(n28440), .A2(n1609), .B1(ram[6011]), .B2(n1610), 
        .ZN(n10252) );
  MOAI22 U19174 ( .A1(n28205), .A2(n1609), .B1(ram[6012]), .B2(n1610), 
        .ZN(n10253) );
  MOAI22 U19175 ( .A1(n27970), .A2(n1609), .B1(ram[6013]), .B2(n1610), 
        .ZN(n10254) );
  MOAI22 U19176 ( .A1(n27735), .A2(n1609), .B1(ram[6014]), .B2(n1610), 
        .ZN(n10255) );
  MOAI22 U19177 ( .A1(n27500), .A2(n1609), .B1(ram[6015]), .B2(n1610), 
        .ZN(n10256) );
  MOAI22 U19178 ( .A1(n29145), .A2(n1611), .B1(ram[6016]), .B2(n1612), 
        .ZN(n10257) );
  MOAI22 U19179 ( .A1(n28910), .A2(n1611), .B1(ram[6017]), .B2(n1612), 
        .ZN(n10258) );
  MOAI22 U19180 ( .A1(n28675), .A2(n1611), .B1(ram[6018]), .B2(n1612), 
        .ZN(n10259) );
  MOAI22 U19181 ( .A1(n28440), .A2(n1611), .B1(ram[6019]), .B2(n1612), 
        .ZN(n10260) );
  MOAI22 U19182 ( .A1(n28205), .A2(n1611), .B1(ram[6020]), .B2(n1612), 
        .ZN(n10261) );
  MOAI22 U19183 ( .A1(n27970), .A2(n1611), .B1(ram[6021]), .B2(n1612), 
        .ZN(n10262) );
  MOAI22 U19184 ( .A1(n27735), .A2(n1611), .B1(ram[6022]), .B2(n1612), 
        .ZN(n10263) );
  MOAI22 U19185 ( .A1(n27500), .A2(n1611), .B1(ram[6023]), .B2(n1612), 
        .ZN(n10264) );
  MOAI22 U19186 ( .A1(n29145), .A2(n1613), .B1(ram[6024]), .B2(n1614), 
        .ZN(n10265) );
  MOAI22 U19187 ( .A1(n28910), .A2(n1613), .B1(ram[6025]), .B2(n1614), 
        .ZN(n10266) );
  MOAI22 U19188 ( .A1(n28675), .A2(n1613), .B1(ram[6026]), .B2(n1614), 
        .ZN(n10267) );
  MOAI22 U19189 ( .A1(n28440), .A2(n1613), .B1(ram[6027]), .B2(n1614), 
        .ZN(n10268) );
  MOAI22 U19190 ( .A1(n28205), .A2(n1613), .B1(ram[6028]), .B2(n1614), 
        .ZN(n10269) );
  MOAI22 U19191 ( .A1(n27970), .A2(n1613), .B1(ram[6029]), .B2(n1614), 
        .ZN(n10270) );
  MOAI22 U19192 ( .A1(n27735), .A2(n1613), .B1(ram[6030]), .B2(n1614), 
        .ZN(n10271) );
  MOAI22 U19193 ( .A1(n27500), .A2(n1613), .B1(ram[6031]), .B2(n1614), 
        .ZN(n10272) );
  MOAI22 U19194 ( .A1(n29146), .A2(n1615), .B1(ram[6032]), .B2(n1616), 
        .ZN(n10273) );
  MOAI22 U19195 ( .A1(n28911), .A2(n1615), .B1(ram[6033]), .B2(n1616), 
        .ZN(n10274) );
  MOAI22 U19196 ( .A1(n28676), .A2(n1615), .B1(ram[6034]), .B2(n1616), 
        .ZN(n10275) );
  MOAI22 U19197 ( .A1(n28441), .A2(n1615), .B1(ram[6035]), .B2(n1616), 
        .ZN(n10276) );
  MOAI22 U19198 ( .A1(n28206), .A2(n1615), .B1(ram[6036]), .B2(n1616), 
        .ZN(n10277) );
  MOAI22 U19199 ( .A1(n27971), .A2(n1615), .B1(ram[6037]), .B2(n1616), 
        .ZN(n10278) );
  MOAI22 U19200 ( .A1(n27736), .A2(n1615), .B1(ram[6038]), .B2(n1616), 
        .ZN(n10279) );
  MOAI22 U19201 ( .A1(n27501), .A2(n1615), .B1(ram[6039]), .B2(n1616), 
        .ZN(n10280) );
  MOAI22 U19202 ( .A1(n29146), .A2(n1617), .B1(ram[6040]), .B2(n1618), 
        .ZN(n10281) );
  MOAI22 U19203 ( .A1(n28911), .A2(n1617), .B1(ram[6041]), .B2(n1618), 
        .ZN(n10282) );
  MOAI22 U19204 ( .A1(n28676), .A2(n1617), .B1(ram[6042]), .B2(n1618), 
        .ZN(n10283) );
  MOAI22 U19205 ( .A1(n28441), .A2(n1617), .B1(ram[6043]), .B2(n1618), 
        .ZN(n10284) );
  MOAI22 U19206 ( .A1(n28206), .A2(n1617), .B1(ram[6044]), .B2(n1618), 
        .ZN(n10285) );
  MOAI22 U19207 ( .A1(n27971), .A2(n1617), .B1(ram[6045]), .B2(n1618), 
        .ZN(n10286) );
  MOAI22 U19208 ( .A1(n27736), .A2(n1617), .B1(ram[6046]), .B2(n1618), 
        .ZN(n10287) );
  MOAI22 U19209 ( .A1(n27501), .A2(n1617), .B1(ram[6047]), .B2(n1618), 
        .ZN(n10288) );
  MOAI22 U19210 ( .A1(n29146), .A2(n1619), .B1(ram[6048]), .B2(n1620), 
        .ZN(n10289) );
  MOAI22 U19211 ( .A1(n28911), .A2(n1619), .B1(ram[6049]), .B2(n1620), 
        .ZN(n10290) );
  MOAI22 U19212 ( .A1(n28676), .A2(n1619), .B1(ram[6050]), .B2(n1620), 
        .ZN(n10291) );
  MOAI22 U19213 ( .A1(n28441), .A2(n1619), .B1(ram[6051]), .B2(n1620), 
        .ZN(n10292) );
  MOAI22 U19214 ( .A1(n28206), .A2(n1619), .B1(ram[6052]), .B2(n1620), 
        .ZN(n10293) );
  MOAI22 U19215 ( .A1(n27971), .A2(n1619), .B1(ram[6053]), .B2(n1620), 
        .ZN(n10294) );
  MOAI22 U19216 ( .A1(n27736), .A2(n1619), .B1(ram[6054]), .B2(n1620), 
        .ZN(n10295) );
  MOAI22 U19217 ( .A1(n27501), .A2(n1619), .B1(ram[6055]), .B2(n1620), 
        .ZN(n10296) );
  MOAI22 U19218 ( .A1(n29146), .A2(n1621), .B1(ram[6056]), .B2(n1622), 
        .ZN(n10297) );
  MOAI22 U19219 ( .A1(n28911), .A2(n1621), .B1(ram[6057]), .B2(n1622), 
        .ZN(n10298) );
  MOAI22 U19220 ( .A1(n28676), .A2(n1621), .B1(ram[6058]), .B2(n1622), 
        .ZN(n10299) );
  MOAI22 U19221 ( .A1(n28441), .A2(n1621), .B1(ram[6059]), .B2(n1622), 
        .ZN(n10300) );
  MOAI22 U19222 ( .A1(n28206), .A2(n1621), .B1(ram[6060]), .B2(n1622), 
        .ZN(n10301) );
  MOAI22 U19223 ( .A1(n27971), .A2(n1621), .B1(ram[6061]), .B2(n1622), 
        .ZN(n10302) );
  MOAI22 U19224 ( .A1(n27736), .A2(n1621), .B1(ram[6062]), .B2(n1622), 
        .ZN(n10303) );
  MOAI22 U19225 ( .A1(n27501), .A2(n1621), .B1(ram[6063]), .B2(n1622), 
        .ZN(n10304) );
  MOAI22 U19226 ( .A1(n29146), .A2(n1623), .B1(ram[6064]), .B2(n1624), 
        .ZN(n10305) );
  MOAI22 U19227 ( .A1(n28911), .A2(n1623), .B1(ram[6065]), .B2(n1624), 
        .ZN(n10306) );
  MOAI22 U19228 ( .A1(n28676), .A2(n1623), .B1(ram[6066]), .B2(n1624), 
        .ZN(n10307) );
  MOAI22 U19229 ( .A1(n28441), .A2(n1623), .B1(ram[6067]), .B2(n1624), 
        .ZN(n10308) );
  MOAI22 U19230 ( .A1(n28206), .A2(n1623), .B1(ram[6068]), .B2(n1624), 
        .ZN(n10309) );
  MOAI22 U19231 ( .A1(n27971), .A2(n1623), .B1(ram[6069]), .B2(n1624), 
        .ZN(n10310) );
  MOAI22 U19232 ( .A1(n27736), .A2(n1623), .B1(ram[6070]), .B2(n1624), 
        .ZN(n10311) );
  MOAI22 U19233 ( .A1(n27501), .A2(n1623), .B1(ram[6071]), .B2(n1624), 
        .ZN(n10312) );
  MOAI22 U19234 ( .A1(n29146), .A2(n1625), .B1(ram[6072]), .B2(n1626), 
        .ZN(n10313) );
  MOAI22 U19235 ( .A1(n28911), .A2(n1625), .B1(ram[6073]), .B2(n1626), 
        .ZN(n10314) );
  MOAI22 U19236 ( .A1(n28676), .A2(n1625), .B1(ram[6074]), .B2(n1626), 
        .ZN(n10315) );
  MOAI22 U19237 ( .A1(n28441), .A2(n1625), .B1(ram[6075]), .B2(n1626), 
        .ZN(n10316) );
  MOAI22 U19238 ( .A1(n28206), .A2(n1625), .B1(ram[6076]), .B2(n1626), 
        .ZN(n10317) );
  MOAI22 U19239 ( .A1(n27971), .A2(n1625), .B1(ram[6077]), .B2(n1626), 
        .ZN(n10318) );
  MOAI22 U19240 ( .A1(n27736), .A2(n1625), .B1(ram[6078]), .B2(n1626), 
        .ZN(n10319) );
  MOAI22 U19241 ( .A1(n27501), .A2(n1625), .B1(ram[6079]), .B2(n1626), 
        .ZN(n10320) );
  MOAI22 U19242 ( .A1(n29146), .A2(n1627), .B1(ram[6080]), .B2(n1628), 
        .ZN(n10321) );
  MOAI22 U19243 ( .A1(n28911), .A2(n1627), .B1(ram[6081]), .B2(n1628), 
        .ZN(n10322) );
  MOAI22 U19244 ( .A1(n28676), .A2(n1627), .B1(ram[6082]), .B2(n1628), 
        .ZN(n10323) );
  MOAI22 U19245 ( .A1(n28441), .A2(n1627), .B1(ram[6083]), .B2(n1628), 
        .ZN(n10324) );
  MOAI22 U19246 ( .A1(n28206), .A2(n1627), .B1(ram[6084]), .B2(n1628), 
        .ZN(n10325) );
  MOAI22 U19247 ( .A1(n27971), .A2(n1627), .B1(ram[6085]), .B2(n1628), 
        .ZN(n10326) );
  MOAI22 U19248 ( .A1(n27736), .A2(n1627), .B1(ram[6086]), .B2(n1628), 
        .ZN(n10327) );
  MOAI22 U19249 ( .A1(n27501), .A2(n1627), .B1(ram[6087]), .B2(n1628), 
        .ZN(n10328) );
  MOAI22 U19250 ( .A1(n29146), .A2(n1629), .B1(ram[6088]), .B2(n1630), 
        .ZN(n10329) );
  MOAI22 U19251 ( .A1(n28911), .A2(n1629), .B1(ram[6089]), .B2(n1630), 
        .ZN(n10330) );
  MOAI22 U19252 ( .A1(n28676), .A2(n1629), .B1(ram[6090]), .B2(n1630), 
        .ZN(n10331) );
  MOAI22 U19253 ( .A1(n28441), .A2(n1629), .B1(ram[6091]), .B2(n1630), 
        .ZN(n10332) );
  MOAI22 U19254 ( .A1(n28206), .A2(n1629), .B1(ram[6092]), .B2(n1630), 
        .ZN(n10333) );
  MOAI22 U19255 ( .A1(n27971), .A2(n1629), .B1(ram[6093]), .B2(n1630), 
        .ZN(n10334) );
  MOAI22 U19256 ( .A1(n27736), .A2(n1629), .B1(ram[6094]), .B2(n1630), 
        .ZN(n10335) );
  MOAI22 U19257 ( .A1(n27501), .A2(n1629), .B1(ram[6095]), .B2(n1630), 
        .ZN(n10336) );
  MOAI22 U19258 ( .A1(n29146), .A2(n1631), .B1(ram[6096]), .B2(n1632), 
        .ZN(n10337) );
  MOAI22 U19259 ( .A1(n28911), .A2(n1631), .B1(ram[6097]), .B2(n1632), 
        .ZN(n10338) );
  MOAI22 U19260 ( .A1(n28676), .A2(n1631), .B1(ram[6098]), .B2(n1632), 
        .ZN(n10339) );
  MOAI22 U19261 ( .A1(n28441), .A2(n1631), .B1(ram[6099]), .B2(n1632), 
        .ZN(n10340) );
  MOAI22 U19262 ( .A1(n28206), .A2(n1631), .B1(ram[6100]), .B2(n1632), 
        .ZN(n10341) );
  MOAI22 U19263 ( .A1(n27971), .A2(n1631), .B1(ram[6101]), .B2(n1632), 
        .ZN(n10342) );
  MOAI22 U19264 ( .A1(n27736), .A2(n1631), .B1(ram[6102]), .B2(n1632), 
        .ZN(n10343) );
  MOAI22 U19265 ( .A1(n27501), .A2(n1631), .B1(ram[6103]), .B2(n1632), 
        .ZN(n10344) );
  MOAI22 U19266 ( .A1(n29146), .A2(n1633), .B1(ram[6104]), .B2(n1634), 
        .ZN(n10345) );
  MOAI22 U19267 ( .A1(n28911), .A2(n1633), .B1(ram[6105]), .B2(n1634), 
        .ZN(n10346) );
  MOAI22 U19268 ( .A1(n28676), .A2(n1633), .B1(ram[6106]), .B2(n1634), 
        .ZN(n10347) );
  MOAI22 U19269 ( .A1(n28441), .A2(n1633), .B1(ram[6107]), .B2(n1634), 
        .ZN(n10348) );
  MOAI22 U19270 ( .A1(n28206), .A2(n1633), .B1(ram[6108]), .B2(n1634), 
        .ZN(n10349) );
  MOAI22 U19271 ( .A1(n27971), .A2(n1633), .B1(ram[6109]), .B2(n1634), 
        .ZN(n10350) );
  MOAI22 U19272 ( .A1(n27736), .A2(n1633), .B1(ram[6110]), .B2(n1634), 
        .ZN(n10351) );
  MOAI22 U19273 ( .A1(n27501), .A2(n1633), .B1(ram[6111]), .B2(n1634), 
        .ZN(n10352) );
  MOAI22 U19274 ( .A1(n29146), .A2(n1635), .B1(ram[6112]), .B2(n1636), 
        .ZN(n10353) );
  MOAI22 U19275 ( .A1(n28911), .A2(n1635), .B1(ram[6113]), .B2(n1636), 
        .ZN(n10354) );
  MOAI22 U19276 ( .A1(n28676), .A2(n1635), .B1(ram[6114]), .B2(n1636), 
        .ZN(n10355) );
  MOAI22 U19277 ( .A1(n28441), .A2(n1635), .B1(ram[6115]), .B2(n1636), 
        .ZN(n10356) );
  MOAI22 U19278 ( .A1(n28206), .A2(n1635), .B1(ram[6116]), .B2(n1636), 
        .ZN(n10357) );
  MOAI22 U19279 ( .A1(n27971), .A2(n1635), .B1(ram[6117]), .B2(n1636), 
        .ZN(n10358) );
  MOAI22 U19280 ( .A1(n27736), .A2(n1635), .B1(ram[6118]), .B2(n1636), 
        .ZN(n10359) );
  MOAI22 U19281 ( .A1(n27501), .A2(n1635), .B1(ram[6119]), .B2(n1636), 
        .ZN(n10360) );
  MOAI22 U19282 ( .A1(n29146), .A2(n1637), .B1(ram[6120]), .B2(n1638), 
        .ZN(n10361) );
  MOAI22 U19283 ( .A1(n28911), .A2(n1637), .B1(ram[6121]), .B2(n1638), 
        .ZN(n10362) );
  MOAI22 U19284 ( .A1(n28676), .A2(n1637), .B1(ram[6122]), .B2(n1638), 
        .ZN(n10363) );
  MOAI22 U19285 ( .A1(n28441), .A2(n1637), .B1(ram[6123]), .B2(n1638), 
        .ZN(n10364) );
  MOAI22 U19286 ( .A1(n28206), .A2(n1637), .B1(ram[6124]), .B2(n1638), 
        .ZN(n10365) );
  MOAI22 U19287 ( .A1(n27971), .A2(n1637), .B1(ram[6125]), .B2(n1638), 
        .ZN(n10366) );
  MOAI22 U19288 ( .A1(n27736), .A2(n1637), .B1(ram[6126]), .B2(n1638), 
        .ZN(n10367) );
  MOAI22 U19289 ( .A1(n27501), .A2(n1637), .B1(ram[6127]), .B2(n1638), 
        .ZN(n10368) );
  MOAI22 U19290 ( .A1(n29146), .A2(n1639), .B1(ram[6128]), .B2(n1640), 
        .ZN(n10369) );
  MOAI22 U19291 ( .A1(n28911), .A2(n1639), .B1(ram[6129]), .B2(n1640), 
        .ZN(n10370) );
  MOAI22 U19292 ( .A1(n28676), .A2(n1639), .B1(ram[6130]), .B2(n1640), 
        .ZN(n10371) );
  MOAI22 U19293 ( .A1(n28441), .A2(n1639), .B1(ram[6131]), .B2(n1640), 
        .ZN(n10372) );
  MOAI22 U19294 ( .A1(n28206), .A2(n1639), .B1(ram[6132]), .B2(n1640), 
        .ZN(n10373) );
  MOAI22 U19295 ( .A1(n27971), .A2(n1639), .B1(ram[6133]), .B2(n1640), 
        .ZN(n10374) );
  MOAI22 U19296 ( .A1(n27736), .A2(n1639), .B1(ram[6134]), .B2(n1640), 
        .ZN(n10375) );
  MOAI22 U19297 ( .A1(n27501), .A2(n1639), .B1(ram[6135]), .B2(n1640), 
        .ZN(n10376) );
  MOAI22 U19298 ( .A1(n29147), .A2(n1641), .B1(ram[6136]), .B2(n1642), 
        .ZN(n10377) );
  MOAI22 U19299 ( .A1(n28912), .A2(n1641), .B1(ram[6137]), .B2(n1642), 
        .ZN(n10378) );
  MOAI22 U19300 ( .A1(n28677), .A2(n1641), .B1(ram[6138]), .B2(n1642), 
        .ZN(n10379) );
  MOAI22 U19301 ( .A1(n28442), .A2(n1641), .B1(ram[6139]), .B2(n1642), 
        .ZN(n10380) );
  MOAI22 U19302 ( .A1(n28207), .A2(n1641), .B1(ram[6140]), .B2(n1642), 
        .ZN(n10381) );
  MOAI22 U19303 ( .A1(n27972), .A2(n1641), .B1(ram[6141]), .B2(n1642), 
        .ZN(n10382) );
  MOAI22 U19304 ( .A1(n27737), .A2(n1641), .B1(ram[6142]), .B2(n1642), 
        .ZN(n10383) );
  MOAI22 U19305 ( .A1(n27502), .A2(n1641), .B1(ram[6143]), .B2(n1642), 
        .ZN(n10384) );
  MOAI22 U19306 ( .A1(n29147), .A2(n1643), .B1(ram[6144]), .B2(n1644), 
        .ZN(n10385) );
  MOAI22 U19307 ( .A1(n28912), .A2(n1643), .B1(ram[6145]), .B2(n1644), 
        .ZN(n10386) );
  MOAI22 U19308 ( .A1(n28677), .A2(n1643), .B1(ram[6146]), .B2(n1644), 
        .ZN(n10387) );
  MOAI22 U19309 ( .A1(n28442), .A2(n1643), .B1(ram[6147]), .B2(n1644), 
        .ZN(n10388) );
  MOAI22 U19310 ( .A1(n28207), .A2(n1643), .B1(ram[6148]), .B2(n1644), 
        .ZN(n10389) );
  MOAI22 U19311 ( .A1(n27972), .A2(n1643), .B1(ram[6149]), .B2(n1644), 
        .ZN(n10390) );
  MOAI22 U19312 ( .A1(n27737), .A2(n1643), .B1(ram[6150]), .B2(n1644), 
        .ZN(n10391) );
  MOAI22 U19313 ( .A1(n27502), .A2(n1643), .B1(ram[6151]), .B2(n1644), 
        .ZN(n10392) );
  MOAI22 U19314 ( .A1(n29147), .A2(n1646), .B1(ram[6152]), .B2(n1647), 
        .ZN(n10393) );
  MOAI22 U19315 ( .A1(n28912), .A2(n1646), .B1(ram[6153]), .B2(n1647), 
        .ZN(n10394) );
  MOAI22 U19316 ( .A1(n28677), .A2(n1646), .B1(ram[6154]), .B2(n1647), 
        .ZN(n10395) );
  MOAI22 U19317 ( .A1(n28442), .A2(n1646), .B1(ram[6155]), .B2(n1647), 
        .ZN(n10396) );
  MOAI22 U19318 ( .A1(n28207), .A2(n1646), .B1(ram[6156]), .B2(n1647), 
        .ZN(n10397) );
  MOAI22 U19319 ( .A1(n27972), .A2(n1646), .B1(ram[6157]), .B2(n1647), 
        .ZN(n10398) );
  MOAI22 U19320 ( .A1(n27737), .A2(n1646), .B1(ram[6158]), .B2(n1647), 
        .ZN(n10399) );
  MOAI22 U19321 ( .A1(n27502), .A2(n1646), .B1(ram[6159]), .B2(n1647), 
        .ZN(n10400) );
  MOAI22 U19322 ( .A1(n29147), .A2(n1648), .B1(ram[6160]), .B2(n1649), 
        .ZN(n10401) );
  MOAI22 U19323 ( .A1(n28912), .A2(n1648), .B1(ram[6161]), .B2(n1649), 
        .ZN(n10402) );
  MOAI22 U19324 ( .A1(n28677), .A2(n1648), .B1(ram[6162]), .B2(n1649), 
        .ZN(n10403) );
  MOAI22 U19325 ( .A1(n28442), .A2(n1648), .B1(ram[6163]), .B2(n1649), 
        .ZN(n10404) );
  MOAI22 U19326 ( .A1(n28207), .A2(n1648), .B1(ram[6164]), .B2(n1649), 
        .ZN(n10405) );
  MOAI22 U19327 ( .A1(n27972), .A2(n1648), .B1(ram[6165]), .B2(n1649), 
        .ZN(n10406) );
  MOAI22 U19328 ( .A1(n27737), .A2(n1648), .B1(ram[6166]), .B2(n1649), 
        .ZN(n10407) );
  MOAI22 U19329 ( .A1(n27502), .A2(n1648), .B1(ram[6167]), .B2(n1649), 
        .ZN(n10408) );
  MOAI22 U19330 ( .A1(n29147), .A2(n1650), .B1(ram[6168]), .B2(n1651), 
        .ZN(n10409) );
  MOAI22 U19331 ( .A1(n28912), .A2(n1650), .B1(ram[6169]), .B2(n1651), 
        .ZN(n10410) );
  MOAI22 U19332 ( .A1(n28677), .A2(n1650), .B1(ram[6170]), .B2(n1651), 
        .ZN(n10411) );
  MOAI22 U19333 ( .A1(n28442), .A2(n1650), .B1(ram[6171]), .B2(n1651), 
        .ZN(n10412) );
  MOAI22 U19334 ( .A1(n28207), .A2(n1650), .B1(ram[6172]), .B2(n1651), 
        .ZN(n10413) );
  MOAI22 U19335 ( .A1(n27972), .A2(n1650), .B1(ram[6173]), .B2(n1651), 
        .ZN(n10414) );
  MOAI22 U19336 ( .A1(n27737), .A2(n1650), .B1(ram[6174]), .B2(n1651), 
        .ZN(n10415) );
  MOAI22 U19337 ( .A1(n27502), .A2(n1650), .B1(ram[6175]), .B2(n1651), 
        .ZN(n10416) );
  MOAI22 U19338 ( .A1(n29147), .A2(n1652), .B1(ram[6176]), .B2(n1653), 
        .ZN(n10417) );
  MOAI22 U19339 ( .A1(n28912), .A2(n1652), .B1(ram[6177]), .B2(n1653), 
        .ZN(n10418) );
  MOAI22 U19340 ( .A1(n28677), .A2(n1652), .B1(ram[6178]), .B2(n1653), 
        .ZN(n10419) );
  MOAI22 U19341 ( .A1(n28442), .A2(n1652), .B1(ram[6179]), .B2(n1653), 
        .ZN(n10420) );
  MOAI22 U19342 ( .A1(n28207), .A2(n1652), .B1(ram[6180]), .B2(n1653), 
        .ZN(n10421) );
  MOAI22 U19343 ( .A1(n27972), .A2(n1652), .B1(ram[6181]), .B2(n1653), 
        .ZN(n10422) );
  MOAI22 U19344 ( .A1(n27737), .A2(n1652), .B1(ram[6182]), .B2(n1653), 
        .ZN(n10423) );
  MOAI22 U19345 ( .A1(n27502), .A2(n1652), .B1(ram[6183]), .B2(n1653), 
        .ZN(n10424) );
  MOAI22 U19346 ( .A1(n29147), .A2(n1654), .B1(ram[6184]), .B2(n1655), 
        .ZN(n10425) );
  MOAI22 U19347 ( .A1(n28912), .A2(n1654), .B1(ram[6185]), .B2(n1655), 
        .ZN(n10426) );
  MOAI22 U19348 ( .A1(n28677), .A2(n1654), .B1(ram[6186]), .B2(n1655), 
        .ZN(n10427) );
  MOAI22 U19349 ( .A1(n28442), .A2(n1654), .B1(ram[6187]), .B2(n1655), 
        .ZN(n10428) );
  MOAI22 U19350 ( .A1(n28207), .A2(n1654), .B1(ram[6188]), .B2(n1655), 
        .ZN(n10429) );
  MOAI22 U19351 ( .A1(n27972), .A2(n1654), .B1(ram[6189]), .B2(n1655), 
        .ZN(n10430) );
  MOAI22 U19352 ( .A1(n27737), .A2(n1654), .B1(ram[6190]), .B2(n1655), 
        .ZN(n10431) );
  MOAI22 U19353 ( .A1(n27502), .A2(n1654), .B1(ram[6191]), .B2(n1655), 
        .ZN(n10432) );
  MOAI22 U19354 ( .A1(n29147), .A2(n1656), .B1(ram[6192]), .B2(n1657), 
        .ZN(n10433) );
  MOAI22 U19355 ( .A1(n28912), .A2(n1656), .B1(ram[6193]), .B2(n1657), 
        .ZN(n10434) );
  MOAI22 U19356 ( .A1(n28677), .A2(n1656), .B1(ram[6194]), .B2(n1657), 
        .ZN(n10435) );
  MOAI22 U19357 ( .A1(n28442), .A2(n1656), .B1(ram[6195]), .B2(n1657), 
        .ZN(n10436) );
  MOAI22 U19358 ( .A1(n28207), .A2(n1656), .B1(ram[6196]), .B2(n1657), 
        .ZN(n10437) );
  MOAI22 U19359 ( .A1(n27972), .A2(n1656), .B1(ram[6197]), .B2(n1657), 
        .ZN(n10438) );
  MOAI22 U19360 ( .A1(n27737), .A2(n1656), .B1(ram[6198]), .B2(n1657), 
        .ZN(n10439) );
  MOAI22 U19361 ( .A1(n27502), .A2(n1656), .B1(ram[6199]), .B2(n1657), 
        .ZN(n10440) );
  MOAI22 U19362 ( .A1(n29147), .A2(n1658), .B1(ram[6200]), .B2(n1659), 
        .ZN(n10441) );
  MOAI22 U19363 ( .A1(n28912), .A2(n1658), .B1(ram[6201]), .B2(n1659), 
        .ZN(n10442) );
  MOAI22 U19364 ( .A1(n28677), .A2(n1658), .B1(ram[6202]), .B2(n1659), 
        .ZN(n10443) );
  MOAI22 U19365 ( .A1(n28442), .A2(n1658), .B1(ram[6203]), .B2(n1659), 
        .ZN(n10444) );
  MOAI22 U19366 ( .A1(n28207), .A2(n1658), .B1(ram[6204]), .B2(n1659), 
        .ZN(n10445) );
  MOAI22 U19367 ( .A1(n27972), .A2(n1658), .B1(ram[6205]), .B2(n1659), 
        .ZN(n10446) );
  MOAI22 U19368 ( .A1(n27737), .A2(n1658), .B1(ram[6206]), .B2(n1659), 
        .ZN(n10447) );
  MOAI22 U19369 ( .A1(n27502), .A2(n1658), .B1(ram[6207]), .B2(n1659), 
        .ZN(n10448) );
  MOAI22 U19370 ( .A1(n29147), .A2(n1660), .B1(ram[6208]), .B2(n1661), 
        .ZN(n10449) );
  MOAI22 U19371 ( .A1(n28912), .A2(n1660), .B1(ram[6209]), .B2(n1661), 
        .ZN(n10450) );
  MOAI22 U19372 ( .A1(n28677), .A2(n1660), .B1(ram[6210]), .B2(n1661), 
        .ZN(n10451) );
  MOAI22 U19373 ( .A1(n28442), .A2(n1660), .B1(ram[6211]), .B2(n1661), 
        .ZN(n10452) );
  MOAI22 U19374 ( .A1(n28207), .A2(n1660), .B1(ram[6212]), .B2(n1661), 
        .ZN(n10453) );
  MOAI22 U19375 ( .A1(n27972), .A2(n1660), .B1(ram[6213]), .B2(n1661), 
        .ZN(n10454) );
  MOAI22 U19376 ( .A1(n27737), .A2(n1660), .B1(ram[6214]), .B2(n1661), 
        .ZN(n10455) );
  MOAI22 U19377 ( .A1(n27502), .A2(n1660), .B1(ram[6215]), .B2(n1661), 
        .ZN(n10456) );
  MOAI22 U19378 ( .A1(n29147), .A2(n1662), .B1(ram[6216]), .B2(n1663), 
        .ZN(n10457) );
  MOAI22 U19379 ( .A1(n28912), .A2(n1662), .B1(ram[6217]), .B2(n1663), 
        .ZN(n10458) );
  MOAI22 U19380 ( .A1(n28677), .A2(n1662), .B1(ram[6218]), .B2(n1663), 
        .ZN(n10459) );
  MOAI22 U19381 ( .A1(n28442), .A2(n1662), .B1(ram[6219]), .B2(n1663), 
        .ZN(n10460) );
  MOAI22 U19382 ( .A1(n28207), .A2(n1662), .B1(ram[6220]), .B2(n1663), 
        .ZN(n10461) );
  MOAI22 U19383 ( .A1(n27972), .A2(n1662), .B1(ram[6221]), .B2(n1663), 
        .ZN(n10462) );
  MOAI22 U19384 ( .A1(n27737), .A2(n1662), .B1(ram[6222]), .B2(n1663), 
        .ZN(n10463) );
  MOAI22 U19385 ( .A1(n27502), .A2(n1662), .B1(ram[6223]), .B2(n1663), 
        .ZN(n10464) );
  MOAI22 U19386 ( .A1(n29147), .A2(n1664), .B1(ram[6224]), .B2(n1665), 
        .ZN(n10465) );
  MOAI22 U19387 ( .A1(n28912), .A2(n1664), .B1(ram[6225]), .B2(n1665), 
        .ZN(n10466) );
  MOAI22 U19388 ( .A1(n28677), .A2(n1664), .B1(ram[6226]), .B2(n1665), 
        .ZN(n10467) );
  MOAI22 U19389 ( .A1(n28442), .A2(n1664), .B1(ram[6227]), .B2(n1665), 
        .ZN(n10468) );
  MOAI22 U19390 ( .A1(n28207), .A2(n1664), .B1(ram[6228]), .B2(n1665), 
        .ZN(n10469) );
  MOAI22 U19391 ( .A1(n27972), .A2(n1664), .B1(ram[6229]), .B2(n1665), 
        .ZN(n10470) );
  MOAI22 U19392 ( .A1(n27737), .A2(n1664), .B1(ram[6230]), .B2(n1665), 
        .ZN(n10471) );
  MOAI22 U19393 ( .A1(n27502), .A2(n1664), .B1(ram[6231]), .B2(n1665), 
        .ZN(n10472) );
  MOAI22 U19394 ( .A1(n29147), .A2(n1666), .B1(ram[6232]), .B2(n1667), 
        .ZN(n10473) );
  MOAI22 U19395 ( .A1(n28912), .A2(n1666), .B1(ram[6233]), .B2(n1667), 
        .ZN(n10474) );
  MOAI22 U19396 ( .A1(n28677), .A2(n1666), .B1(ram[6234]), .B2(n1667), 
        .ZN(n10475) );
  MOAI22 U19397 ( .A1(n28442), .A2(n1666), .B1(ram[6235]), .B2(n1667), 
        .ZN(n10476) );
  MOAI22 U19398 ( .A1(n28207), .A2(n1666), .B1(ram[6236]), .B2(n1667), 
        .ZN(n10477) );
  MOAI22 U19399 ( .A1(n27972), .A2(n1666), .B1(ram[6237]), .B2(n1667), 
        .ZN(n10478) );
  MOAI22 U19400 ( .A1(n27737), .A2(n1666), .B1(ram[6238]), .B2(n1667), 
        .ZN(n10479) );
  MOAI22 U19401 ( .A1(n27502), .A2(n1666), .B1(ram[6239]), .B2(n1667), 
        .ZN(n10480) );
  MOAI22 U19402 ( .A1(n29148), .A2(n1668), .B1(ram[6240]), .B2(n1669), 
        .ZN(n10481) );
  MOAI22 U19403 ( .A1(n28913), .A2(n1668), .B1(ram[6241]), .B2(n1669), 
        .ZN(n10482) );
  MOAI22 U19404 ( .A1(n28678), .A2(n1668), .B1(ram[6242]), .B2(n1669), 
        .ZN(n10483) );
  MOAI22 U19405 ( .A1(n28443), .A2(n1668), .B1(ram[6243]), .B2(n1669), 
        .ZN(n10484) );
  MOAI22 U19406 ( .A1(n28208), .A2(n1668), .B1(ram[6244]), .B2(n1669), 
        .ZN(n10485) );
  MOAI22 U19407 ( .A1(n27973), .A2(n1668), .B1(ram[6245]), .B2(n1669), 
        .ZN(n10486) );
  MOAI22 U19408 ( .A1(n27738), .A2(n1668), .B1(ram[6246]), .B2(n1669), 
        .ZN(n10487) );
  MOAI22 U19409 ( .A1(n27503), .A2(n1668), .B1(ram[6247]), .B2(n1669), 
        .ZN(n10488) );
  MOAI22 U19410 ( .A1(n29148), .A2(n1670), .B1(ram[6248]), .B2(n1671), 
        .ZN(n10489) );
  MOAI22 U19411 ( .A1(n28913), .A2(n1670), .B1(ram[6249]), .B2(n1671), 
        .ZN(n10490) );
  MOAI22 U19412 ( .A1(n28678), .A2(n1670), .B1(ram[6250]), .B2(n1671), 
        .ZN(n10491) );
  MOAI22 U19413 ( .A1(n28443), .A2(n1670), .B1(ram[6251]), .B2(n1671), 
        .ZN(n10492) );
  MOAI22 U19414 ( .A1(n28208), .A2(n1670), .B1(ram[6252]), .B2(n1671), 
        .ZN(n10493) );
  MOAI22 U19415 ( .A1(n27973), .A2(n1670), .B1(ram[6253]), .B2(n1671), 
        .ZN(n10494) );
  MOAI22 U19416 ( .A1(n27738), .A2(n1670), .B1(ram[6254]), .B2(n1671), 
        .ZN(n10495) );
  MOAI22 U19417 ( .A1(n27503), .A2(n1670), .B1(ram[6255]), .B2(n1671), 
        .ZN(n10496) );
  MOAI22 U19418 ( .A1(n29148), .A2(n1672), .B1(ram[6256]), .B2(n1673), 
        .ZN(n10497) );
  MOAI22 U19419 ( .A1(n28913), .A2(n1672), .B1(ram[6257]), .B2(n1673), 
        .ZN(n10498) );
  MOAI22 U19420 ( .A1(n28678), .A2(n1672), .B1(ram[6258]), .B2(n1673), 
        .ZN(n10499) );
  MOAI22 U19421 ( .A1(n28443), .A2(n1672), .B1(ram[6259]), .B2(n1673), 
        .ZN(n10500) );
  MOAI22 U19422 ( .A1(n28208), .A2(n1672), .B1(ram[6260]), .B2(n1673), 
        .ZN(n10501) );
  MOAI22 U19423 ( .A1(n27973), .A2(n1672), .B1(ram[6261]), .B2(n1673), 
        .ZN(n10502) );
  MOAI22 U19424 ( .A1(n27738), .A2(n1672), .B1(ram[6262]), .B2(n1673), 
        .ZN(n10503) );
  MOAI22 U19425 ( .A1(n27503), .A2(n1672), .B1(ram[6263]), .B2(n1673), 
        .ZN(n10504) );
  MOAI22 U19426 ( .A1(n29148), .A2(n1674), .B1(ram[6264]), .B2(n1675), 
        .ZN(n10505) );
  MOAI22 U19427 ( .A1(n28913), .A2(n1674), .B1(ram[6265]), .B2(n1675), 
        .ZN(n10506) );
  MOAI22 U19428 ( .A1(n28678), .A2(n1674), .B1(ram[6266]), .B2(n1675), 
        .ZN(n10507) );
  MOAI22 U19429 ( .A1(n28443), .A2(n1674), .B1(ram[6267]), .B2(n1675), 
        .ZN(n10508) );
  MOAI22 U19430 ( .A1(n28208), .A2(n1674), .B1(ram[6268]), .B2(n1675), 
        .ZN(n10509) );
  MOAI22 U19431 ( .A1(n27973), .A2(n1674), .B1(ram[6269]), .B2(n1675), 
        .ZN(n10510) );
  MOAI22 U19432 ( .A1(n27738), .A2(n1674), .B1(ram[6270]), .B2(n1675), 
        .ZN(n10511) );
  MOAI22 U19433 ( .A1(n27503), .A2(n1674), .B1(ram[6271]), .B2(n1675), 
        .ZN(n10512) );
  MOAI22 U19434 ( .A1(n29148), .A2(n1676), .B1(ram[6272]), .B2(n1677), 
        .ZN(n10513) );
  MOAI22 U19435 ( .A1(n28913), .A2(n1676), .B1(ram[6273]), .B2(n1677), 
        .ZN(n10514) );
  MOAI22 U19436 ( .A1(n28678), .A2(n1676), .B1(ram[6274]), .B2(n1677), 
        .ZN(n10515) );
  MOAI22 U19437 ( .A1(n28443), .A2(n1676), .B1(ram[6275]), .B2(n1677), 
        .ZN(n10516) );
  MOAI22 U19438 ( .A1(n28208), .A2(n1676), .B1(ram[6276]), .B2(n1677), 
        .ZN(n10517) );
  MOAI22 U19439 ( .A1(n27973), .A2(n1676), .B1(ram[6277]), .B2(n1677), 
        .ZN(n10518) );
  MOAI22 U19440 ( .A1(n27738), .A2(n1676), .B1(ram[6278]), .B2(n1677), 
        .ZN(n10519) );
  MOAI22 U19441 ( .A1(n27503), .A2(n1676), .B1(ram[6279]), .B2(n1677), 
        .ZN(n10520) );
  MOAI22 U19442 ( .A1(n29148), .A2(n1678), .B1(ram[6280]), .B2(n1679), 
        .ZN(n10521) );
  MOAI22 U19443 ( .A1(n28913), .A2(n1678), .B1(ram[6281]), .B2(n1679), 
        .ZN(n10522) );
  MOAI22 U19444 ( .A1(n28678), .A2(n1678), .B1(ram[6282]), .B2(n1679), 
        .ZN(n10523) );
  MOAI22 U19445 ( .A1(n28443), .A2(n1678), .B1(ram[6283]), .B2(n1679), 
        .ZN(n10524) );
  MOAI22 U19446 ( .A1(n28208), .A2(n1678), .B1(ram[6284]), .B2(n1679), 
        .ZN(n10525) );
  MOAI22 U19447 ( .A1(n27973), .A2(n1678), .B1(ram[6285]), .B2(n1679), 
        .ZN(n10526) );
  MOAI22 U19448 ( .A1(n27738), .A2(n1678), .B1(ram[6286]), .B2(n1679), 
        .ZN(n10527) );
  MOAI22 U19449 ( .A1(n27503), .A2(n1678), .B1(ram[6287]), .B2(n1679), 
        .ZN(n10528) );
  MOAI22 U19450 ( .A1(n29148), .A2(n1680), .B1(ram[6288]), .B2(n1681), 
        .ZN(n10529) );
  MOAI22 U19451 ( .A1(n28913), .A2(n1680), .B1(ram[6289]), .B2(n1681), 
        .ZN(n10530) );
  MOAI22 U19452 ( .A1(n28678), .A2(n1680), .B1(ram[6290]), .B2(n1681), 
        .ZN(n10531) );
  MOAI22 U19453 ( .A1(n28443), .A2(n1680), .B1(ram[6291]), .B2(n1681), 
        .ZN(n10532) );
  MOAI22 U19454 ( .A1(n28208), .A2(n1680), .B1(ram[6292]), .B2(n1681), 
        .ZN(n10533) );
  MOAI22 U19455 ( .A1(n27973), .A2(n1680), .B1(ram[6293]), .B2(n1681), 
        .ZN(n10534) );
  MOAI22 U19456 ( .A1(n27738), .A2(n1680), .B1(ram[6294]), .B2(n1681), 
        .ZN(n10535) );
  MOAI22 U19457 ( .A1(n27503), .A2(n1680), .B1(ram[6295]), .B2(n1681), 
        .ZN(n10536) );
  MOAI22 U19458 ( .A1(n29148), .A2(n1682), .B1(ram[6296]), .B2(n1683), 
        .ZN(n10537) );
  MOAI22 U19459 ( .A1(n28913), .A2(n1682), .B1(ram[6297]), .B2(n1683), 
        .ZN(n10538) );
  MOAI22 U19460 ( .A1(n28678), .A2(n1682), .B1(ram[6298]), .B2(n1683), 
        .ZN(n10539) );
  MOAI22 U19461 ( .A1(n28443), .A2(n1682), .B1(ram[6299]), .B2(n1683), 
        .ZN(n10540) );
  MOAI22 U19462 ( .A1(n28208), .A2(n1682), .B1(ram[6300]), .B2(n1683), 
        .ZN(n10541) );
  MOAI22 U19463 ( .A1(n27973), .A2(n1682), .B1(ram[6301]), .B2(n1683), 
        .ZN(n10542) );
  MOAI22 U19464 ( .A1(n27738), .A2(n1682), .B1(ram[6302]), .B2(n1683), 
        .ZN(n10543) );
  MOAI22 U19465 ( .A1(n27503), .A2(n1682), .B1(ram[6303]), .B2(n1683), 
        .ZN(n10544) );
  MOAI22 U19466 ( .A1(n29148), .A2(n1684), .B1(ram[6304]), .B2(n1685), 
        .ZN(n10545) );
  MOAI22 U19467 ( .A1(n28913), .A2(n1684), .B1(ram[6305]), .B2(n1685), 
        .ZN(n10546) );
  MOAI22 U19468 ( .A1(n28678), .A2(n1684), .B1(ram[6306]), .B2(n1685), 
        .ZN(n10547) );
  MOAI22 U19469 ( .A1(n28443), .A2(n1684), .B1(ram[6307]), .B2(n1685), 
        .ZN(n10548) );
  MOAI22 U19470 ( .A1(n28208), .A2(n1684), .B1(ram[6308]), .B2(n1685), 
        .ZN(n10549) );
  MOAI22 U19471 ( .A1(n27973), .A2(n1684), .B1(ram[6309]), .B2(n1685), 
        .ZN(n10550) );
  MOAI22 U19472 ( .A1(n27738), .A2(n1684), .B1(ram[6310]), .B2(n1685), 
        .ZN(n10551) );
  MOAI22 U19473 ( .A1(n27503), .A2(n1684), .B1(ram[6311]), .B2(n1685), 
        .ZN(n10552) );
  MOAI22 U19474 ( .A1(n29148), .A2(n1686), .B1(ram[6312]), .B2(n1687), 
        .ZN(n10553) );
  MOAI22 U19475 ( .A1(n28913), .A2(n1686), .B1(ram[6313]), .B2(n1687), 
        .ZN(n10554) );
  MOAI22 U19476 ( .A1(n28678), .A2(n1686), .B1(ram[6314]), .B2(n1687), 
        .ZN(n10555) );
  MOAI22 U19477 ( .A1(n28443), .A2(n1686), .B1(ram[6315]), .B2(n1687), 
        .ZN(n10556) );
  MOAI22 U19478 ( .A1(n28208), .A2(n1686), .B1(ram[6316]), .B2(n1687), 
        .ZN(n10557) );
  MOAI22 U19479 ( .A1(n27973), .A2(n1686), .B1(ram[6317]), .B2(n1687), 
        .ZN(n10558) );
  MOAI22 U19480 ( .A1(n27738), .A2(n1686), .B1(ram[6318]), .B2(n1687), 
        .ZN(n10559) );
  MOAI22 U19481 ( .A1(n27503), .A2(n1686), .B1(ram[6319]), .B2(n1687), 
        .ZN(n10560) );
  MOAI22 U19482 ( .A1(n29148), .A2(n1688), .B1(ram[6320]), .B2(n1689), 
        .ZN(n10561) );
  MOAI22 U19483 ( .A1(n28913), .A2(n1688), .B1(ram[6321]), .B2(n1689), 
        .ZN(n10562) );
  MOAI22 U19484 ( .A1(n28678), .A2(n1688), .B1(ram[6322]), .B2(n1689), 
        .ZN(n10563) );
  MOAI22 U19485 ( .A1(n28443), .A2(n1688), .B1(ram[6323]), .B2(n1689), 
        .ZN(n10564) );
  MOAI22 U19486 ( .A1(n28208), .A2(n1688), .B1(ram[6324]), .B2(n1689), 
        .ZN(n10565) );
  MOAI22 U19487 ( .A1(n27973), .A2(n1688), .B1(ram[6325]), .B2(n1689), 
        .ZN(n10566) );
  MOAI22 U19488 ( .A1(n27738), .A2(n1688), .B1(ram[6326]), .B2(n1689), 
        .ZN(n10567) );
  MOAI22 U19489 ( .A1(n27503), .A2(n1688), .B1(ram[6327]), .B2(n1689), 
        .ZN(n10568) );
  MOAI22 U19490 ( .A1(n29148), .A2(n1690), .B1(ram[6328]), .B2(n1691), 
        .ZN(n10569) );
  MOAI22 U19491 ( .A1(n28913), .A2(n1690), .B1(ram[6329]), .B2(n1691), 
        .ZN(n10570) );
  MOAI22 U19492 ( .A1(n28678), .A2(n1690), .B1(ram[6330]), .B2(n1691), 
        .ZN(n10571) );
  MOAI22 U19493 ( .A1(n28443), .A2(n1690), .B1(ram[6331]), .B2(n1691), 
        .ZN(n10572) );
  MOAI22 U19494 ( .A1(n28208), .A2(n1690), .B1(ram[6332]), .B2(n1691), 
        .ZN(n10573) );
  MOAI22 U19495 ( .A1(n27973), .A2(n1690), .B1(ram[6333]), .B2(n1691), 
        .ZN(n10574) );
  MOAI22 U19496 ( .A1(n27738), .A2(n1690), .B1(ram[6334]), .B2(n1691), 
        .ZN(n10575) );
  MOAI22 U19497 ( .A1(n27503), .A2(n1690), .B1(ram[6335]), .B2(n1691), 
        .ZN(n10576) );
  MOAI22 U19498 ( .A1(n29148), .A2(n1692), .B1(ram[6336]), .B2(n1693), 
        .ZN(n10577) );
  MOAI22 U19499 ( .A1(n28913), .A2(n1692), .B1(ram[6337]), .B2(n1693), 
        .ZN(n10578) );
  MOAI22 U19500 ( .A1(n28678), .A2(n1692), .B1(ram[6338]), .B2(n1693), 
        .ZN(n10579) );
  MOAI22 U19501 ( .A1(n28443), .A2(n1692), .B1(ram[6339]), .B2(n1693), 
        .ZN(n10580) );
  MOAI22 U19502 ( .A1(n28208), .A2(n1692), .B1(ram[6340]), .B2(n1693), 
        .ZN(n10581) );
  MOAI22 U19503 ( .A1(n27973), .A2(n1692), .B1(ram[6341]), .B2(n1693), 
        .ZN(n10582) );
  MOAI22 U19504 ( .A1(n27738), .A2(n1692), .B1(ram[6342]), .B2(n1693), 
        .ZN(n10583) );
  MOAI22 U19505 ( .A1(n27503), .A2(n1692), .B1(ram[6343]), .B2(n1693), 
        .ZN(n10584) );
  MOAI22 U19506 ( .A1(n29149), .A2(n1694), .B1(ram[6344]), .B2(n1695), 
        .ZN(n10585) );
  MOAI22 U19507 ( .A1(n28914), .A2(n1694), .B1(ram[6345]), .B2(n1695), 
        .ZN(n10586) );
  MOAI22 U19508 ( .A1(n28679), .A2(n1694), .B1(ram[6346]), .B2(n1695), 
        .ZN(n10587) );
  MOAI22 U19509 ( .A1(n28444), .A2(n1694), .B1(ram[6347]), .B2(n1695), 
        .ZN(n10588) );
  MOAI22 U19510 ( .A1(n28209), .A2(n1694), .B1(ram[6348]), .B2(n1695), 
        .ZN(n10589) );
  MOAI22 U19511 ( .A1(n27974), .A2(n1694), .B1(ram[6349]), .B2(n1695), 
        .ZN(n10590) );
  MOAI22 U19512 ( .A1(n27739), .A2(n1694), .B1(ram[6350]), .B2(n1695), 
        .ZN(n10591) );
  MOAI22 U19513 ( .A1(n27504), .A2(n1694), .B1(ram[6351]), .B2(n1695), 
        .ZN(n10592) );
  MOAI22 U19514 ( .A1(n29149), .A2(n1696), .B1(ram[6352]), .B2(n1697), 
        .ZN(n10593) );
  MOAI22 U19515 ( .A1(n28914), .A2(n1696), .B1(ram[6353]), .B2(n1697), 
        .ZN(n10594) );
  MOAI22 U19516 ( .A1(n28679), .A2(n1696), .B1(ram[6354]), .B2(n1697), 
        .ZN(n10595) );
  MOAI22 U19517 ( .A1(n28444), .A2(n1696), .B1(ram[6355]), .B2(n1697), 
        .ZN(n10596) );
  MOAI22 U19518 ( .A1(n28209), .A2(n1696), .B1(ram[6356]), .B2(n1697), 
        .ZN(n10597) );
  MOAI22 U19519 ( .A1(n27974), .A2(n1696), .B1(ram[6357]), .B2(n1697), 
        .ZN(n10598) );
  MOAI22 U19520 ( .A1(n27739), .A2(n1696), .B1(ram[6358]), .B2(n1697), 
        .ZN(n10599) );
  MOAI22 U19521 ( .A1(n27504), .A2(n1696), .B1(ram[6359]), .B2(n1697), 
        .ZN(n10600) );
  MOAI22 U19522 ( .A1(n29149), .A2(n1698), .B1(ram[6360]), .B2(n1699), 
        .ZN(n10601) );
  MOAI22 U19523 ( .A1(n28914), .A2(n1698), .B1(ram[6361]), .B2(n1699), 
        .ZN(n10602) );
  MOAI22 U19524 ( .A1(n28679), .A2(n1698), .B1(ram[6362]), .B2(n1699), 
        .ZN(n10603) );
  MOAI22 U19525 ( .A1(n28444), .A2(n1698), .B1(ram[6363]), .B2(n1699), 
        .ZN(n10604) );
  MOAI22 U19526 ( .A1(n28209), .A2(n1698), .B1(ram[6364]), .B2(n1699), 
        .ZN(n10605) );
  MOAI22 U19527 ( .A1(n27974), .A2(n1698), .B1(ram[6365]), .B2(n1699), 
        .ZN(n10606) );
  MOAI22 U19528 ( .A1(n27739), .A2(n1698), .B1(ram[6366]), .B2(n1699), 
        .ZN(n10607) );
  MOAI22 U19529 ( .A1(n27504), .A2(n1698), .B1(ram[6367]), .B2(n1699), 
        .ZN(n10608) );
  MOAI22 U19530 ( .A1(n29149), .A2(n1700), .B1(ram[6368]), .B2(n1701), 
        .ZN(n10609) );
  MOAI22 U19531 ( .A1(n28914), .A2(n1700), .B1(ram[6369]), .B2(n1701), 
        .ZN(n10610) );
  MOAI22 U19532 ( .A1(n28679), .A2(n1700), .B1(ram[6370]), .B2(n1701), 
        .ZN(n10611) );
  MOAI22 U19533 ( .A1(n28444), .A2(n1700), .B1(ram[6371]), .B2(n1701), 
        .ZN(n10612) );
  MOAI22 U19534 ( .A1(n28209), .A2(n1700), .B1(ram[6372]), .B2(n1701), 
        .ZN(n10613) );
  MOAI22 U19535 ( .A1(n27974), .A2(n1700), .B1(ram[6373]), .B2(n1701), 
        .ZN(n10614) );
  MOAI22 U19536 ( .A1(n27739), .A2(n1700), .B1(ram[6374]), .B2(n1701), 
        .ZN(n10615) );
  MOAI22 U19537 ( .A1(n27504), .A2(n1700), .B1(ram[6375]), .B2(n1701), 
        .ZN(n10616) );
  MOAI22 U19538 ( .A1(n29149), .A2(n1702), .B1(ram[6376]), .B2(n1703), 
        .ZN(n10617) );
  MOAI22 U19539 ( .A1(n28914), .A2(n1702), .B1(ram[6377]), .B2(n1703), 
        .ZN(n10618) );
  MOAI22 U19540 ( .A1(n28679), .A2(n1702), .B1(ram[6378]), .B2(n1703), 
        .ZN(n10619) );
  MOAI22 U19541 ( .A1(n28444), .A2(n1702), .B1(ram[6379]), .B2(n1703), 
        .ZN(n10620) );
  MOAI22 U19542 ( .A1(n28209), .A2(n1702), .B1(ram[6380]), .B2(n1703), 
        .ZN(n10621) );
  MOAI22 U19543 ( .A1(n27974), .A2(n1702), .B1(ram[6381]), .B2(n1703), 
        .ZN(n10622) );
  MOAI22 U19544 ( .A1(n27739), .A2(n1702), .B1(ram[6382]), .B2(n1703), 
        .ZN(n10623) );
  MOAI22 U19545 ( .A1(n27504), .A2(n1702), .B1(ram[6383]), .B2(n1703), 
        .ZN(n10624) );
  MOAI22 U19546 ( .A1(n29149), .A2(n1704), .B1(ram[6384]), .B2(n1705), 
        .ZN(n10625) );
  MOAI22 U19547 ( .A1(n28914), .A2(n1704), .B1(ram[6385]), .B2(n1705), 
        .ZN(n10626) );
  MOAI22 U19548 ( .A1(n28679), .A2(n1704), .B1(ram[6386]), .B2(n1705), 
        .ZN(n10627) );
  MOAI22 U19549 ( .A1(n28444), .A2(n1704), .B1(ram[6387]), .B2(n1705), 
        .ZN(n10628) );
  MOAI22 U19550 ( .A1(n28209), .A2(n1704), .B1(ram[6388]), .B2(n1705), 
        .ZN(n10629) );
  MOAI22 U19551 ( .A1(n27974), .A2(n1704), .B1(ram[6389]), .B2(n1705), 
        .ZN(n10630) );
  MOAI22 U19552 ( .A1(n27739), .A2(n1704), .B1(ram[6390]), .B2(n1705), 
        .ZN(n10631) );
  MOAI22 U19553 ( .A1(n27504), .A2(n1704), .B1(ram[6391]), .B2(n1705), 
        .ZN(n10632) );
  MOAI22 U19554 ( .A1(n29149), .A2(n1706), .B1(ram[6392]), .B2(n1707), 
        .ZN(n10633) );
  MOAI22 U19555 ( .A1(n28914), .A2(n1706), .B1(ram[6393]), .B2(n1707), 
        .ZN(n10634) );
  MOAI22 U19556 ( .A1(n28679), .A2(n1706), .B1(ram[6394]), .B2(n1707), 
        .ZN(n10635) );
  MOAI22 U19557 ( .A1(n28444), .A2(n1706), .B1(ram[6395]), .B2(n1707), 
        .ZN(n10636) );
  MOAI22 U19558 ( .A1(n28209), .A2(n1706), .B1(ram[6396]), .B2(n1707), 
        .ZN(n10637) );
  MOAI22 U19559 ( .A1(n27974), .A2(n1706), .B1(ram[6397]), .B2(n1707), 
        .ZN(n10638) );
  MOAI22 U19560 ( .A1(n27739), .A2(n1706), .B1(ram[6398]), .B2(n1707), 
        .ZN(n10639) );
  MOAI22 U19561 ( .A1(n27504), .A2(n1706), .B1(ram[6399]), .B2(n1707), 
        .ZN(n10640) );
  MOAI22 U19562 ( .A1(n29149), .A2(n1708), .B1(ram[6400]), .B2(n1709), 
        .ZN(n10641) );
  MOAI22 U19563 ( .A1(n28914), .A2(n1708), .B1(ram[6401]), .B2(n1709), 
        .ZN(n10642) );
  MOAI22 U19564 ( .A1(n28679), .A2(n1708), .B1(ram[6402]), .B2(n1709), 
        .ZN(n10643) );
  MOAI22 U19565 ( .A1(n28444), .A2(n1708), .B1(ram[6403]), .B2(n1709), 
        .ZN(n10644) );
  MOAI22 U19566 ( .A1(n28209), .A2(n1708), .B1(ram[6404]), .B2(n1709), 
        .ZN(n10645) );
  MOAI22 U19567 ( .A1(n27974), .A2(n1708), .B1(ram[6405]), .B2(n1709), 
        .ZN(n10646) );
  MOAI22 U19568 ( .A1(n27739), .A2(n1708), .B1(ram[6406]), .B2(n1709), 
        .ZN(n10647) );
  MOAI22 U19569 ( .A1(n27504), .A2(n1708), .B1(ram[6407]), .B2(n1709), 
        .ZN(n10648) );
  MOAI22 U19570 ( .A1(n29149), .A2(n1710), .B1(ram[6408]), .B2(n1711), 
        .ZN(n10649) );
  MOAI22 U19571 ( .A1(n28914), .A2(n1710), .B1(ram[6409]), .B2(n1711), 
        .ZN(n10650) );
  MOAI22 U19572 ( .A1(n28679), .A2(n1710), .B1(ram[6410]), .B2(n1711), 
        .ZN(n10651) );
  MOAI22 U19573 ( .A1(n28444), .A2(n1710), .B1(ram[6411]), .B2(n1711), 
        .ZN(n10652) );
  MOAI22 U19574 ( .A1(n28209), .A2(n1710), .B1(ram[6412]), .B2(n1711), 
        .ZN(n10653) );
  MOAI22 U19575 ( .A1(n27974), .A2(n1710), .B1(ram[6413]), .B2(n1711), 
        .ZN(n10654) );
  MOAI22 U19576 ( .A1(n27739), .A2(n1710), .B1(ram[6414]), .B2(n1711), 
        .ZN(n10655) );
  MOAI22 U19577 ( .A1(n27504), .A2(n1710), .B1(ram[6415]), .B2(n1711), 
        .ZN(n10656) );
  MOAI22 U19578 ( .A1(n29149), .A2(n1712), .B1(ram[6416]), .B2(n1713), 
        .ZN(n10657) );
  MOAI22 U19579 ( .A1(n28914), .A2(n1712), .B1(ram[6417]), .B2(n1713), 
        .ZN(n10658) );
  MOAI22 U19580 ( .A1(n28679), .A2(n1712), .B1(ram[6418]), .B2(n1713), 
        .ZN(n10659) );
  MOAI22 U19581 ( .A1(n28444), .A2(n1712), .B1(ram[6419]), .B2(n1713), 
        .ZN(n10660) );
  MOAI22 U19582 ( .A1(n28209), .A2(n1712), .B1(ram[6420]), .B2(n1713), 
        .ZN(n10661) );
  MOAI22 U19583 ( .A1(n27974), .A2(n1712), .B1(ram[6421]), .B2(n1713), 
        .ZN(n10662) );
  MOAI22 U19584 ( .A1(n27739), .A2(n1712), .B1(ram[6422]), .B2(n1713), 
        .ZN(n10663) );
  MOAI22 U19585 ( .A1(n27504), .A2(n1712), .B1(ram[6423]), .B2(n1713), 
        .ZN(n10664) );
  MOAI22 U19586 ( .A1(n29149), .A2(n1714), .B1(ram[6424]), .B2(n1715), 
        .ZN(n10665) );
  MOAI22 U19587 ( .A1(n28914), .A2(n1714), .B1(ram[6425]), .B2(n1715), 
        .ZN(n10666) );
  MOAI22 U19588 ( .A1(n28679), .A2(n1714), .B1(ram[6426]), .B2(n1715), 
        .ZN(n10667) );
  MOAI22 U19589 ( .A1(n28444), .A2(n1714), .B1(ram[6427]), .B2(n1715), 
        .ZN(n10668) );
  MOAI22 U19590 ( .A1(n28209), .A2(n1714), .B1(ram[6428]), .B2(n1715), 
        .ZN(n10669) );
  MOAI22 U19591 ( .A1(n27974), .A2(n1714), .B1(ram[6429]), .B2(n1715), 
        .ZN(n10670) );
  MOAI22 U19592 ( .A1(n27739), .A2(n1714), .B1(ram[6430]), .B2(n1715), 
        .ZN(n10671) );
  MOAI22 U19593 ( .A1(n27504), .A2(n1714), .B1(ram[6431]), .B2(n1715), 
        .ZN(n10672) );
  MOAI22 U19594 ( .A1(n29149), .A2(n1716), .B1(ram[6432]), .B2(n1717), 
        .ZN(n10673) );
  MOAI22 U19595 ( .A1(n28914), .A2(n1716), .B1(ram[6433]), .B2(n1717), 
        .ZN(n10674) );
  MOAI22 U19596 ( .A1(n28679), .A2(n1716), .B1(ram[6434]), .B2(n1717), 
        .ZN(n10675) );
  MOAI22 U19597 ( .A1(n28444), .A2(n1716), .B1(ram[6435]), .B2(n1717), 
        .ZN(n10676) );
  MOAI22 U19598 ( .A1(n28209), .A2(n1716), .B1(ram[6436]), .B2(n1717), 
        .ZN(n10677) );
  MOAI22 U19599 ( .A1(n27974), .A2(n1716), .B1(ram[6437]), .B2(n1717), 
        .ZN(n10678) );
  MOAI22 U19600 ( .A1(n27739), .A2(n1716), .B1(ram[6438]), .B2(n1717), 
        .ZN(n10679) );
  MOAI22 U19601 ( .A1(n27504), .A2(n1716), .B1(ram[6439]), .B2(n1717), 
        .ZN(n10680) );
  MOAI22 U19602 ( .A1(n29149), .A2(n1718), .B1(ram[6440]), .B2(n1719), 
        .ZN(n10681) );
  MOAI22 U19603 ( .A1(n28914), .A2(n1718), .B1(ram[6441]), .B2(n1719), 
        .ZN(n10682) );
  MOAI22 U19604 ( .A1(n28679), .A2(n1718), .B1(ram[6442]), .B2(n1719), 
        .ZN(n10683) );
  MOAI22 U19605 ( .A1(n28444), .A2(n1718), .B1(ram[6443]), .B2(n1719), 
        .ZN(n10684) );
  MOAI22 U19606 ( .A1(n28209), .A2(n1718), .B1(ram[6444]), .B2(n1719), 
        .ZN(n10685) );
  MOAI22 U19607 ( .A1(n27974), .A2(n1718), .B1(ram[6445]), .B2(n1719), 
        .ZN(n10686) );
  MOAI22 U19608 ( .A1(n27739), .A2(n1718), .B1(ram[6446]), .B2(n1719), 
        .ZN(n10687) );
  MOAI22 U19609 ( .A1(n27504), .A2(n1718), .B1(ram[6447]), .B2(n1719), 
        .ZN(n10688) );
  MOAI22 U19610 ( .A1(n29150), .A2(n1720), .B1(ram[6448]), .B2(n1721), 
        .ZN(n10689) );
  MOAI22 U19611 ( .A1(n28915), .A2(n1720), .B1(ram[6449]), .B2(n1721), 
        .ZN(n10690) );
  MOAI22 U19612 ( .A1(n28680), .A2(n1720), .B1(ram[6450]), .B2(n1721), 
        .ZN(n10691) );
  MOAI22 U19613 ( .A1(n28445), .A2(n1720), .B1(ram[6451]), .B2(n1721), 
        .ZN(n10692) );
  MOAI22 U19614 ( .A1(n28210), .A2(n1720), .B1(ram[6452]), .B2(n1721), 
        .ZN(n10693) );
  MOAI22 U19615 ( .A1(n27975), .A2(n1720), .B1(ram[6453]), .B2(n1721), 
        .ZN(n10694) );
  MOAI22 U19616 ( .A1(n27740), .A2(n1720), .B1(ram[6454]), .B2(n1721), 
        .ZN(n10695) );
  MOAI22 U19617 ( .A1(n27505), .A2(n1720), .B1(ram[6455]), .B2(n1721), 
        .ZN(n10696) );
  MOAI22 U19618 ( .A1(n29150), .A2(n1722), .B1(ram[6456]), .B2(n1723), 
        .ZN(n10697) );
  MOAI22 U19619 ( .A1(n28915), .A2(n1722), .B1(ram[6457]), .B2(n1723), 
        .ZN(n10698) );
  MOAI22 U19620 ( .A1(n28680), .A2(n1722), .B1(ram[6458]), .B2(n1723), 
        .ZN(n10699) );
  MOAI22 U19621 ( .A1(n28445), .A2(n1722), .B1(ram[6459]), .B2(n1723), 
        .ZN(n10700) );
  MOAI22 U19622 ( .A1(n28210), .A2(n1722), .B1(ram[6460]), .B2(n1723), 
        .ZN(n10701) );
  MOAI22 U19623 ( .A1(n27975), .A2(n1722), .B1(ram[6461]), .B2(n1723), 
        .ZN(n10702) );
  MOAI22 U19624 ( .A1(n27740), .A2(n1722), .B1(ram[6462]), .B2(n1723), 
        .ZN(n10703) );
  MOAI22 U19625 ( .A1(n27505), .A2(n1722), .B1(ram[6463]), .B2(n1723), 
        .ZN(n10704) );
  MOAI22 U19626 ( .A1(n29150), .A2(n1724), .B1(ram[6464]), .B2(n1725), 
        .ZN(n10705) );
  MOAI22 U19627 ( .A1(n28915), .A2(n1724), .B1(ram[6465]), .B2(n1725), 
        .ZN(n10706) );
  MOAI22 U19628 ( .A1(n28680), .A2(n1724), .B1(ram[6466]), .B2(n1725), 
        .ZN(n10707) );
  MOAI22 U19629 ( .A1(n28445), .A2(n1724), .B1(ram[6467]), .B2(n1725), 
        .ZN(n10708) );
  MOAI22 U19630 ( .A1(n28210), .A2(n1724), .B1(ram[6468]), .B2(n1725), 
        .ZN(n10709) );
  MOAI22 U19631 ( .A1(n27975), .A2(n1724), .B1(ram[6469]), .B2(n1725), 
        .ZN(n10710) );
  MOAI22 U19632 ( .A1(n27740), .A2(n1724), .B1(ram[6470]), .B2(n1725), 
        .ZN(n10711) );
  MOAI22 U19633 ( .A1(n27505), .A2(n1724), .B1(ram[6471]), .B2(n1725), 
        .ZN(n10712) );
  MOAI22 U19634 ( .A1(n29150), .A2(n1726), .B1(ram[6472]), .B2(n1727), 
        .ZN(n10713) );
  MOAI22 U19635 ( .A1(n28915), .A2(n1726), .B1(ram[6473]), .B2(n1727), 
        .ZN(n10714) );
  MOAI22 U19636 ( .A1(n28680), .A2(n1726), .B1(ram[6474]), .B2(n1727), 
        .ZN(n10715) );
  MOAI22 U19637 ( .A1(n28445), .A2(n1726), .B1(ram[6475]), .B2(n1727), 
        .ZN(n10716) );
  MOAI22 U19638 ( .A1(n28210), .A2(n1726), .B1(ram[6476]), .B2(n1727), 
        .ZN(n10717) );
  MOAI22 U19639 ( .A1(n27975), .A2(n1726), .B1(ram[6477]), .B2(n1727), 
        .ZN(n10718) );
  MOAI22 U19640 ( .A1(n27740), .A2(n1726), .B1(ram[6478]), .B2(n1727), 
        .ZN(n10719) );
  MOAI22 U19641 ( .A1(n27505), .A2(n1726), .B1(ram[6479]), .B2(n1727), 
        .ZN(n10720) );
  MOAI22 U19642 ( .A1(n29150), .A2(n1728), .B1(ram[6480]), .B2(n1729), 
        .ZN(n10721) );
  MOAI22 U19643 ( .A1(n28915), .A2(n1728), .B1(ram[6481]), .B2(n1729), 
        .ZN(n10722) );
  MOAI22 U19644 ( .A1(n28680), .A2(n1728), .B1(ram[6482]), .B2(n1729), 
        .ZN(n10723) );
  MOAI22 U19645 ( .A1(n28445), .A2(n1728), .B1(ram[6483]), .B2(n1729), 
        .ZN(n10724) );
  MOAI22 U19646 ( .A1(n28210), .A2(n1728), .B1(ram[6484]), .B2(n1729), 
        .ZN(n10725) );
  MOAI22 U19647 ( .A1(n27975), .A2(n1728), .B1(ram[6485]), .B2(n1729), 
        .ZN(n10726) );
  MOAI22 U19648 ( .A1(n27740), .A2(n1728), .B1(ram[6486]), .B2(n1729), 
        .ZN(n10727) );
  MOAI22 U19649 ( .A1(n27505), .A2(n1728), .B1(ram[6487]), .B2(n1729), 
        .ZN(n10728) );
  MOAI22 U19650 ( .A1(n29150), .A2(n1730), .B1(ram[6488]), .B2(n1731), 
        .ZN(n10729) );
  MOAI22 U19651 ( .A1(n28915), .A2(n1730), .B1(ram[6489]), .B2(n1731), 
        .ZN(n10730) );
  MOAI22 U19652 ( .A1(n28680), .A2(n1730), .B1(ram[6490]), .B2(n1731), 
        .ZN(n10731) );
  MOAI22 U19653 ( .A1(n28445), .A2(n1730), .B1(ram[6491]), .B2(n1731), 
        .ZN(n10732) );
  MOAI22 U19654 ( .A1(n28210), .A2(n1730), .B1(ram[6492]), .B2(n1731), 
        .ZN(n10733) );
  MOAI22 U19655 ( .A1(n27975), .A2(n1730), .B1(ram[6493]), .B2(n1731), 
        .ZN(n10734) );
  MOAI22 U19656 ( .A1(n27740), .A2(n1730), .B1(ram[6494]), .B2(n1731), 
        .ZN(n10735) );
  MOAI22 U19657 ( .A1(n27505), .A2(n1730), .B1(ram[6495]), .B2(n1731), 
        .ZN(n10736) );
  MOAI22 U19658 ( .A1(n29150), .A2(n1732), .B1(ram[6496]), .B2(n1733), 
        .ZN(n10737) );
  MOAI22 U19659 ( .A1(n28915), .A2(n1732), .B1(ram[6497]), .B2(n1733), 
        .ZN(n10738) );
  MOAI22 U19660 ( .A1(n28680), .A2(n1732), .B1(ram[6498]), .B2(n1733), 
        .ZN(n10739) );
  MOAI22 U19661 ( .A1(n28445), .A2(n1732), .B1(ram[6499]), .B2(n1733), 
        .ZN(n10740) );
  MOAI22 U19662 ( .A1(n28210), .A2(n1732), .B1(ram[6500]), .B2(n1733), 
        .ZN(n10741) );
  MOAI22 U19663 ( .A1(n27975), .A2(n1732), .B1(ram[6501]), .B2(n1733), 
        .ZN(n10742) );
  MOAI22 U19664 ( .A1(n27740), .A2(n1732), .B1(ram[6502]), .B2(n1733), 
        .ZN(n10743) );
  MOAI22 U19665 ( .A1(n27505), .A2(n1732), .B1(ram[6503]), .B2(n1733), 
        .ZN(n10744) );
  MOAI22 U19666 ( .A1(n29150), .A2(n1734), .B1(ram[6504]), .B2(n1735), 
        .ZN(n10745) );
  MOAI22 U19667 ( .A1(n28915), .A2(n1734), .B1(ram[6505]), .B2(n1735), 
        .ZN(n10746) );
  MOAI22 U19668 ( .A1(n28680), .A2(n1734), .B1(ram[6506]), .B2(n1735), 
        .ZN(n10747) );
  MOAI22 U19669 ( .A1(n28445), .A2(n1734), .B1(ram[6507]), .B2(n1735), 
        .ZN(n10748) );
  MOAI22 U19670 ( .A1(n28210), .A2(n1734), .B1(ram[6508]), .B2(n1735), 
        .ZN(n10749) );
  MOAI22 U19671 ( .A1(n27975), .A2(n1734), .B1(ram[6509]), .B2(n1735), 
        .ZN(n10750) );
  MOAI22 U19672 ( .A1(n27740), .A2(n1734), .B1(ram[6510]), .B2(n1735), 
        .ZN(n10751) );
  MOAI22 U19673 ( .A1(n27505), .A2(n1734), .B1(ram[6511]), .B2(n1735), 
        .ZN(n10752) );
  MOAI22 U19674 ( .A1(n29150), .A2(n1736), .B1(ram[6512]), .B2(n1737), 
        .ZN(n10753) );
  MOAI22 U19675 ( .A1(n28915), .A2(n1736), .B1(ram[6513]), .B2(n1737), 
        .ZN(n10754) );
  MOAI22 U19676 ( .A1(n28680), .A2(n1736), .B1(ram[6514]), .B2(n1737), 
        .ZN(n10755) );
  MOAI22 U19677 ( .A1(n28445), .A2(n1736), .B1(ram[6515]), .B2(n1737), 
        .ZN(n10756) );
  MOAI22 U19678 ( .A1(n28210), .A2(n1736), .B1(ram[6516]), .B2(n1737), 
        .ZN(n10757) );
  MOAI22 U19679 ( .A1(n27975), .A2(n1736), .B1(ram[6517]), .B2(n1737), 
        .ZN(n10758) );
  MOAI22 U19680 ( .A1(n27740), .A2(n1736), .B1(ram[6518]), .B2(n1737), 
        .ZN(n10759) );
  MOAI22 U19681 ( .A1(n27505), .A2(n1736), .B1(ram[6519]), .B2(n1737), 
        .ZN(n10760) );
  MOAI22 U19682 ( .A1(n29150), .A2(n1738), .B1(ram[6520]), .B2(n1739), 
        .ZN(n10761) );
  MOAI22 U19683 ( .A1(n28915), .A2(n1738), .B1(ram[6521]), .B2(n1739), 
        .ZN(n10762) );
  MOAI22 U19684 ( .A1(n28680), .A2(n1738), .B1(ram[6522]), .B2(n1739), 
        .ZN(n10763) );
  MOAI22 U19685 ( .A1(n28445), .A2(n1738), .B1(ram[6523]), .B2(n1739), 
        .ZN(n10764) );
  MOAI22 U19686 ( .A1(n28210), .A2(n1738), .B1(ram[6524]), .B2(n1739), 
        .ZN(n10765) );
  MOAI22 U19687 ( .A1(n27975), .A2(n1738), .B1(ram[6525]), .B2(n1739), 
        .ZN(n10766) );
  MOAI22 U19688 ( .A1(n27740), .A2(n1738), .B1(ram[6526]), .B2(n1739), 
        .ZN(n10767) );
  MOAI22 U19689 ( .A1(n27505), .A2(n1738), .B1(ram[6527]), .B2(n1739), 
        .ZN(n10768) );
  MOAI22 U19690 ( .A1(n29150), .A2(n1740), .B1(ram[6528]), .B2(n1741), 
        .ZN(n10769) );
  MOAI22 U19691 ( .A1(n28915), .A2(n1740), .B1(ram[6529]), .B2(n1741), 
        .ZN(n10770) );
  MOAI22 U19692 ( .A1(n28680), .A2(n1740), .B1(ram[6530]), .B2(n1741), 
        .ZN(n10771) );
  MOAI22 U19693 ( .A1(n28445), .A2(n1740), .B1(ram[6531]), .B2(n1741), 
        .ZN(n10772) );
  MOAI22 U19694 ( .A1(n28210), .A2(n1740), .B1(ram[6532]), .B2(n1741), 
        .ZN(n10773) );
  MOAI22 U19695 ( .A1(n27975), .A2(n1740), .B1(ram[6533]), .B2(n1741), 
        .ZN(n10774) );
  MOAI22 U19696 ( .A1(n27740), .A2(n1740), .B1(ram[6534]), .B2(n1741), 
        .ZN(n10775) );
  MOAI22 U19697 ( .A1(n27505), .A2(n1740), .B1(ram[6535]), .B2(n1741), 
        .ZN(n10776) );
  MOAI22 U19698 ( .A1(n29150), .A2(n1742), .B1(ram[6536]), .B2(n1743), 
        .ZN(n10777) );
  MOAI22 U19699 ( .A1(n28915), .A2(n1742), .B1(ram[6537]), .B2(n1743), 
        .ZN(n10778) );
  MOAI22 U19700 ( .A1(n28680), .A2(n1742), .B1(ram[6538]), .B2(n1743), 
        .ZN(n10779) );
  MOAI22 U19701 ( .A1(n28445), .A2(n1742), .B1(ram[6539]), .B2(n1743), 
        .ZN(n10780) );
  MOAI22 U19702 ( .A1(n28210), .A2(n1742), .B1(ram[6540]), .B2(n1743), 
        .ZN(n10781) );
  MOAI22 U19703 ( .A1(n27975), .A2(n1742), .B1(ram[6541]), .B2(n1743), 
        .ZN(n10782) );
  MOAI22 U19704 ( .A1(n27740), .A2(n1742), .B1(ram[6542]), .B2(n1743), 
        .ZN(n10783) );
  MOAI22 U19705 ( .A1(n27505), .A2(n1742), .B1(ram[6543]), .B2(n1743), 
        .ZN(n10784) );
  MOAI22 U19706 ( .A1(n29150), .A2(n1744), .B1(ram[6544]), .B2(n1745), 
        .ZN(n10785) );
  MOAI22 U19707 ( .A1(n28915), .A2(n1744), .B1(ram[6545]), .B2(n1745), 
        .ZN(n10786) );
  MOAI22 U19708 ( .A1(n28680), .A2(n1744), .B1(ram[6546]), .B2(n1745), 
        .ZN(n10787) );
  MOAI22 U19709 ( .A1(n28445), .A2(n1744), .B1(ram[6547]), .B2(n1745), 
        .ZN(n10788) );
  MOAI22 U19710 ( .A1(n28210), .A2(n1744), .B1(ram[6548]), .B2(n1745), 
        .ZN(n10789) );
  MOAI22 U19711 ( .A1(n27975), .A2(n1744), .B1(ram[6549]), .B2(n1745), 
        .ZN(n10790) );
  MOAI22 U19712 ( .A1(n27740), .A2(n1744), .B1(ram[6550]), .B2(n1745), 
        .ZN(n10791) );
  MOAI22 U19713 ( .A1(n27505), .A2(n1744), .B1(ram[6551]), .B2(n1745), 
        .ZN(n10792) );
  MOAI22 U19714 ( .A1(n29151), .A2(n1746), .B1(ram[6552]), .B2(n1747), 
        .ZN(n10793) );
  MOAI22 U19715 ( .A1(n28916), .A2(n1746), .B1(ram[6553]), .B2(n1747), 
        .ZN(n10794) );
  MOAI22 U19716 ( .A1(n28681), .A2(n1746), .B1(ram[6554]), .B2(n1747), 
        .ZN(n10795) );
  MOAI22 U19717 ( .A1(n28446), .A2(n1746), .B1(ram[6555]), .B2(n1747), 
        .ZN(n10796) );
  MOAI22 U19718 ( .A1(n28211), .A2(n1746), .B1(ram[6556]), .B2(n1747), 
        .ZN(n10797) );
  MOAI22 U19719 ( .A1(n27976), .A2(n1746), .B1(ram[6557]), .B2(n1747), 
        .ZN(n10798) );
  MOAI22 U19720 ( .A1(n27741), .A2(n1746), .B1(ram[6558]), .B2(n1747), 
        .ZN(n10799) );
  MOAI22 U19721 ( .A1(n27506), .A2(n1746), .B1(ram[6559]), .B2(n1747), 
        .ZN(n10800) );
  MOAI22 U19722 ( .A1(n29151), .A2(n1748), .B1(ram[6560]), .B2(n1749), 
        .ZN(n10801) );
  MOAI22 U19723 ( .A1(n28916), .A2(n1748), .B1(ram[6561]), .B2(n1749), 
        .ZN(n10802) );
  MOAI22 U19724 ( .A1(n28681), .A2(n1748), .B1(ram[6562]), .B2(n1749), 
        .ZN(n10803) );
  MOAI22 U19725 ( .A1(n28446), .A2(n1748), .B1(ram[6563]), .B2(n1749), 
        .ZN(n10804) );
  MOAI22 U19726 ( .A1(n28211), .A2(n1748), .B1(ram[6564]), .B2(n1749), 
        .ZN(n10805) );
  MOAI22 U19727 ( .A1(n27976), .A2(n1748), .B1(ram[6565]), .B2(n1749), 
        .ZN(n10806) );
  MOAI22 U19728 ( .A1(n27741), .A2(n1748), .B1(ram[6566]), .B2(n1749), 
        .ZN(n10807) );
  MOAI22 U19729 ( .A1(n27506), .A2(n1748), .B1(ram[6567]), .B2(n1749), 
        .ZN(n10808) );
  MOAI22 U19730 ( .A1(n29151), .A2(n1750), .B1(ram[6568]), .B2(n1751), 
        .ZN(n10809) );
  MOAI22 U19731 ( .A1(n28916), .A2(n1750), .B1(ram[6569]), .B2(n1751), 
        .ZN(n10810) );
  MOAI22 U19732 ( .A1(n28681), .A2(n1750), .B1(ram[6570]), .B2(n1751), 
        .ZN(n10811) );
  MOAI22 U19733 ( .A1(n28446), .A2(n1750), .B1(ram[6571]), .B2(n1751), 
        .ZN(n10812) );
  MOAI22 U19734 ( .A1(n28211), .A2(n1750), .B1(ram[6572]), .B2(n1751), 
        .ZN(n10813) );
  MOAI22 U19735 ( .A1(n27976), .A2(n1750), .B1(ram[6573]), .B2(n1751), 
        .ZN(n10814) );
  MOAI22 U19736 ( .A1(n27741), .A2(n1750), .B1(ram[6574]), .B2(n1751), 
        .ZN(n10815) );
  MOAI22 U19737 ( .A1(n27506), .A2(n1750), .B1(ram[6575]), .B2(n1751), 
        .ZN(n10816) );
  MOAI22 U19738 ( .A1(n29151), .A2(n1752), .B1(ram[6576]), .B2(n1753), 
        .ZN(n10817) );
  MOAI22 U19739 ( .A1(n28916), .A2(n1752), .B1(ram[6577]), .B2(n1753), 
        .ZN(n10818) );
  MOAI22 U19740 ( .A1(n28681), .A2(n1752), .B1(ram[6578]), .B2(n1753), 
        .ZN(n10819) );
  MOAI22 U19741 ( .A1(n28446), .A2(n1752), .B1(ram[6579]), .B2(n1753), 
        .ZN(n10820) );
  MOAI22 U19742 ( .A1(n28211), .A2(n1752), .B1(ram[6580]), .B2(n1753), 
        .ZN(n10821) );
  MOAI22 U19743 ( .A1(n27976), .A2(n1752), .B1(ram[6581]), .B2(n1753), 
        .ZN(n10822) );
  MOAI22 U19744 ( .A1(n27741), .A2(n1752), .B1(ram[6582]), .B2(n1753), 
        .ZN(n10823) );
  MOAI22 U19745 ( .A1(n27506), .A2(n1752), .B1(ram[6583]), .B2(n1753), 
        .ZN(n10824) );
  MOAI22 U19746 ( .A1(n29151), .A2(n1754), .B1(ram[6584]), .B2(n1755), 
        .ZN(n10825) );
  MOAI22 U19747 ( .A1(n28916), .A2(n1754), .B1(ram[6585]), .B2(n1755), 
        .ZN(n10826) );
  MOAI22 U19748 ( .A1(n28681), .A2(n1754), .B1(ram[6586]), .B2(n1755), 
        .ZN(n10827) );
  MOAI22 U19749 ( .A1(n28446), .A2(n1754), .B1(ram[6587]), .B2(n1755), 
        .ZN(n10828) );
  MOAI22 U19750 ( .A1(n28211), .A2(n1754), .B1(ram[6588]), .B2(n1755), 
        .ZN(n10829) );
  MOAI22 U19751 ( .A1(n27976), .A2(n1754), .B1(ram[6589]), .B2(n1755), 
        .ZN(n10830) );
  MOAI22 U19752 ( .A1(n27741), .A2(n1754), .B1(ram[6590]), .B2(n1755), 
        .ZN(n10831) );
  MOAI22 U19753 ( .A1(n27506), .A2(n1754), .B1(ram[6591]), .B2(n1755), 
        .ZN(n10832) );
  MOAI22 U19754 ( .A1(n29151), .A2(n1756), .B1(ram[6592]), .B2(n1757), 
        .ZN(n10833) );
  MOAI22 U19755 ( .A1(n28916), .A2(n1756), .B1(ram[6593]), .B2(n1757), 
        .ZN(n10834) );
  MOAI22 U19756 ( .A1(n28681), .A2(n1756), .B1(ram[6594]), .B2(n1757), 
        .ZN(n10835) );
  MOAI22 U19757 ( .A1(n28446), .A2(n1756), .B1(ram[6595]), .B2(n1757), 
        .ZN(n10836) );
  MOAI22 U19758 ( .A1(n28211), .A2(n1756), .B1(ram[6596]), .B2(n1757), 
        .ZN(n10837) );
  MOAI22 U19759 ( .A1(n27976), .A2(n1756), .B1(ram[6597]), .B2(n1757), 
        .ZN(n10838) );
  MOAI22 U19760 ( .A1(n27741), .A2(n1756), .B1(ram[6598]), .B2(n1757), 
        .ZN(n10839) );
  MOAI22 U19761 ( .A1(n27506), .A2(n1756), .B1(ram[6599]), .B2(n1757), 
        .ZN(n10840) );
  MOAI22 U19762 ( .A1(n29151), .A2(n1758), .B1(ram[6600]), .B2(n1759), 
        .ZN(n10841) );
  MOAI22 U19763 ( .A1(n28916), .A2(n1758), .B1(ram[6601]), .B2(n1759), 
        .ZN(n10842) );
  MOAI22 U19764 ( .A1(n28681), .A2(n1758), .B1(ram[6602]), .B2(n1759), 
        .ZN(n10843) );
  MOAI22 U19765 ( .A1(n28446), .A2(n1758), .B1(ram[6603]), .B2(n1759), 
        .ZN(n10844) );
  MOAI22 U19766 ( .A1(n28211), .A2(n1758), .B1(ram[6604]), .B2(n1759), 
        .ZN(n10845) );
  MOAI22 U19767 ( .A1(n27976), .A2(n1758), .B1(ram[6605]), .B2(n1759), 
        .ZN(n10846) );
  MOAI22 U19768 ( .A1(n27741), .A2(n1758), .B1(ram[6606]), .B2(n1759), 
        .ZN(n10847) );
  MOAI22 U19769 ( .A1(n27506), .A2(n1758), .B1(ram[6607]), .B2(n1759), 
        .ZN(n10848) );
  MOAI22 U19770 ( .A1(n29151), .A2(n1760), .B1(ram[6608]), .B2(n1761), 
        .ZN(n10849) );
  MOAI22 U19771 ( .A1(n28916), .A2(n1760), .B1(ram[6609]), .B2(n1761), 
        .ZN(n10850) );
  MOAI22 U19772 ( .A1(n28681), .A2(n1760), .B1(ram[6610]), .B2(n1761), 
        .ZN(n10851) );
  MOAI22 U19773 ( .A1(n28446), .A2(n1760), .B1(ram[6611]), .B2(n1761), 
        .ZN(n10852) );
  MOAI22 U19774 ( .A1(n28211), .A2(n1760), .B1(ram[6612]), .B2(n1761), 
        .ZN(n10853) );
  MOAI22 U19775 ( .A1(n27976), .A2(n1760), .B1(ram[6613]), .B2(n1761), 
        .ZN(n10854) );
  MOAI22 U19776 ( .A1(n27741), .A2(n1760), .B1(ram[6614]), .B2(n1761), 
        .ZN(n10855) );
  MOAI22 U19777 ( .A1(n27506), .A2(n1760), .B1(ram[6615]), .B2(n1761), 
        .ZN(n10856) );
  MOAI22 U19778 ( .A1(n29151), .A2(n1762), .B1(ram[6616]), .B2(n1763), 
        .ZN(n10857) );
  MOAI22 U19779 ( .A1(n28916), .A2(n1762), .B1(ram[6617]), .B2(n1763), 
        .ZN(n10858) );
  MOAI22 U19780 ( .A1(n28681), .A2(n1762), .B1(ram[6618]), .B2(n1763), 
        .ZN(n10859) );
  MOAI22 U19781 ( .A1(n28446), .A2(n1762), .B1(ram[6619]), .B2(n1763), 
        .ZN(n10860) );
  MOAI22 U19782 ( .A1(n28211), .A2(n1762), .B1(ram[6620]), .B2(n1763), 
        .ZN(n10861) );
  MOAI22 U19783 ( .A1(n27976), .A2(n1762), .B1(ram[6621]), .B2(n1763), 
        .ZN(n10862) );
  MOAI22 U19784 ( .A1(n27741), .A2(n1762), .B1(ram[6622]), .B2(n1763), 
        .ZN(n10863) );
  MOAI22 U19785 ( .A1(n27506), .A2(n1762), .B1(ram[6623]), .B2(n1763), 
        .ZN(n10864) );
  MOAI22 U19786 ( .A1(n29151), .A2(n1764), .B1(ram[6624]), .B2(n1765), 
        .ZN(n10865) );
  MOAI22 U19787 ( .A1(n28916), .A2(n1764), .B1(ram[6625]), .B2(n1765), 
        .ZN(n10866) );
  MOAI22 U19788 ( .A1(n28681), .A2(n1764), .B1(ram[6626]), .B2(n1765), 
        .ZN(n10867) );
  MOAI22 U19789 ( .A1(n28446), .A2(n1764), .B1(ram[6627]), .B2(n1765), 
        .ZN(n10868) );
  MOAI22 U19790 ( .A1(n28211), .A2(n1764), .B1(ram[6628]), .B2(n1765), 
        .ZN(n10869) );
  MOAI22 U19791 ( .A1(n27976), .A2(n1764), .B1(ram[6629]), .B2(n1765), 
        .ZN(n10870) );
  MOAI22 U19792 ( .A1(n27741), .A2(n1764), .B1(ram[6630]), .B2(n1765), 
        .ZN(n10871) );
  MOAI22 U19793 ( .A1(n27506), .A2(n1764), .B1(ram[6631]), .B2(n1765), 
        .ZN(n10872) );
  MOAI22 U19794 ( .A1(n29151), .A2(n1766), .B1(ram[6632]), .B2(n1767), 
        .ZN(n10873) );
  MOAI22 U19795 ( .A1(n28916), .A2(n1766), .B1(ram[6633]), .B2(n1767), 
        .ZN(n10874) );
  MOAI22 U19796 ( .A1(n28681), .A2(n1766), .B1(ram[6634]), .B2(n1767), 
        .ZN(n10875) );
  MOAI22 U19797 ( .A1(n28446), .A2(n1766), .B1(ram[6635]), .B2(n1767), 
        .ZN(n10876) );
  MOAI22 U19798 ( .A1(n28211), .A2(n1766), .B1(ram[6636]), .B2(n1767), 
        .ZN(n10877) );
  MOAI22 U19799 ( .A1(n27976), .A2(n1766), .B1(ram[6637]), .B2(n1767), 
        .ZN(n10878) );
  MOAI22 U19800 ( .A1(n27741), .A2(n1766), .B1(ram[6638]), .B2(n1767), 
        .ZN(n10879) );
  MOAI22 U19801 ( .A1(n27506), .A2(n1766), .B1(ram[6639]), .B2(n1767), 
        .ZN(n10880) );
  MOAI22 U19802 ( .A1(n29151), .A2(n1768), .B1(ram[6640]), .B2(n1769), 
        .ZN(n10881) );
  MOAI22 U19803 ( .A1(n28916), .A2(n1768), .B1(ram[6641]), .B2(n1769), 
        .ZN(n10882) );
  MOAI22 U19804 ( .A1(n28681), .A2(n1768), .B1(ram[6642]), .B2(n1769), 
        .ZN(n10883) );
  MOAI22 U19805 ( .A1(n28446), .A2(n1768), .B1(ram[6643]), .B2(n1769), 
        .ZN(n10884) );
  MOAI22 U19806 ( .A1(n28211), .A2(n1768), .B1(ram[6644]), .B2(n1769), 
        .ZN(n10885) );
  MOAI22 U19807 ( .A1(n27976), .A2(n1768), .B1(ram[6645]), .B2(n1769), 
        .ZN(n10886) );
  MOAI22 U19808 ( .A1(n27741), .A2(n1768), .B1(ram[6646]), .B2(n1769), 
        .ZN(n10887) );
  MOAI22 U19809 ( .A1(n27506), .A2(n1768), .B1(ram[6647]), .B2(n1769), 
        .ZN(n10888) );
  MOAI22 U19810 ( .A1(n29151), .A2(n1770), .B1(ram[6648]), .B2(n1771), 
        .ZN(n10889) );
  MOAI22 U19811 ( .A1(n28916), .A2(n1770), .B1(ram[6649]), .B2(n1771), 
        .ZN(n10890) );
  MOAI22 U19812 ( .A1(n28681), .A2(n1770), .B1(ram[6650]), .B2(n1771), 
        .ZN(n10891) );
  MOAI22 U19813 ( .A1(n28446), .A2(n1770), .B1(ram[6651]), .B2(n1771), 
        .ZN(n10892) );
  MOAI22 U19814 ( .A1(n28211), .A2(n1770), .B1(ram[6652]), .B2(n1771), 
        .ZN(n10893) );
  MOAI22 U19815 ( .A1(n27976), .A2(n1770), .B1(ram[6653]), .B2(n1771), 
        .ZN(n10894) );
  MOAI22 U19816 ( .A1(n27741), .A2(n1770), .B1(ram[6654]), .B2(n1771), 
        .ZN(n10895) );
  MOAI22 U19817 ( .A1(n27506), .A2(n1770), .B1(ram[6655]), .B2(n1771), 
        .ZN(n10896) );
  MOAI22 U19818 ( .A1(n29152), .A2(n1772), .B1(ram[6656]), .B2(n1773), 
        .ZN(n10897) );
  MOAI22 U19819 ( .A1(n28917), .A2(n1772), .B1(ram[6657]), .B2(n1773), 
        .ZN(n10898) );
  MOAI22 U19820 ( .A1(n28682), .A2(n1772), .B1(ram[6658]), .B2(n1773), 
        .ZN(n10899) );
  MOAI22 U19821 ( .A1(n28447), .A2(n1772), .B1(ram[6659]), .B2(n1773), 
        .ZN(n10900) );
  MOAI22 U19822 ( .A1(n28212), .A2(n1772), .B1(ram[6660]), .B2(n1773), 
        .ZN(n10901) );
  MOAI22 U19823 ( .A1(n27977), .A2(n1772), .B1(ram[6661]), .B2(n1773), 
        .ZN(n10902) );
  MOAI22 U19824 ( .A1(n27742), .A2(n1772), .B1(ram[6662]), .B2(n1773), 
        .ZN(n10903) );
  MOAI22 U19825 ( .A1(n27507), .A2(n1772), .B1(ram[6663]), .B2(n1773), 
        .ZN(n10904) );
  MOAI22 U19826 ( .A1(n29152), .A2(n1775), .B1(ram[6664]), .B2(n1776), 
        .ZN(n10905) );
  MOAI22 U19827 ( .A1(n28917), .A2(n1775), .B1(ram[6665]), .B2(n1776), 
        .ZN(n10906) );
  MOAI22 U19828 ( .A1(n28682), .A2(n1775), .B1(ram[6666]), .B2(n1776), 
        .ZN(n10907) );
  MOAI22 U19829 ( .A1(n28447), .A2(n1775), .B1(ram[6667]), .B2(n1776), 
        .ZN(n10908) );
  MOAI22 U19830 ( .A1(n28212), .A2(n1775), .B1(ram[6668]), .B2(n1776), 
        .ZN(n10909) );
  MOAI22 U19831 ( .A1(n27977), .A2(n1775), .B1(ram[6669]), .B2(n1776), 
        .ZN(n10910) );
  MOAI22 U19832 ( .A1(n27742), .A2(n1775), .B1(ram[6670]), .B2(n1776), 
        .ZN(n10911) );
  MOAI22 U19833 ( .A1(n27507), .A2(n1775), .B1(ram[6671]), .B2(n1776), 
        .ZN(n10912) );
  MOAI22 U19834 ( .A1(n29152), .A2(n1777), .B1(ram[6672]), .B2(n1778), 
        .ZN(n10913) );
  MOAI22 U19835 ( .A1(n28917), .A2(n1777), .B1(ram[6673]), .B2(n1778), 
        .ZN(n10914) );
  MOAI22 U19836 ( .A1(n28682), .A2(n1777), .B1(ram[6674]), .B2(n1778), 
        .ZN(n10915) );
  MOAI22 U19837 ( .A1(n28447), .A2(n1777), .B1(ram[6675]), .B2(n1778), 
        .ZN(n10916) );
  MOAI22 U19838 ( .A1(n28212), .A2(n1777), .B1(ram[6676]), .B2(n1778), 
        .ZN(n10917) );
  MOAI22 U19839 ( .A1(n27977), .A2(n1777), .B1(ram[6677]), .B2(n1778), 
        .ZN(n10918) );
  MOAI22 U19840 ( .A1(n27742), .A2(n1777), .B1(ram[6678]), .B2(n1778), 
        .ZN(n10919) );
  MOAI22 U19841 ( .A1(n27507), .A2(n1777), .B1(ram[6679]), .B2(n1778), 
        .ZN(n10920) );
  MOAI22 U19842 ( .A1(n29152), .A2(n1779), .B1(ram[6680]), .B2(n1780), 
        .ZN(n10921) );
  MOAI22 U19843 ( .A1(n28917), .A2(n1779), .B1(ram[6681]), .B2(n1780), 
        .ZN(n10922) );
  MOAI22 U19844 ( .A1(n28682), .A2(n1779), .B1(ram[6682]), .B2(n1780), 
        .ZN(n10923) );
  MOAI22 U19845 ( .A1(n28447), .A2(n1779), .B1(ram[6683]), .B2(n1780), 
        .ZN(n10924) );
  MOAI22 U19846 ( .A1(n28212), .A2(n1779), .B1(ram[6684]), .B2(n1780), 
        .ZN(n10925) );
  MOAI22 U19847 ( .A1(n27977), .A2(n1779), .B1(ram[6685]), .B2(n1780), 
        .ZN(n10926) );
  MOAI22 U19848 ( .A1(n27742), .A2(n1779), .B1(ram[6686]), .B2(n1780), 
        .ZN(n10927) );
  MOAI22 U19849 ( .A1(n27507), .A2(n1779), .B1(ram[6687]), .B2(n1780), 
        .ZN(n10928) );
  MOAI22 U19850 ( .A1(n29152), .A2(n1781), .B1(ram[6688]), .B2(n1782), 
        .ZN(n10929) );
  MOAI22 U19851 ( .A1(n28917), .A2(n1781), .B1(ram[6689]), .B2(n1782), 
        .ZN(n10930) );
  MOAI22 U19852 ( .A1(n28682), .A2(n1781), .B1(ram[6690]), .B2(n1782), 
        .ZN(n10931) );
  MOAI22 U19853 ( .A1(n28447), .A2(n1781), .B1(ram[6691]), .B2(n1782), 
        .ZN(n10932) );
  MOAI22 U19854 ( .A1(n28212), .A2(n1781), .B1(ram[6692]), .B2(n1782), 
        .ZN(n10933) );
  MOAI22 U19855 ( .A1(n27977), .A2(n1781), .B1(ram[6693]), .B2(n1782), 
        .ZN(n10934) );
  MOAI22 U19856 ( .A1(n27742), .A2(n1781), .B1(ram[6694]), .B2(n1782), 
        .ZN(n10935) );
  MOAI22 U19857 ( .A1(n27507), .A2(n1781), .B1(ram[6695]), .B2(n1782), 
        .ZN(n10936) );
  MOAI22 U19858 ( .A1(n29152), .A2(n1783), .B1(ram[6696]), .B2(n1784), 
        .ZN(n10937) );
  MOAI22 U19859 ( .A1(n28917), .A2(n1783), .B1(ram[6697]), .B2(n1784), 
        .ZN(n10938) );
  MOAI22 U19860 ( .A1(n28682), .A2(n1783), .B1(ram[6698]), .B2(n1784), 
        .ZN(n10939) );
  MOAI22 U19861 ( .A1(n28447), .A2(n1783), .B1(ram[6699]), .B2(n1784), 
        .ZN(n10940) );
  MOAI22 U19862 ( .A1(n28212), .A2(n1783), .B1(ram[6700]), .B2(n1784), 
        .ZN(n10941) );
  MOAI22 U19863 ( .A1(n27977), .A2(n1783), .B1(ram[6701]), .B2(n1784), 
        .ZN(n10942) );
  MOAI22 U19864 ( .A1(n27742), .A2(n1783), .B1(ram[6702]), .B2(n1784), 
        .ZN(n10943) );
  MOAI22 U19865 ( .A1(n27507), .A2(n1783), .B1(ram[6703]), .B2(n1784), 
        .ZN(n10944) );
  MOAI22 U19866 ( .A1(n29152), .A2(n1785), .B1(ram[6704]), .B2(n1786), 
        .ZN(n10945) );
  MOAI22 U19867 ( .A1(n28917), .A2(n1785), .B1(ram[6705]), .B2(n1786), 
        .ZN(n10946) );
  MOAI22 U19868 ( .A1(n28682), .A2(n1785), .B1(ram[6706]), .B2(n1786), 
        .ZN(n10947) );
  MOAI22 U19869 ( .A1(n28447), .A2(n1785), .B1(ram[6707]), .B2(n1786), 
        .ZN(n10948) );
  MOAI22 U19870 ( .A1(n28212), .A2(n1785), .B1(ram[6708]), .B2(n1786), 
        .ZN(n10949) );
  MOAI22 U19871 ( .A1(n27977), .A2(n1785), .B1(ram[6709]), .B2(n1786), 
        .ZN(n10950) );
  MOAI22 U19872 ( .A1(n27742), .A2(n1785), .B1(ram[6710]), .B2(n1786), 
        .ZN(n10951) );
  MOAI22 U19873 ( .A1(n27507), .A2(n1785), .B1(ram[6711]), .B2(n1786), 
        .ZN(n10952) );
  MOAI22 U19874 ( .A1(n29152), .A2(n1787), .B1(ram[6712]), .B2(n1788), 
        .ZN(n10953) );
  MOAI22 U19875 ( .A1(n28917), .A2(n1787), .B1(ram[6713]), .B2(n1788), 
        .ZN(n10954) );
  MOAI22 U19876 ( .A1(n28682), .A2(n1787), .B1(ram[6714]), .B2(n1788), 
        .ZN(n10955) );
  MOAI22 U19877 ( .A1(n28447), .A2(n1787), .B1(ram[6715]), .B2(n1788), 
        .ZN(n10956) );
  MOAI22 U19878 ( .A1(n28212), .A2(n1787), .B1(ram[6716]), .B2(n1788), 
        .ZN(n10957) );
  MOAI22 U19879 ( .A1(n27977), .A2(n1787), .B1(ram[6717]), .B2(n1788), 
        .ZN(n10958) );
  MOAI22 U19880 ( .A1(n27742), .A2(n1787), .B1(ram[6718]), .B2(n1788), 
        .ZN(n10959) );
  MOAI22 U19881 ( .A1(n27507), .A2(n1787), .B1(ram[6719]), .B2(n1788), 
        .ZN(n10960) );
  MOAI22 U19882 ( .A1(n29152), .A2(n1789), .B1(ram[6720]), .B2(n1790), 
        .ZN(n10961) );
  MOAI22 U19883 ( .A1(n28917), .A2(n1789), .B1(ram[6721]), .B2(n1790), 
        .ZN(n10962) );
  MOAI22 U19884 ( .A1(n28682), .A2(n1789), .B1(ram[6722]), .B2(n1790), 
        .ZN(n10963) );
  MOAI22 U19885 ( .A1(n28447), .A2(n1789), .B1(ram[6723]), .B2(n1790), 
        .ZN(n10964) );
  MOAI22 U19886 ( .A1(n28212), .A2(n1789), .B1(ram[6724]), .B2(n1790), 
        .ZN(n10965) );
  MOAI22 U19887 ( .A1(n27977), .A2(n1789), .B1(ram[6725]), .B2(n1790), 
        .ZN(n10966) );
  MOAI22 U19888 ( .A1(n27742), .A2(n1789), .B1(ram[6726]), .B2(n1790), 
        .ZN(n10967) );
  MOAI22 U19889 ( .A1(n27507), .A2(n1789), .B1(ram[6727]), .B2(n1790), 
        .ZN(n10968) );
  MOAI22 U19890 ( .A1(n29152), .A2(n1791), .B1(ram[6728]), .B2(n1792), 
        .ZN(n10969) );
  MOAI22 U19891 ( .A1(n28917), .A2(n1791), .B1(ram[6729]), .B2(n1792), 
        .ZN(n10970) );
  MOAI22 U19892 ( .A1(n28682), .A2(n1791), .B1(ram[6730]), .B2(n1792), 
        .ZN(n10971) );
  MOAI22 U19893 ( .A1(n28447), .A2(n1791), .B1(ram[6731]), .B2(n1792), 
        .ZN(n10972) );
  MOAI22 U19894 ( .A1(n28212), .A2(n1791), .B1(ram[6732]), .B2(n1792), 
        .ZN(n10973) );
  MOAI22 U19895 ( .A1(n27977), .A2(n1791), .B1(ram[6733]), .B2(n1792), 
        .ZN(n10974) );
  MOAI22 U19896 ( .A1(n27742), .A2(n1791), .B1(ram[6734]), .B2(n1792), 
        .ZN(n10975) );
  MOAI22 U19897 ( .A1(n27507), .A2(n1791), .B1(ram[6735]), .B2(n1792), 
        .ZN(n10976) );
  MOAI22 U19898 ( .A1(n29152), .A2(n1793), .B1(ram[6736]), .B2(n1794), 
        .ZN(n10977) );
  MOAI22 U19899 ( .A1(n28917), .A2(n1793), .B1(ram[6737]), .B2(n1794), 
        .ZN(n10978) );
  MOAI22 U19900 ( .A1(n28682), .A2(n1793), .B1(ram[6738]), .B2(n1794), 
        .ZN(n10979) );
  MOAI22 U19901 ( .A1(n28447), .A2(n1793), .B1(ram[6739]), .B2(n1794), 
        .ZN(n10980) );
  MOAI22 U19902 ( .A1(n28212), .A2(n1793), .B1(ram[6740]), .B2(n1794), 
        .ZN(n10981) );
  MOAI22 U19903 ( .A1(n27977), .A2(n1793), .B1(ram[6741]), .B2(n1794), 
        .ZN(n10982) );
  MOAI22 U19904 ( .A1(n27742), .A2(n1793), .B1(ram[6742]), .B2(n1794), 
        .ZN(n10983) );
  MOAI22 U19905 ( .A1(n27507), .A2(n1793), .B1(ram[6743]), .B2(n1794), 
        .ZN(n10984) );
  MOAI22 U19906 ( .A1(n29152), .A2(n1795), .B1(ram[6744]), .B2(n1796), 
        .ZN(n10985) );
  MOAI22 U19907 ( .A1(n28917), .A2(n1795), .B1(ram[6745]), .B2(n1796), 
        .ZN(n10986) );
  MOAI22 U19908 ( .A1(n28682), .A2(n1795), .B1(ram[6746]), .B2(n1796), 
        .ZN(n10987) );
  MOAI22 U19909 ( .A1(n28447), .A2(n1795), .B1(ram[6747]), .B2(n1796), 
        .ZN(n10988) );
  MOAI22 U19910 ( .A1(n28212), .A2(n1795), .B1(ram[6748]), .B2(n1796), 
        .ZN(n10989) );
  MOAI22 U19911 ( .A1(n27977), .A2(n1795), .B1(ram[6749]), .B2(n1796), 
        .ZN(n10990) );
  MOAI22 U19912 ( .A1(n27742), .A2(n1795), .B1(ram[6750]), .B2(n1796), 
        .ZN(n10991) );
  MOAI22 U19913 ( .A1(n27507), .A2(n1795), .B1(ram[6751]), .B2(n1796), 
        .ZN(n10992) );
  MOAI22 U19914 ( .A1(n29152), .A2(n1797), .B1(ram[6752]), .B2(n1798), 
        .ZN(n10993) );
  MOAI22 U19915 ( .A1(n28917), .A2(n1797), .B1(ram[6753]), .B2(n1798), 
        .ZN(n10994) );
  MOAI22 U19916 ( .A1(n28682), .A2(n1797), .B1(ram[6754]), .B2(n1798), 
        .ZN(n10995) );
  MOAI22 U19917 ( .A1(n28447), .A2(n1797), .B1(ram[6755]), .B2(n1798), 
        .ZN(n10996) );
  MOAI22 U19918 ( .A1(n28212), .A2(n1797), .B1(ram[6756]), .B2(n1798), 
        .ZN(n10997) );
  MOAI22 U19919 ( .A1(n27977), .A2(n1797), .B1(ram[6757]), .B2(n1798), 
        .ZN(n10998) );
  MOAI22 U19920 ( .A1(n27742), .A2(n1797), .B1(ram[6758]), .B2(n1798), 
        .ZN(n10999) );
  MOAI22 U19921 ( .A1(n27507), .A2(n1797), .B1(ram[6759]), .B2(n1798), 
        .ZN(n11000) );
  MOAI22 U19922 ( .A1(n29153), .A2(n1799), .B1(ram[6760]), .B2(n1800), 
        .ZN(n11001) );
  MOAI22 U19923 ( .A1(n28918), .A2(n1799), .B1(ram[6761]), .B2(n1800), 
        .ZN(n11002) );
  MOAI22 U19924 ( .A1(n28683), .A2(n1799), .B1(ram[6762]), .B2(n1800), 
        .ZN(n11003) );
  MOAI22 U19925 ( .A1(n28448), .A2(n1799), .B1(ram[6763]), .B2(n1800), 
        .ZN(n11004) );
  MOAI22 U19926 ( .A1(n28213), .A2(n1799), .B1(ram[6764]), .B2(n1800), 
        .ZN(n11005) );
  MOAI22 U19927 ( .A1(n27978), .A2(n1799), .B1(ram[6765]), .B2(n1800), 
        .ZN(n11006) );
  MOAI22 U19928 ( .A1(n27743), .A2(n1799), .B1(ram[6766]), .B2(n1800), 
        .ZN(n11007) );
  MOAI22 U19929 ( .A1(n27508), .A2(n1799), .B1(ram[6767]), .B2(n1800), 
        .ZN(n11008) );
  MOAI22 U19930 ( .A1(n29153), .A2(n1801), .B1(ram[6768]), .B2(n1802), 
        .ZN(n11009) );
  MOAI22 U19931 ( .A1(n28918), .A2(n1801), .B1(ram[6769]), .B2(n1802), 
        .ZN(n11010) );
  MOAI22 U19932 ( .A1(n28683), .A2(n1801), .B1(ram[6770]), .B2(n1802), 
        .ZN(n11011) );
  MOAI22 U19933 ( .A1(n28448), .A2(n1801), .B1(ram[6771]), .B2(n1802), 
        .ZN(n11012) );
  MOAI22 U19934 ( .A1(n28213), .A2(n1801), .B1(ram[6772]), .B2(n1802), 
        .ZN(n11013) );
  MOAI22 U19935 ( .A1(n27978), .A2(n1801), .B1(ram[6773]), .B2(n1802), 
        .ZN(n11014) );
  MOAI22 U19936 ( .A1(n27743), .A2(n1801), .B1(ram[6774]), .B2(n1802), 
        .ZN(n11015) );
  MOAI22 U19937 ( .A1(n27508), .A2(n1801), .B1(ram[6775]), .B2(n1802), 
        .ZN(n11016) );
  MOAI22 U19938 ( .A1(n29153), .A2(n1803), .B1(ram[6776]), .B2(n1804), 
        .ZN(n11017) );
  MOAI22 U19939 ( .A1(n28918), .A2(n1803), .B1(ram[6777]), .B2(n1804), 
        .ZN(n11018) );
  MOAI22 U19940 ( .A1(n28683), .A2(n1803), .B1(ram[6778]), .B2(n1804), 
        .ZN(n11019) );
  MOAI22 U19941 ( .A1(n28448), .A2(n1803), .B1(ram[6779]), .B2(n1804), 
        .ZN(n11020) );
  MOAI22 U19942 ( .A1(n28213), .A2(n1803), .B1(ram[6780]), .B2(n1804), 
        .ZN(n11021) );
  MOAI22 U19943 ( .A1(n27978), .A2(n1803), .B1(ram[6781]), .B2(n1804), 
        .ZN(n11022) );
  MOAI22 U19944 ( .A1(n27743), .A2(n1803), .B1(ram[6782]), .B2(n1804), 
        .ZN(n11023) );
  MOAI22 U19945 ( .A1(n27508), .A2(n1803), .B1(ram[6783]), .B2(n1804), 
        .ZN(n11024) );
  MOAI22 U19946 ( .A1(n29153), .A2(n1805), .B1(ram[6784]), .B2(n1806), 
        .ZN(n11025) );
  MOAI22 U19947 ( .A1(n28918), .A2(n1805), .B1(ram[6785]), .B2(n1806), 
        .ZN(n11026) );
  MOAI22 U19948 ( .A1(n28683), .A2(n1805), .B1(ram[6786]), .B2(n1806), 
        .ZN(n11027) );
  MOAI22 U19949 ( .A1(n28448), .A2(n1805), .B1(ram[6787]), .B2(n1806), 
        .ZN(n11028) );
  MOAI22 U19950 ( .A1(n28213), .A2(n1805), .B1(ram[6788]), .B2(n1806), 
        .ZN(n11029) );
  MOAI22 U19951 ( .A1(n27978), .A2(n1805), .B1(ram[6789]), .B2(n1806), 
        .ZN(n11030) );
  MOAI22 U19952 ( .A1(n27743), .A2(n1805), .B1(ram[6790]), .B2(n1806), 
        .ZN(n11031) );
  MOAI22 U19953 ( .A1(n27508), .A2(n1805), .B1(ram[6791]), .B2(n1806), 
        .ZN(n11032) );
  MOAI22 U19954 ( .A1(n29153), .A2(n1807), .B1(ram[6792]), .B2(n1808), 
        .ZN(n11033) );
  MOAI22 U19955 ( .A1(n28918), .A2(n1807), .B1(ram[6793]), .B2(n1808), 
        .ZN(n11034) );
  MOAI22 U19956 ( .A1(n28683), .A2(n1807), .B1(ram[6794]), .B2(n1808), 
        .ZN(n11035) );
  MOAI22 U19957 ( .A1(n28448), .A2(n1807), .B1(ram[6795]), .B2(n1808), 
        .ZN(n11036) );
  MOAI22 U19958 ( .A1(n28213), .A2(n1807), .B1(ram[6796]), .B2(n1808), 
        .ZN(n11037) );
  MOAI22 U19959 ( .A1(n27978), .A2(n1807), .B1(ram[6797]), .B2(n1808), 
        .ZN(n11038) );
  MOAI22 U19960 ( .A1(n27743), .A2(n1807), .B1(ram[6798]), .B2(n1808), 
        .ZN(n11039) );
  MOAI22 U19961 ( .A1(n27508), .A2(n1807), .B1(ram[6799]), .B2(n1808), 
        .ZN(n11040) );
  MOAI22 U19962 ( .A1(n29153), .A2(n1809), .B1(ram[6800]), .B2(n1810), 
        .ZN(n11041) );
  MOAI22 U19963 ( .A1(n28918), .A2(n1809), .B1(ram[6801]), .B2(n1810), 
        .ZN(n11042) );
  MOAI22 U19964 ( .A1(n28683), .A2(n1809), .B1(ram[6802]), .B2(n1810), 
        .ZN(n11043) );
  MOAI22 U19965 ( .A1(n28448), .A2(n1809), .B1(ram[6803]), .B2(n1810), 
        .ZN(n11044) );
  MOAI22 U19966 ( .A1(n28213), .A2(n1809), .B1(ram[6804]), .B2(n1810), 
        .ZN(n11045) );
  MOAI22 U19967 ( .A1(n27978), .A2(n1809), .B1(ram[6805]), .B2(n1810), 
        .ZN(n11046) );
  MOAI22 U19968 ( .A1(n27743), .A2(n1809), .B1(ram[6806]), .B2(n1810), 
        .ZN(n11047) );
  MOAI22 U19969 ( .A1(n27508), .A2(n1809), .B1(ram[6807]), .B2(n1810), 
        .ZN(n11048) );
  MOAI22 U19970 ( .A1(n29153), .A2(n1811), .B1(ram[6808]), .B2(n1812), 
        .ZN(n11049) );
  MOAI22 U19971 ( .A1(n28918), .A2(n1811), .B1(ram[6809]), .B2(n1812), 
        .ZN(n11050) );
  MOAI22 U19972 ( .A1(n28683), .A2(n1811), .B1(ram[6810]), .B2(n1812), 
        .ZN(n11051) );
  MOAI22 U19973 ( .A1(n28448), .A2(n1811), .B1(ram[6811]), .B2(n1812), 
        .ZN(n11052) );
  MOAI22 U19974 ( .A1(n28213), .A2(n1811), .B1(ram[6812]), .B2(n1812), 
        .ZN(n11053) );
  MOAI22 U19975 ( .A1(n27978), .A2(n1811), .B1(ram[6813]), .B2(n1812), 
        .ZN(n11054) );
  MOAI22 U19976 ( .A1(n27743), .A2(n1811), .B1(ram[6814]), .B2(n1812), 
        .ZN(n11055) );
  MOAI22 U19977 ( .A1(n27508), .A2(n1811), .B1(ram[6815]), .B2(n1812), 
        .ZN(n11056) );
  MOAI22 U19978 ( .A1(n29153), .A2(n1813), .B1(ram[6816]), .B2(n1814), 
        .ZN(n11057) );
  MOAI22 U19979 ( .A1(n28918), .A2(n1813), .B1(ram[6817]), .B2(n1814), 
        .ZN(n11058) );
  MOAI22 U19980 ( .A1(n28683), .A2(n1813), .B1(ram[6818]), .B2(n1814), 
        .ZN(n11059) );
  MOAI22 U19981 ( .A1(n28448), .A2(n1813), .B1(ram[6819]), .B2(n1814), 
        .ZN(n11060) );
  MOAI22 U19982 ( .A1(n28213), .A2(n1813), .B1(ram[6820]), .B2(n1814), 
        .ZN(n11061) );
  MOAI22 U19983 ( .A1(n27978), .A2(n1813), .B1(ram[6821]), .B2(n1814), 
        .ZN(n11062) );
  MOAI22 U19984 ( .A1(n27743), .A2(n1813), .B1(ram[6822]), .B2(n1814), 
        .ZN(n11063) );
  MOAI22 U19985 ( .A1(n27508), .A2(n1813), .B1(ram[6823]), .B2(n1814), 
        .ZN(n11064) );
  MOAI22 U19986 ( .A1(n29153), .A2(n1815), .B1(ram[6824]), .B2(n1816), 
        .ZN(n11065) );
  MOAI22 U19987 ( .A1(n28918), .A2(n1815), .B1(ram[6825]), .B2(n1816), 
        .ZN(n11066) );
  MOAI22 U19988 ( .A1(n28683), .A2(n1815), .B1(ram[6826]), .B2(n1816), 
        .ZN(n11067) );
  MOAI22 U19989 ( .A1(n28448), .A2(n1815), .B1(ram[6827]), .B2(n1816), 
        .ZN(n11068) );
  MOAI22 U19990 ( .A1(n28213), .A2(n1815), .B1(ram[6828]), .B2(n1816), 
        .ZN(n11069) );
  MOAI22 U19991 ( .A1(n27978), .A2(n1815), .B1(ram[6829]), .B2(n1816), 
        .ZN(n11070) );
  MOAI22 U19992 ( .A1(n27743), .A2(n1815), .B1(ram[6830]), .B2(n1816), 
        .ZN(n11071) );
  MOAI22 U19993 ( .A1(n27508), .A2(n1815), .B1(ram[6831]), .B2(n1816), 
        .ZN(n11072) );
  MOAI22 U19994 ( .A1(n29153), .A2(n1817), .B1(ram[6832]), .B2(n1818), 
        .ZN(n11073) );
  MOAI22 U19995 ( .A1(n28918), .A2(n1817), .B1(ram[6833]), .B2(n1818), 
        .ZN(n11074) );
  MOAI22 U19996 ( .A1(n28683), .A2(n1817), .B1(ram[6834]), .B2(n1818), 
        .ZN(n11075) );
  MOAI22 U19997 ( .A1(n28448), .A2(n1817), .B1(ram[6835]), .B2(n1818), 
        .ZN(n11076) );
  MOAI22 U19998 ( .A1(n28213), .A2(n1817), .B1(ram[6836]), .B2(n1818), 
        .ZN(n11077) );
  MOAI22 U19999 ( .A1(n27978), .A2(n1817), .B1(ram[6837]), .B2(n1818), 
        .ZN(n11078) );
  MOAI22 U20000 ( .A1(n27743), .A2(n1817), .B1(ram[6838]), .B2(n1818), 
        .ZN(n11079) );
  MOAI22 U20001 ( .A1(n27508), .A2(n1817), .B1(ram[6839]), .B2(n1818), 
        .ZN(n11080) );
  MOAI22 U20002 ( .A1(n29153), .A2(n1819), .B1(ram[6840]), .B2(n1820), 
        .ZN(n11081) );
  MOAI22 U20003 ( .A1(n28918), .A2(n1819), .B1(ram[6841]), .B2(n1820), 
        .ZN(n11082) );
  MOAI22 U20004 ( .A1(n28683), .A2(n1819), .B1(ram[6842]), .B2(n1820), 
        .ZN(n11083) );
  MOAI22 U20005 ( .A1(n28448), .A2(n1819), .B1(ram[6843]), .B2(n1820), 
        .ZN(n11084) );
  MOAI22 U20006 ( .A1(n28213), .A2(n1819), .B1(ram[6844]), .B2(n1820), 
        .ZN(n11085) );
  MOAI22 U20007 ( .A1(n27978), .A2(n1819), .B1(ram[6845]), .B2(n1820), 
        .ZN(n11086) );
  MOAI22 U20008 ( .A1(n27743), .A2(n1819), .B1(ram[6846]), .B2(n1820), 
        .ZN(n11087) );
  MOAI22 U20009 ( .A1(n27508), .A2(n1819), .B1(ram[6847]), .B2(n1820), 
        .ZN(n11088) );
  MOAI22 U20010 ( .A1(n29153), .A2(n1821), .B1(ram[6848]), .B2(n1822), 
        .ZN(n11089) );
  MOAI22 U20011 ( .A1(n28918), .A2(n1821), .B1(ram[6849]), .B2(n1822), 
        .ZN(n11090) );
  MOAI22 U20012 ( .A1(n28683), .A2(n1821), .B1(ram[6850]), .B2(n1822), 
        .ZN(n11091) );
  MOAI22 U20013 ( .A1(n28448), .A2(n1821), .B1(ram[6851]), .B2(n1822), 
        .ZN(n11092) );
  MOAI22 U20014 ( .A1(n28213), .A2(n1821), .B1(ram[6852]), .B2(n1822), 
        .ZN(n11093) );
  MOAI22 U20015 ( .A1(n27978), .A2(n1821), .B1(ram[6853]), .B2(n1822), 
        .ZN(n11094) );
  MOAI22 U20016 ( .A1(n27743), .A2(n1821), .B1(ram[6854]), .B2(n1822), 
        .ZN(n11095) );
  MOAI22 U20017 ( .A1(n27508), .A2(n1821), .B1(ram[6855]), .B2(n1822), 
        .ZN(n11096) );
  MOAI22 U20018 ( .A1(n29153), .A2(n1823), .B1(ram[6856]), .B2(n1824), 
        .ZN(n11097) );
  MOAI22 U20019 ( .A1(n28918), .A2(n1823), .B1(ram[6857]), .B2(n1824), 
        .ZN(n11098) );
  MOAI22 U20020 ( .A1(n28683), .A2(n1823), .B1(ram[6858]), .B2(n1824), 
        .ZN(n11099) );
  MOAI22 U20021 ( .A1(n28448), .A2(n1823), .B1(ram[6859]), .B2(n1824), 
        .ZN(n11100) );
  MOAI22 U20022 ( .A1(n28213), .A2(n1823), .B1(ram[6860]), .B2(n1824), 
        .ZN(n11101) );
  MOAI22 U20023 ( .A1(n27978), .A2(n1823), .B1(ram[6861]), .B2(n1824), 
        .ZN(n11102) );
  MOAI22 U20024 ( .A1(n27743), .A2(n1823), .B1(ram[6862]), .B2(n1824), 
        .ZN(n11103) );
  MOAI22 U20025 ( .A1(n27508), .A2(n1823), .B1(ram[6863]), .B2(n1824), 
        .ZN(n11104) );
  MOAI22 U20026 ( .A1(n29154), .A2(n1825), .B1(ram[6864]), .B2(n1826), 
        .ZN(n11105) );
  MOAI22 U20027 ( .A1(n28919), .A2(n1825), .B1(ram[6865]), .B2(n1826), 
        .ZN(n11106) );
  MOAI22 U20028 ( .A1(n28684), .A2(n1825), .B1(ram[6866]), .B2(n1826), 
        .ZN(n11107) );
  MOAI22 U20029 ( .A1(n28449), .A2(n1825), .B1(ram[6867]), .B2(n1826), 
        .ZN(n11108) );
  MOAI22 U20030 ( .A1(n28214), .A2(n1825), .B1(ram[6868]), .B2(n1826), 
        .ZN(n11109) );
  MOAI22 U20031 ( .A1(n27979), .A2(n1825), .B1(ram[6869]), .B2(n1826), 
        .ZN(n11110) );
  MOAI22 U20032 ( .A1(n27744), .A2(n1825), .B1(ram[6870]), .B2(n1826), 
        .ZN(n11111) );
  MOAI22 U20033 ( .A1(n27509), .A2(n1825), .B1(ram[6871]), .B2(n1826), 
        .ZN(n11112) );
  MOAI22 U20034 ( .A1(n29154), .A2(n1827), .B1(ram[6872]), .B2(n1828), 
        .ZN(n11113) );
  MOAI22 U20035 ( .A1(n28919), .A2(n1827), .B1(ram[6873]), .B2(n1828), 
        .ZN(n11114) );
  MOAI22 U20036 ( .A1(n28684), .A2(n1827), .B1(ram[6874]), .B2(n1828), 
        .ZN(n11115) );
  MOAI22 U20037 ( .A1(n28449), .A2(n1827), .B1(ram[6875]), .B2(n1828), 
        .ZN(n11116) );
  MOAI22 U20038 ( .A1(n28214), .A2(n1827), .B1(ram[6876]), .B2(n1828), 
        .ZN(n11117) );
  MOAI22 U20039 ( .A1(n27979), .A2(n1827), .B1(ram[6877]), .B2(n1828), 
        .ZN(n11118) );
  MOAI22 U20040 ( .A1(n27744), .A2(n1827), .B1(ram[6878]), .B2(n1828), 
        .ZN(n11119) );
  MOAI22 U20041 ( .A1(n27509), .A2(n1827), .B1(ram[6879]), .B2(n1828), 
        .ZN(n11120) );
  MOAI22 U20042 ( .A1(n29154), .A2(n1829), .B1(ram[6880]), .B2(n1830), 
        .ZN(n11121) );
  MOAI22 U20043 ( .A1(n28919), .A2(n1829), .B1(ram[6881]), .B2(n1830), 
        .ZN(n11122) );
  MOAI22 U20044 ( .A1(n28684), .A2(n1829), .B1(ram[6882]), .B2(n1830), 
        .ZN(n11123) );
  MOAI22 U20045 ( .A1(n28449), .A2(n1829), .B1(ram[6883]), .B2(n1830), 
        .ZN(n11124) );
  MOAI22 U20046 ( .A1(n28214), .A2(n1829), .B1(ram[6884]), .B2(n1830), 
        .ZN(n11125) );
  MOAI22 U20047 ( .A1(n27979), .A2(n1829), .B1(ram[6885]), .B2(n1830), 
        .ZN(n11126) );
  MOAI22 U20048 ( .A1(n27744), .A2(n1829), .B1(ram[6886]), .B2(n1830), 
        .ZN(n11127) );
  MOAI22 U20049 ( .A1(n27509), .A2(n1829), .B1(ram[6887]), .B2(n1830), 
        .ZN(n11128) );
  MOAI22 U20050 ( .A1(n29154), .A2(n1831), .B1(ram[6888]), .B2(n1832), 
        .ZN(n11129) );
  MOAI22 U20051 ( .A1(n28919), .A2(n1831), .B1(ram[6889]), .B2(n1832), 
        .ZN(n11130) );
  MOAI22 U20052 ( .A1(n28684), .A2(n1831), .B1(ram[6890]), .B2(n1832), 
        .ZN(n11131) );
  MOAI22 U20053 ( .A1(n28449), .A2(n1831), .B1(ram[6891]), .B2(n1832), 
        .ZN(n11132) );
  MOAI22 U20054 ( .A1(n28214), .A2(n1831), .B1(ram[6892]), .B2(n1832), 
        .ZN(n11133) );
  MOAI22 U20055 ( .A1(n27979), .A2(n1831), .B1(ram[6893]), .B2(n1832), 
        .ZN(n11134) );
  MOAI22 U20056 ( .A1(n27744), .A2(n1831), .B1(ram[6894]), .B2(n1832), 
        .ZN(n11135) );
  MOAI22 U20057 ( .A1(n27509), .A2(n1831), .B1(ram[6895]), .B2(n1832), 
        .ZN(n11136) );
  MOAI22 U20058 ( .A1(n29154), .A2(n1833), .B1(ram[6896]), .B2(n1834), 
        .ZN(n11137) );
  MOAI22 U20059 ( .A1(n28919), .A2(n1833), .B1(ram[6897]), .B2(n1834), 
        .ZN(n11138) );
  MOAI22 U20060 ( .A1(n28684), .A2(n1833), .B1(ram[6898]), .B2(n1834), 
        .ZN(n11139) );
  MOAI22 U20061 ( .A1(n28449), .A2(n1833), .B1(ram[6899]), .B2(n1834), 
        .ZN(n11140) );
  MOAI22 U20062 ( .A1(n28214), .A2(n1833), .B1(ram[6900]), .B2(n1834), 
        .ZN(n11141) );
  MOAI22 U20063 ( .A1(n27979), .A2(n1833), .B1(ram[6901]), .B2(n1834), 
        .ZN(n11142) );
  MOAI22 U20064 ( .A1(n27744), .A2(n1833), .B1(ram[6902]), .B2(n1834), 
        .ZN(n11143) );
  MOAI22 U20065 ( .A1(n27509), .A2(n1833), .B1(ram[6903]), .B2(n1834), 
        .ZN(n11144) );
  MOAI22 U20066 ( .A1(n29154), .A2(n1835), .B1(ram[6904]), .B2(n1836), 
        .ZN(n11145) );
  MOAI22 U20067 ( .A1(n28919), .A2(n1835), .B1(ram[6905]), .B2(n1836), 
        .ZN(n11146) );
  MOAI22 U20068 ( .A1(n28684), .A2(n1835), .B1(ram[6906]), .B2(n1836), 
        .ZN(n11147) );
  MOAI22 U20069 ( .A1(n28449), .A2(n1835), .B1(ram[6907]), .B2(n1836), 
        .ZN(n11148) );
  MOAI22 U20070 ( .A1(n28214), .A2(n1835), .B1(ram[6908]), .B2(n1836), 
        .ZN(n11149) );
  MOAI22 U20071 ( .A1(n27979), .A2(n1835), .B1(ram[6909]), .B2(n1836), 
        .ZN(n11150) );
  MOAI22 U20072 ( .A1(n27744), .A2(n1835), .B1(ram[6910]), .B2(n1836), 
        .ZN(n11151) );
  MOAI22 U20073 ( .A1(n27509), .A2(n1835), .B1(ram[6911]), .B2(n1836), 
        .ZN(n11152) );
  MOAI22 U20074 ( .A1(n29154), .A2(n1837), .B1(ram[6912]), .B2(n1838), 
        .ZN(n11153) );
  MOAI22 U20075 ( .A1(n28919), .A2(n1837), .B1(ram[6913]), .B2(n1838), 
        .ZN(n11154) );
  MOAI22 U20076 ( .A1(n28684), .A2(n1837), .B1(ram[6914]), .B2(n1838), 
        .ZN(n11155) );
  MOAI22 U20077 ( .A1(n28449), .A2(n1837), .B1(ram[6915]), .B2(n1838), 
        .ZN(n11156) );
  MOAI22 U20078 ( .A1(n28214), .A2(n1837), .B1(ram[6916]), .B2(n1838), 
        .ZN(n11157) );
  MOAI22 U20079 ( .A1(n27979), .A2(n1837), .B1(ram[6917]), .B2(n1838), 
        .ZN(n11158) );
  MOAI22 U20080 ( .A1(n27744), .A2(n1837), .B1(ram[6918]), .B2(n1838), 
        .ZN(n11159) );
  MOAI22 U20081 ( .A1(n27509), .A2(n1837), .B1(ram[6919]), .B2(n1838), 
        .ZN(n11160) );
  MOAI22 U20082 ( .A1(n29154), .A2(n1839), .B1(ram[6920]), .B2(n1840), 
        .ZN(n11161) );
  MOAI22 U20083 ( .A1(n28919), .A2(n1839), .B1(ram[6921]), .B2(n1840), 
        .ZN(n11162) );
  MOAI22 U20084 ( .A1(n28684), .A2(n1839), .B1(ram[6922]), .B2(n1840), 
        .ZN(n11163) );
  MOAI22 U20085 ( .A1(n28449), .A2(n1839), .B1(ram[6923]), .B2(n1840), 
        .ZN(n11164) );
  MOAI22 U20086 ( .A1(n28214), .A2(n1839), .B1(ram[6924]), .B2(n1840), 
        .ZN(n11165) );
  MOAI22 U20087 ( .A1(n27979), .A2(n1839), .B1(ram[6925]), .B2(n1840), 
        .ZN(n11166) );
  MOAI22 U20088 ( .A1(n27744), .A2(n1839), .B1(ram[6926]), .B2(n1840), 
        .ZN(n11167) );
  MOAI22 U20089 ( .A1(n27509), .A2(n1839), .B1(ram[6927]), .B2(n1840), 
        .ZN(n11168) );
  MOAI22 U20090 ( .A1(n29154), .A2(n1841), .B1(ram[6928]), .B2(n1842), 
        .ZN(n11169) );
  MOAI22 U20091 ( .A1(n28919), .A2(n1841), .B1(ram[6929]), .B2(n1842), 
        .ZN(n11170) );
  MOAI22 U20092 ( .A1(n28684), .A2(n1841), .B1(ram[6930]), .B2(n1842), 
        .ZN(n11171) );
  MOAI22 U20093 ( .A1(n28449), .A2(n1841), .B1(ram[6931]), .B2(n1842), 
        .ZN(n11172) );
  MOAI22 U20094 ( .A1(n28214), .A2(n1841), .B1(ram[6932]), .B2(n1842), 
        .ZN(n11173) );
  MOAI22 U20095 ( .A1(n27979), .A2(n1841), .B1(ram[6933]), .B2(n1842), 
        .ZN(n11174) );
  MOAI22 U20096 ( .A1(n27744), .A2(n1841), .B1(ram[6934]), .B2(n1842), 
        .ZN(n11175) );
  MOAI22 U20097 ( .A1(n27509), .A2(n1841), .B1(ram[6935]), .B2(n1842), 
        .ZN(n11176) );
  MOAI22 U20098 ( .A1(n29154), .A2(n1843), .B1(ram[6936]), .B2(n1844), 
        .ZN(n11177) );
  MOAI22 U20099 ( .A1(n28919), .A2(n1843), .B1(ram[6937]), .B2(n1844), 
        .ZN(n11178) );
  MOAI22 U20100 ( .A1(n28684), .A2(n1843), .B1(ram[6938]), .B2(n1844), 
        .ZN(n11179) );
  MOAI22 U20101 ( .A1(n28449), .A2(n1843), .B1(ram[6939]), .B2(n1844), 
        .ZN(n11180) );
  MOAI22 U20102 ( .A1(n28214), .A2(n1843), .B1(ram[6940]), .B2(n1844), 
        .ZN(n11181) );
  MOAI22 U20103 ( .A1(n27979), .A2(n1843), .B1(ram[6941]), .B2(n1844), 
        .ZN(n11182) );
  MOAI22 U20104 ( .A1(n27744), .A2(n1843), .B1(ram[6942]), .B2(n1844), 
        .ZN(n11183) );
  MOAI22 U20105 ( .A1(n27509), .A2(n1843), .B1(ram[6943]), .B2(n1844), 
        .ZN(n11184) );
  MOAI22 U20106 ( .A1(n29154), .A2(n1845), .B1(ram[6944]), .B2(n1846), 
        .ZN(n11185) );
  MOAI22 U20107 ( .A1(n28919), .A2(n1845), .B1(ram[6945]), .B2(n1846), 
        .ZN(n11186) );
  MOAI22 U20108 ( .A1(n28684), .A2(n1845), .B1(ram[6946]), .B2(n1846), 
        .ZN(n11187) );
  MOAI22 U20109 ( .A1(n28449), .A2(n1845), .B1(ram[6947]), .B2(n1846), 
        .ZN(n11188) );
  MOAI22 U20110 ( .A1(n28214), .A2(n1845), .B1(ram[6948]), .B2(n1846), 
        .ZN(n11189) );
  MOAI22 U20111 ( .A1(n27979), .A2(n1845), .B1(ram[6949]), .B2(n1846), 
        .ZN(n11190) );
  MOAI22 U20112 ( .A1(n27744), .A2(n1845), .B1(ram[6950]), .B2(n1846), 
        .ZN(n11191) );
  MOAI22 U20113 ( .A1(n27509), .A2(n1845), .B1(ram[6951]), .B2(n1846), 
        .ZN(n11192) );
  MOAI22 U20114 ( .A1(n29154), .A2(n1847), .B1(ram[6952]), .B2(n1848), 
        .ZN(n11193) );
  MOAI22 U20115 ( .A1(n28919), .A2(n1847), .B1(ram[6953]), .B2(n1848), 
        .ZN(n11194) );
  MOAI22 U20116 ( .A1(n28684), .A2(n1847), .B1(ram[6954]), .B2(n1848), 
        .ZN(n11195) );
  MOAI22 U20117 ( .A1(n28449), .A2(n1847), .B1(ram[6955]), .B2(n1848), 
        .ZN(n11196) );
  MOAI22 U20118 ( .A1(n28214), .A2(n1847), .B1(ram[6956]), .B2(n1848), 
        .ZN(n11197) );
  MOAI22 U20119 ( .A1(n27979), .A2(n1847), .B1(ram[6957]), .B2(n1848), 
        .ZN(n11198) );
  MOAI22 U20120 ( .A1(n27744), .A2(n1847), .B1(ram[6958]), .B2(n1848), 
        .ZN(n11199) );
  MOAI22 U20121 ( .A1(n27509), .A2(n1847), .B1(ram[6959]), .B2(n1848), 
        .ZN(n11200) );
  MOAI22 U20122 ( .A1(n29154), .A2(n1849), .B1(ram[6960]), .B2(n1850), 
        .ZN(n11201) );
  MOAI22 U20123 ( .A1(n28919), .A2(n1849), .B1(ram[6961]), .B2(n1850), 
        .ZN(n11202) );
  MOAI22 U20124 ( .A1(n28684), .A2(n1849), .B1(ram[6962]), .B2(n1850), 
        .ZN(n11203) );
  MOAI22 U20125 ( .A1(n28449), .A2(n1849), .B1(ram[6963]), .B2(n1850), 
        .ZN(n11204) );
  MOAI22 U20126 ( .A1(n28214), .A2(n1849), .B1(ram[6964]), .B2(n1850), 
        .ZN(n11205) );
  MOAI22 U20127 ( .A1(n27979), .A2(n1849), .B1(ram[6965]), .B2(n1850), 
        .ZN(n11206) );
  MOAI22 U20128 ( .A1(n27744), .A2(n1849), .B1(ram[6966]), .B2(n1850), 
        .ZN(n11207) );
  MOAI22 U20129 ( .A1(n27509), .A2(n1849), .B1(ram[6967]), .B2(n1850), 
        .ZN(n11208) );
  MOAI22 U20130 ( .A1(n29155), .A2(n1851), .B1(ram[6968]), .B2(n1852), 
        .ZN(n11209) );
  MOAI22 U20131 ( .A1(n28920), .A2(n1851), .B1(ram[6969]), .B2(n1852), 
        .ZN(n11210) );
  MOAI22 U20132 ( .A1(n28685), .A2(n1851), .B1(ram[6970]), .B2(n1852), 
        .ZN(n11211) );
  MOAI22 U20133 ( .A1(n28450), .A2(n1851), .B1(ram[6971]), .B2(n1852), 
        .ZN(n11212) );
  MOAI22 U20134 ( .A1(n28215), .A2(n1851), .B1(ram[6972]), .B2(n1852), 
        .ZN(n11213) );
  MOAI22 U20135 ( .A1(n27980), .A2(n1851), .B1(ram[6973]), .B2(n1852), 
        .ZN(n11214) );
  MOAI22 U20136 ( .A1(n27745), .A2(n1851), .B1(ram[6974]), .B2(n1852), 
        .ZN(n11215) );
  MOAI22 U20137 ( .A1(n27510), .A2(n1851), .B1(ram[6975]), .B2(n1852), 
        .ZN(n11216) );
  MOAI22 U20138 ( .A1(n29155), .A2(n1853), .B1(ram[6976]), .B2(n1854), 
        .ZN(n11217) );
  MOAI22 U20139 ( .A1(n28920), .A2(n1853), .B1(ram[6977]), .B2(n1854), 
        .ZN(n11218) );
  MOAI22 U20140 ( .A1(n28685), .A2(n1853), .B1(ram[6978]), .B2(n1854), 
        .ZN(n11219) );
  MOAI22 U20141 ( .A1(n28450), .A2(n1853), .B1(ram[6979]), .B2(n1854), 
        .ZN(n11220) );
  MOAI22 U20142 ( .A1(n28215), .A2(n1853), .B1(ram[6980]), .B2(n1854), 
        .ZN(n11221) );
  MOAI22 U20143 ( .A1(n27980), .A2(n1853), .B1(ram[6981]), .B2(n1854), 
        .ZN(n11222) );
  MOAI22 U20144 ( .A1(n27745), .A2(n1853), .B1(ram[6982]), .B2(n1854), 
        .ZN(n11223) );
  MOAI22 U20145 ( .A1(n27510), .A2(n1853), .B1(ram[6983]), .B2(n1854), 
        .ZN(n11224) );
  MOAI22 U20146 ( .A1(n29155), .A2(n1855), .B1(ram[6984]), .B2(n1856), 
        .ZN(n11225) );
  MOAI22 U20147 ( .A1(n28920), .A2(n1855), .B1(ram[6985]), .B2(n1856), 
        .ZN(n11226) );
  MOAI22 U20148 ( .A1(n28685), .A2(n1855), .B1(ram[6986]), .B2(n1856), 
        .ZN(n11227) );
  MOAI22 U20149 ( .A1(n28450), .A2(n1855), .B1(ram[6987]), .B2(n1856), 
        .ZN(n11228) );
  MOAI22 U20150 ( .A1(n28215), .A2(n1855), .B1(ram[6988]), .B2(n1856), 
        .ZN(n11229) );
  MOAI22 U20151 ( .A1(n27980), .A2(n1855), .B1(ram[6989]), .B2(n1856), 
        .ZN(n11230) );
  MOAI22 U20152 ( .A1(n27745), .A2(n1855), .B1(ram[6990]), .B2(n1856), 
        .ZN(n11231) );
  MOAI22 U20153 ( .A1(n27510), .A2(n1855), .B1(ram[6991]), .B2(n1856), 
        .ZN(n11232) );
  MOAI22 U20154 ( .A1(n29155), .A2(n1857), .B1(ram[6992]), .B2(n1858), 
        .ZN(n11233) );
  MOAI22 U20155 ( .A1(n28920), .A2(n1857), .B1(ram[6993]), .B2(n1858), 
        .ZN(n11234) );
  MOAI22 U20156 ( .A1(n28685), .A2(n1857), .B1(ram[6994]), .B2(n1858), 
        .ZN(n11235) );
  MOAI22 U20157 ( .A1(n28450), .A2(n1857), .B1(ram[6995]), .B2(n1858), 
        .ZN(n11236) );
  MOAI22 U20158 ( .A1(n28215), .A2(n1857), .B1(ram[6996]), .B2(n1858), 
        .ZN(n11237) );
  MOAI22 U20159 ( .A1(n27980), .A2(n1857), .B1(ram[6997]), .B2(n1858), 
        .ZN(n11238) );
  MOAI22 U20160 ( .A1(n27745), .A2(n1857), .B1(ram[6998]), .B2(n1858), 
        .ZN(n11239) );
  MOAI22 U20161 ( .A1(n27510), .A2(n1857), .B1(ram[6999]), .B2(n1858), 
        .ZN(n11240) );
  MOAI22 U20162 ( .A1(n29155), .A2(n1859), .B1(ram[7000]), .B2(n1860), 
        .ZN(n11241) );
  MOAI22 U20163 ( .A1(n28920), .A2(n1859), .B1(ram[7001]), .B2(n1860), 
        .ZN(n11242) );
  MOAI22 U20164 ( .A1(n28685), .A2(n1859), .B1(ram[7002]), .B2(n1860), 
        .ZN(n11243) );
  MOAI22 U20165 ( .A1(n28450), .A2(n1859), .B1(ram[7003]), .B2(n1860), 
        .ZN(n11244) );
  MOAI22 U20166 ( .A1(n28215), .A2(n1859), .B1(ram[7004]), .B2(n1860), 
        .ZN(n11245) );
  MOAI22 U20167 ( .A1(n27980), .A2(n1859), .B1(ram[7005]), .B2(n1860), 
        .ZN(n11246) );
  MOAI22 U20168 ( .A1(n27745), .A2(n1859), .B1(ram[7006]), .B2(n1860), 
        .ZN(n11247) );
  MOAI22 U20169 ( .A1(n27510), .A2(n1859), .B1(ram[7007]), .B2(n1860), 
        .ZN(n11248) );
  MOAI22 U20170 ( .A1(n29155), .A2(n1861), .B1(ram[7008]), .B2(n1862), 
        .ZN(n11249) );
  MOAI22 U20171 ( .A1(n28920), .A2(n1861), .B1(ram[7009]), .B2(n1862), 
        .ZN(n11250) );
  MOAI22 U20172 ( .A1(n28685), .A2(n1861), .B1(ram[7010]), .B2(n1862), 
        .ZN(n11251) );
  MOAI22 U20173 ( .A1(n28450), .A2(n1861), .B1(ram[7011]), .B2(n1862), 
        .ZN(n11252) );
  MOAI22 U20174 ( .A1(n28215), .A2(n1861), .B1(ram[7012]), .B2(n1862), 
        .ZN(n11253) );
  MOAI22 U20175 ( .A1(n27980), .A2(n1861), .B1(ram[7013]), .B2(n1862), 
        .ZN(n11254) );
  MOAI22 U20176 ( .A1(n27745), .A2(n1861), .B1(ram[7014]), .B2(n1862), 
        .ZN(n11255) );
  MOAI22 U20177 ( .A1(n27510), .A2(n1861), .B1(ram[7015]), .B2(n1862), 
        .ZN(n11256) );
  MOAI22 U20178 ( .A1(n29155), .A2(n1863), .B1(ram[7016]), .B2(n1864), 
        .ZN(n11257) );
  MOAI22 U20179 ( .A1(n28920), .A2(n1863), .B1(ram[7017]), .B2(n1864), 
        .ZN(n11258) );
  MOAI22 U20180 ( .A1(n28685), .A2(n1863), .B1(ram[7018]), .B2(n1864), 
        .ZN(n11259) );
  MOAI22 U20181 ( .A1(n28450), .A2(n1863), .B1(ram[7019]), .B2(n1864), 
        .ZN(n11260) );
  MOAI22 U20182 ( .A1(n28215), .A2(n1863), .B1(ram[7020]), .B2(n1864), 
        .ZN(n11261) );
  MOAI22 U20183 ( .A1(n27980), .A2(n1863), .B1(ram[7021]), .B2(n1864), 
        .ZN(n11262) );
  MOAI22 U20184 ( .A1(n27745), .A2(n1863), .B1(ram[7022]), .B2(n1864), 
        .ZN(n11263) );
  MOAI22 U20185 ( .A1(n27510), .A2(n1863), .B1(ram[7023]), .B2(n1864), 
        .ZN(n11264) );
  MOAI22 U20186 ( .A1(n29155), .A2(n1865), .B1(ram[7024]), .B2(n1866), 
        .ZN(n11265) );
  MOAI22 U20187 ( .A1(n28920), .A2(n1865), .B1(ram[7025]), .B2(n1866), 
        .ZN(n11266) );
  MOAI22 U20188 ( .A1(n28685), .A2(n1865), .B1(ram[7026]), .B2(n1866), 
        .ZN(n11267) );
  MOAI22 U20189 ( .A1(n28450), .A2(n1865), .B1(ram[7027]), .B2(n1866), 
        .ZN(n11268) );
  MOAI22 U20190 ( .A1(n28215), .A2(n1865), .B1(ram[7028]), .B2(n1866), 
        .ZN(n11269) );
  MOAI22 U20191 ( .A1(n27980), .A2(n1865), .B1(ram[7029]), .B2(n1866), 
        .ZN(n11270) );
  MOAI22 U20192 ( .A1(n27745), .A2(n1865), .B1(ram[7030]), .B2(n1866), 
        .ZN(n11271) );
  MOAI22 U20193 ( .A1(n27510), .A2(n1865), .B1(ram[7031]), .B2(n1866), 
        .ZN(n11272) );
  MOAI22 U20194 ( .A1(n29155), .A2(n1867), .B1(ram[7032]), .B2(n1868), 
        .ZN(n11273) );
  MOAI22 U20195 ( .A1(n28920), .A2(n1867), .B1(ram[7033]), .B2(n1868), 
        .ZN(n11274) );
  MOAI22 U20196 ( .A1(n28685), .A2(n1867), .B1(ram[7034]), .B2(n1868), 
        .ZN(n11275) );
  MOAI22 U20197 ( .A1(n28450), .A2(n1867), .B1(ram[7035]), .B2(n1868), 
        .ZN(n11276) );
  MOAI22 U20198 ( .A1(n28215), .A2(n1867), .B1(ram[7036]), .B2(n1868), 
        .ZN(n11277) );
  MOAI22 U20199 ( .A1(n27980), .A2(n1867), .B1(ram[7037]), .B2(n1868), 
        .ZN(n11278) );
  MOAI22 U20200 ( .A1(n27745), .A2(n1867), .B1(ram[7038]), .B2(n1868), 
        .ZN(n11279) );
  MOAI22 U20201 ( .A1(n27510), .A2(n1867), .B1(ram[7039]), .B2(n1868), 
        .ZN(n11280) );
  MOAI22 U20202 ( .A1(n29155), .A2(n1869), .B1(ram[7040]), .B2(n1870), 
        .ZN(n11281) );
  MOAI22 U20203 ( .A1(n28920), .A2(n1869), .B1(ram[7041]), .B2(n1870), 
        .ZN(n11282) );
  MOAI22 U20204 ( .A1(n28685), .A2(n1869), .B1(ram[7042]), .B2(n1870), 
        .ZN(n11283) );
  MOAI22 U20205 ( .A1(n28450), .A2(n1869), .B1(ram[7043]), .B2(n1870), 
        .ZN(n11284) );
  MOAI22 U20206 ( .A1(n28215), .A2(n1869), .B1(ram[7044]), .B2(n1870), 
        .ZN(n11285) );
  MOAI22 U20207 ( .A1(n27980), .A2(n1869), .B1(ram[7045]), .B2(n1870), 
        .ZN(n11286) );
  MOAI22 U20208 ( .A1(n27745), .A2(n1869), .B1(ram[7046]), .B2(n1870), 
        .ZN(n11287) );
  MOAI22 U20209 ( .A1(n27510), .A2(n1869), .B1(ram[7047]), .B2(n1870), 
        .ZN(n11288) );
  MOAI22 U20210 ( .A1(n29155), .A2(n1871), .B1(ram[7048]), .B2(n1872), 
        .ZN(n11289) );
  MOAI22 U20211 ( .A1(n28920), .A2(n1871), .B1(ram[7049]), .B2(n1872), 
        .ZN(n11290) );
  MOAI22 U20212 ( .A1(n28685), .A2(n1871), .B1(ram[7050]), .B2(n1872), 
        .ZN(n11291) );
  MOAI22 U20213 ( .A1(n28450), .A2(n1871), .B1(ram[7051]), .B2(n1872), 
        .ZN(n11292) );
  MOAI22 U20214 ( .A1(n28215), .A2(n1871), .B1(ram[7052]), .B2(n1872), 
        .ZN(n11293) );
  MOAI22 U20215 ( .A1(n27980), .A2(n1871), .B1(ram[7053]), .B2(n1872), 
        .ZN(n11294) );
  MOAI22 U20216 ( .A1(n27745), .A2(n1871), .B1(ram[7054]), .B2(n1872), 
        .ZN(n11295) );
  MOAI22 U20217 ( .A1(n27510), .A2(n1871), .B1(ram[7055]), .B2(n1872), 
        .ZN(n11296) );
  MOAI22 U20218 ( .A1(n29155), .A2(n1873), .B1(ram[7056]), .B2(n1874), 
        .ZN(n11297) );
  MOAI22 U20219 ( .A1(n28920), .A2(n1873), .B1(ram[7057]), .B2(n1874), 
        .ZN(n11298) );
  MOAI22 U20220 ( .A1(n28685), .A2(n1873), .B1(ram[7058]), .B2(n1874), 
        .ZN(n11299) );
  MOAI22 U20221 ( .A1(n28450), .A2(n1873), .B1(ram[7059]), .B2(n1874), 
        .ZN(n11300) );
  MOAI22 U20222 ( .A1(n28215), .A2(n1873), .B1(ram[7060]), .B2(n1874), 
        .ZN(n11301) );
  MOAI22 U20223 ( .A1(n27980), .A2(n1873), .B1(ram[7061]), .B2(n1874), 
        .ZN(n11302) );
  MOAI22 U20224 ( .A1(n27745), .A2(n1873), .B1(ram[7062]), .B2(n1874), 
        .ZN(n11303) );
  MOAI22 U20225 ( .A1(n27510), .A2(n1873), .B1(ram[7063]), .B2(n1874), 
        .ZN(n11304) );
  MOAI22 U20226 ( .A1(n29155), .A2(n1875), .B1(ram[7064]), .B2(n1876), 
        .ZN(n11305) );
  MOAI22 U20227 ( .A1(n28920), .A2(n1875), .B1(ram[7065]), .B2(n1876), 
        .ZN(n11306) );
  MOAI22 U20228 ( .A1(n28685), .A2(n1875), .B1(ram[7066]), .B2(n1876), 
        .ZN(n11307) );
  MOAI22 U20229 ( .A1(n28450), .A2(n1875), .B1(ram[7067]), .B2(n1876), 
        .ZN(n11308) );
  MOAI22 U20230 ( .A1(n28215), .A2(n1875), .B1(ram[7068]), .B2(n1876), 
        .ZN(n11309) );
  MOAI22 U20231 ( .A1(n27980), .A2(n1875), .B1(ram[7069]), .B2(n1876), 
        .ZN(n11310) );
  MOAI22 U20232 ( .A1(n27745), .A2(n1875), .B1(ram[7070]), .B2(n1876), 
        .ZN(n11311) );
  MOAI22 U20233 ( .A1(n27510), .A2(n1875), .B1(ram[7071]), .B2(n1876), 
        .ZN(n11312) );
  MOAI22 U20234 ( .A1(n29156), .A2(n1877), .B1(ram[7072]), .B2(n1878), 
        .ZN(n11313) );
  MOAI22 U20235 ( .A1(n28921), .A2(n1877), .B1(ram[7073]), .B2(n1878), 
        .ZN(n11314) );
  MOAI22 U20236 ( .A1(n28686), .A2(n1877), .B1(ram[7074]), .B2(n1878), 
        .ZN(n11315) );
  MOAI22 U20237 ( .A1(n28451), .A2(n1877), .B1(ram[7075]), .B2(n1878), 
        .ZN(n11316) );
  MOAI22 U20238 ( .A1(n28216), .A2(n1877), .B1(ram[7076]), .B2(n1878), 
        .ZN(n11317) );
  MOAI22 U20239 ( .A1(n27981), .A2(n1877), .B1(ram[7077]), .B2(n1878), 
        .ZN(n11318) );
  MOAI22 U20240 ( .A1(n27746), .A2(n1877), .B1(ram[7078]), .B2(n1878), 
        .ZN(n11319) );
  MOAI22 U20241 ( .A1(n27511), .A2(n1877), .B1(ram[7079]), .B2(n1878), 
        .ZN(n11320) );
  MOAI22 U20242 ( .A1(n29156), .A2(n1879), .B1(ram[7080]), .B2(n1880), 
        .ZN(n11321) );
  MOAI22 U20243 ( .A1(n28921), .A2(n1879), .B1(ram[7081]), .B2(n1880), 
        .ZN(n11322) );
  MOAI22 U20244 ( .A1(n28686), .A2(n1879), .B1(ram[7082]), .B2(n1880), 
        .ZN(n11323) );
  MOAI22 U20245 ( .A1(n28451), .A2(n1879), .B1(ram[7083]), .B2(n1880), 
        .ZN(n11324) );
  MOAI22 U20246 ( .A1(n28216), .A2(n1879), .B1(ram[7084]), .B2(n1880), 
        .ZN(n11325) );
  MOAI22 U20247 ( .A1(n27981), .A2(n1879), .B1(ram[7085]), .B2(n1880), 
        .ZN(n11326) );
  MOAI22 U20248 ( .A1(n27746), .A2(n1879), .B1(ram[7086]), .B2(n1880), 
        .ZN(n11327) );
  MOAI22 U20249 ( .A1(n27511), .A2(n1879), .B1(ram[7087]), .B2(n1880), 
        .ZN(n11328) );
  MOAI22 U20250 ( .A1(n29156), .A2(n1881), .B1(ram[7088]), .B2(n1882), 
        .ZN(n11329) );
  MOAI22 U20251 ( .A1(n28921), .A2(n1881), .B1(ram[7089]), .B2(n1882), 
        .ZN(n11330) );
  MOAI22 U20252 ( .A1(n28686), .A2(n1881), .B1(ram[7090]), .B2(n1882), 
        .ZN(n11331) );
  MOAI22 U20253 ( .A1(n28451), .A2(n1881), .B1(ram[7091]), .B2(n1882), 
        .ZN(n11332) );
  MOAI22 U20254 ( .A1(n28216), .A2(n1881), .B1(ram[7092]), .B2(n1882), 
        .ZN(n11333) );
  MOAI22 U20255 ( .A1(n27981), .A2(n1881), .B1(ram[7093]), .B2(n1882), 
        .ZN(n11334) );
  MOAI22 U20256 ( .A1(n27746), .A2(n1881), .B1(ram[7094]), .B2(n1882), 
        .ZN(n11335) );
  MOAI22 U20257 ( .A1(n27511), .A2(n1881), .B1(ram[7095]), .B2(n1882), 
        .ZN(n11336) );
  MOAI22 U20258 ( .A1(n29156), .A2(n1883), .B1(ram[7096]), .B2(n1884), 
        .ZN(n11337) );
  MOAI22 U20259 ( .A1(n28921), .A2(n1883), .B1(ram[7097]), .B2(n1884), 
        .ZN(n11338) );
  MOAI22 U20260 ( .A1(n28686), .A2(n1883), .B1(ram[7098]), .B2(n1884), 
        .ZN(n11339) );
  MOAI22 U20261 ( .A1(n28451), .A2(n1883), .B1(ram[7099]), .B2(n1884), 
        .ZN(n11340) );
  MOAI22 U20262 ( .A1(n28216), .A2(n1883), .B1(ram[7100]), .B2(n1884), 
        .ZN(n11341) );
  MOAI22 U20263 ( .A1(n27981), .A2(n1883), .B1(ram[7101]), .B2(n1884), 
        .ZN(n11342) );
  MOAI22 U20264 ( .A1(n27746), .A2(n1883), .B1(ram[7102]), .B2(n1884), 
        .ZN(n11343) );
  MOAI22 U20265 ( .A1(n27511), .A2(n1883), .B1(ram[7103]), .B2(n1884), 
        .ZN(n11344) );
  MOAI22 U20266 ( .A1(n29156), .A2(n1885), .B1(ram[7104]), .B2(n1886), 
        .ZN(n11345) );
  MOAI22 U20267 ( .A1(n28921), .A2(n1885), .B1(ram[7105]), .B2(n1886), 
        .ZN(n11346) );
  MOAI22 U20268 ( .A1(n28686), .A2(n1885), .B1(ram[7106]), .B2(n1886), 
        .ZN(n11347) );
  MOAI22 U20269 ( .A1(n28451), .A2(n1885), .B1(ram[7107]), .B2(n1886), 
        .ZN(n11348) );
  MOAI22 U20270 ( .A1(n28216), .A2(n1885), .B1(ram[7108]), .B2(n1886), 
        .ZN(n11349) );
  MOAI22 U20271 ( .A1(n27981), .A2(n1885), .B1(ram[7109]), .B2(n1886), 
        .ZN(n11350) );
  MOAI22 U20272 ( .A1(n27746), .A2(n1885), .B1(ram[7110]), .B2(n1886), 
        .ZN(n11351) );
  MOAI22 U20273 ( .A1(n27511), .A2(n1885), .B1(ram[7111]), .B2(n1886), 
        .ZN(n11352) );
  MOAI22 U20274 ( .A1(n29156), .A2(n1887), .B1(ram[7112]), .B2(n1888), 
        .ZN(n11353) );
  MOAI22 U20275 ( .A1(n28921), .A2(n1887), .B1(ram[7113]), .B2(n1888), 
        .ZN(n11354) );
  MOAI22 U20276 ( .A1(n28686), .A2(n1887), .B1(ram[7114]), .B2(n1888), 
        .ZN(n11355) );
  MOAI22 U20277 ( .A1(n28451), .A2(n1887), .B1(ram[7115]), .B2(n1888), 
        .ZN(n11356) );
  MOAI22 U20278 ( .A1(n28216), .A2(n1887), .B1(ram[7116]), .B2(n1888), 
        .ZN(n11357) );
  MOAI22 U20279 ( .A1(n27981), .A2(n1887), .B1(ram[7117]), .B2(n1888), 
        .ZN(n11358) );
  MOAI22 U20280 ( .A1(n27746), .A2(n1887), .B1(ram[7118]), .B2(n1888), 
        .ZN(n11359) );
  MOAI22 U20281 ( .A1(n27511), .A2(n1887), .B1(ram[7119]), .B2(n1888), 
        .ZN(n11360) );
  MOAI22 U20282 ( .A1(n29156), .A2(n1889), .B1(ram[7120]), .B2(n1890), 
        .ZN(n11361) );
  MOAI22 U20283 ( .A1(n28921), .A2(n1889), .B1(ram[7121]), .B2(n1890), 
        .ZN(n11362) );
  MOAI22 U20284 ( .A1(n28686), .A2(n1889), .B1(ram[7122]), .B2(n1890), 
        .ZN(n11363) );
  MOAI22 U20285 ( .A1(n28451), .A2(n1889), .B1(ram[7123]), .B2(n1890), 
        .ZN(n11364) );
  MOAI22 U20286 ( .A1(n28216), .A2(n1889), .B1(ram[7124]), .B2(n1890), 
        .ZN(n11365) );
  MOAI22 U20287 ( .A1(n27981), .A2(n1889), .B1(ram[7125]), .B2(n1890), 
        .ZN(n11366) );
  MOAI22 U20288 ( .A1(n27746), .A2(n1889), .B1(ram[7126]), .B2(n1890), 
        .ZN(n11367) );
  MOAI22 U20289 ( .A1(n27511), .A2(n1889), .B1(ram[7127]), .B2(n1890), 
        .ZN(n11368) );
  MOAI22 U20290 ( .A1(n29156), .A2(n1891), .B1(ram[7128]), .B2(n1892), 
        .ZN(n11369) );
  MOAI22 U20291 ( .A1(n28921), .A2(n1891), .B1(ram[7129]), .B2(n1892), 
        .ZN(n11370) );
  MOAI22 U20292 ( .A1(n28686), .A2(n1891), .B1(ram[7130]), .B2(n1892), 
        .ZN(n11371) );
  MOAI22 U20293 ( .A1(n28451), .A2(n1891), .B1(ram[7131]), .B2(n1892), 
        .ZN(n11372) );
  MOAI22 U20294 ( .A1(n28216), .A2(n1891), .B1(ram[7132]), .B2(n1892), 
        .ZN(n11373) );
  MOAI22 U20295 ( .A1(n27981), .A2(n1891), .B1(ram[7133]), .B2(n1892), 
        .ZN(n11374) );
  MOAI22 U20296 ( .A1(n27746), .A2(n1891), .B1(ram[7134]), .B2(n1892), 
        .ZN(n11375) );
  MOAI22 U20297 ( .A1(n27511), .A2(n1891), .B1(ram[7135]), .B2(n1892), 
        .ZN(n11376) );
  MOAI22 U20298 ( .A1(n29156), .A2(n1893), .B1(ram[7136]), .B2(n1894), 
        .ZN(n11377) );
  MOAI22 U20299 ( .A1(n28921), .A2(n1893), .B1(ram[7137]), .B2(n1894), 
        .ZN(n11378) );
  MOAI22 U20300 ( .A1(n28686), .A2(n1893), .B1(ram[7138]), .B2(n1894), 
        .ZN(n11379) );
  MOAI22 U20301 ( .A1(n28451), .A2(n1893), .B1(ram[7139]), .B2(n1894), 
        .ZN(n11380) );
  MOAI22 U20302 ( .A1(n28216), .A2(n1893), .B1(ram[7140]), .B2(n1894), 
        .ZN(n11381) );
  MOAI22 U20303 ( .A1(n27981), .A2(n1893), .B1(ram[7141]), .B2(n1894), 
        .ZN(n11382) );
  MOAI22 U20304 ( .A1(n27746), .A2(n1893), .B1(ram[7142]), .B2(n1894), 
        .ZN(n11383) );
  MOAI22 U20305 ( .A1(n27511), .A2(n1893), .B1(ram[7143]), .B2(n1894), 
        .ZN(n11384) );
  MOAI22 U20306 ( .A1(n29156), .A2(n1895), .B1(ram[7144]), .B2(n1896), 
        .ZN(n11385) );
  MOAI22 U20307 ( .A1(n28921), .A2(n1895), .B1(ram[7145]), .B2(n1896), 
        .ZN(n11386) );
  MOAI22 U20308 ( .A1(n28686), .A2(n1895), .B1(ram[7146]), .B2(n1896), 
        .ZN(n11387) );
  MOAI22 U20309 ( .A1(n28451), .A2(n1895), .B1(ram[7147]), .B2(n1896), 
        .ZN(n11388) );
  MOAI22 U20310 ( .A1(n28216), .A2(n1895), .B1(ram[7148]), .B2(n1896), 
        .ZN(n11389) );
  MOAI22 U20311 ( .A1(n27981), .A2(n1895), .B1(ram[7149]), .B2(n1896), 
        .ZN(n11390) );
  MOAI22 U20312 ( .A1(n27746), .A2(n1895), .B1(ram[7150]), .B2(n1896), 
        .ZN(n11391) );
  MOAI22 U20313 ( .A1(n27511), .A2(n1895), .B1(ram[7151]), .B2(n1896), 
        .ZN(n11392) );
  MOAI22 U20314 ( .A1(n29156), .A2(n1897), .B1(ram[7152]), .B2(n1898), 
        .ZN(n11393) );
  MOAI22 U20315 ( .A1(n28921), .A2(n1897), .B1(ram[7153]), .B2(n1898), 
        .ZN(n11394) );
  MOAI22 U20316 ( .A1(n28686), .A2(n1897), .B1(ram[7154]), .B2(n1898), 
        .ZN(n11395) );
  MOAI22 U20317 ( .A1(n28451), .A2(n1897), .B1(ram[7155]), .B2(n1898), 
        .ZN(n11396) );
  MOAI22 U20318 ( .A1(n28216), .A2(n1897), .B1(ram[7156]), .B2(n1898), 
        .ZN(n11397) );
  MOAI22 U20319 ( .A1(n27981), .A2(n1897), .B1(ram[7157]), .B2(n1898), 
        .ZN(n11398) );
  MOAI22 U20320 ( .A1(n27746), .A2(n1897), .B1(ram[7158]), .B2(n1898), 
        .ZN(n11399) );
  MOAI22 U20321 ( .A1(n27511), .A2(n1897), .B1(ram[7159]), .B2(n1898), 
        .ZN(n11400) );
  MOAI22 U20322 ( .A1(n29156), .A2(n1899), .B1(ram[7160]), .B2(n1900), 
        .ZN(n11401) );
  MOAI22 U20323 ( .A1(n28921), .A2(n1899), .B1(ram[7161]), .B2(n1900), 
        .ZN(n11402) );
  MOAI22 U20324 ( .A1(n28686), .A2(n1899), .B1(ram[7162]), .B2(n1900), 
        .ZN(n11403) );
  MOAI22 U20325 ( .A1(n28451), .A2(n1899), .B1(ram[7163]), .B2(n1900), 
        .ZN(n11404) );
  MOAI22 U20326 ( .A1(n28216), .A2(n1899), .B1(ram[7164]), .B2(n1900), 
        .ZN(n11405) );
  MOAI22 U20327 ( .A1(n27981), .A2(n1899), .B1(ram[7165]), .B2(n1900), 
        .ZN(n11406) );
  MOAI22 U20328 ( .A1(n27746), .A2(n1899), .B1(ram[7166]), .B2(n1900), 
        .ZN(n11407) );
  MOAI22 U20329 ( .A1(n27511), .A2(n1899), .B1(ram[7167]), .B2(n1900), 
        .ZN(n11408) );
  MOAI22 U20330 ( .A1(n29156), .A2(n1901), .B1(ram[7168]), .B2(n1902), 
        .ZN(n11409) );
  MOAI22 U20331 ( .A1(n28921), .A2(n1901), .B1(ram[7169]), .B2(n1902), 
        .ZN(n11410) );
  MOAI22 U20332 ( .A1(n28686), .A2(n1901), .B1(ram[7170]), .B2(n1902), 
        .ZN(n11411) );
  MOAI22 U20333 ( .A1(n28451), .A2(n1901), .B1(ram[7171]), .B2(n1902), 
        .ZN(n11412) );
  MOAI22 U20334 ( .A1(n28216), .A2(n1901), .B1(ram[7172]), .B2(n1902), 
        .ZN(n11413) );
  MOAI22 U20335 ( .A1(n27981), .A2(n1901), .B1(ram[7173]), .B2(n1902), 
        .ZN(n11414) );
  MOAI22 U20336 ( .A1(n27746), .A2(n1901), .B1(ram[7174]), .B2(n1902), 
        .ZN(n11415) );
  MOAI22 U20337 ( .A1(n27511), .A2(n1901), .B1(ram[7175]), .B2(n1902), 
        .ZN(n11416) );
  MOAI22 U20338 ( .A1(n29157), .A2(n1904), .B1(ram[7176]), .B2(n1905), 
        .ZN(n11417) );
  MOAI22 U20339 ( .A1(n28922), .A2(n1904), .B1(ram[7177]), .B2(n1905), 
        .ZN(n11418) );
  MOAI22 U20340 ( .A1(n28687), .A2(n1904), .B1(ram[7178]), .B2(n1905), 
        .ZN(n11419) );
  MOAI22 U20341 ( .A1(n28452), .A2(n1904), .B1(ram[7179]), .B2(n1905), 
        .ZN(n11420) );
  MOAI22 U20342 ( .A1(n28217), .A2(n1904), .B1(ram[7180]), .B2(n1905), 
        .ZN(n11421) );
  MOAI22 U20343 ( .A1(n27982), .A2(n1904), .B1(ram[7181]), .B2(n1905), 
        .ZN(n11422) );
  MOAI22 U20344 ( .A1(n27747), .A2(n1904), .B1(ram[7182]), .B2(n1905), 
        .ZN(n11423) );
  MOAI22 U20345 ( .A1(n27512), .A2(n1904), .B1(ram[7183]), .B2(n1905), 
        .ZN(n11424) );
  MOAI22 U20346 ( .A1(n29157), .A2(n1906), .B1(ram[7184]), .B2(n1907), 
        .ZN(n11425) );
  MOAI22 U20347 ( .A1(n28922), .A2(n1906), .B1(ram[7185]), .B2(n1907), 
        .ZN(n11426) );
  MOAI22 U20348 ( .A1(n28687), .A2(n1906), .B1(ram[7186]), .B2(n1907), 
        .ZN(n11427) );
  MOAI22 U20349 ( .A1(n28452), .A2(n1906), .B1(ram[7187]), .B2(n1907), 
        .ZN(n11428) );
  MOAI22 U20350 ( .A1(n28217), .A2(n1906), .B1(ram[7188]), .B2(n1907), 
        .ZN(n11429) );
  MOAI22 U20351 ( .A1(n27982), .A2(n1906), .B1(ram[7189]), .B2(n1907), 
        .ZN(n11430) );
  MOAI22 U20352 ( .A1(n27747), .A2(n1906), .B1(ram[7190]), .B2(n1907), 
        .ZN(n11431) );
  MOAI22 U20353 ( .A1(n27512), .A2(n1906), .B1(ram[7191]), .B2(n1907), 
        .ZN(n11432) );
  MOAI22 U20354 ( .A1(n29157), .A2(n1908), .B1(ram[7192]), .B2(n1909), 
        .ZN(n11433) );
  MOAI22 U20355 ( .A1(n28922), .A2(n1908), .B1(ram[7193]), .B2(n1909), 
        .ZN(n11434) );
  MOAI22 U20356 ( .A1(n28687), .A2(n1908), .B1(ram[7194]), .B2(n1909), 
        .ZN(n11435) );
  MOAI22 U20357 ( .A1(n28452), .A2(n1908), .B1(ram[7195]), .B2(n1909), 
        .ZN(n11436) );
  MOAI22 U20358 ( .A1(n28217), .A2(n1908), .B1(ram[7196]), .B2(n1909), 
        .ZN(n11437) );
  MOAI22 U20359 ( .A1(n27982), .A2(n1908), .B1(ram[7197]), .B2(n1909), 
        .ZN(n11438) );
  MOAI22 U20360 ( .A1(n27747), .A2(n1908), .B1(ram[7198]), .B2(n1909), 
        .ZN(n11439) );
  MOAI22 U20361 ( .A1(n27512), .A2(n1908), .B1(ram[7199]), .B2(n1909), 
        .ZN(n11440) );
  MOAI22 U20362 ( .A1(n29157), .A2(n1910), .B1(ram[7200]), .B2(n1911), 
        .ZN(n11441) );
  MOAI22 U20363 ( .A1(n28922), .A2(n1910), .B1(ram[7201]), .B2(n1911), 
        .ZN(n11442) );
  MOAI22 U20364 ( .A1(n28687), .A2(n1910), .B1(ram[7202]), .B2(n1911), 
        .ZN(n11443) );
  MOAI22 U20365 ( .A1(n28452), .A2(n1910), .B1(ram[7203]), .B2(n1911), 
        .ZN(n11444) );
  MOAI22 U20366 ( .A1(n28217), .A2(n1910), .B1(ram[7204]), .B2(n1911), 
        .ZN(n11445) );
  MOAI22 U20367 ( .A1(n27982), .A2(n1910), .B1(ram[7205]), .B2(n1911), 
        .ZN(n11446) );
  MOAI22 U20368 ( .A1(n27747), .A2(n1910), .B1(ram[7206]), .B2(n1911), 
        .ZN(n11447) );
  MOAI22 U20369 ( .A1(n27512), .A2(n1910), .B1(ram[7207]), .B2(n1911), 
        .ZN(n11448) );
  MOAI22 U20370 ( .A1(n29157), .A2(n1912), .B1(ram[7208]), .B2(n1913), 
        .ZN(n11449) );
  MOAI22 U20371 ( .A1(n28922), .A2(n1912), .B1(ram[7209]), .B2(n1913), 
        .ZN(n11450) );
  MOAI22 U20372 ( .A1(n28687), .A2(n1912), .B1(ram[7210]), .B2(n1913), 
        .ZN(n11451) );
  MOAI22 U20373 ( .A1(n28452), .A2(n1912), .B1(ram[7211]), .B2(n1913), 
        .ZN(n11452) );
  MOAI22 U20374 ( .A1(n28217), .A2(n1912), .B1(ram[7212]), .B2(n1913), 
        .ZN(n11453) );
  MOAI22 U20375 ( .A1(n27982), .A2(n1912), .B1(ram[7213]), .B2(n1913), 
        .ZN(n11454) );
  MOAI22 U20376 ( .A1(n27747), .A2(n1912), .B1(ram[7214]), .B2(n1913), 
        .ZN(n11455) );
  MOAI22 U20377 ( .A1(n27512), .A2(n1912), .B1(ram[7215]), .B2(n1913), 
        .ZN(n11456) );
  MOAI22 U20378 ( .A1(n29157), .A2(n1914), .B1(ram[7216]), .B2(n1915), 
        .ZN(n11457) );
  MOAI22 U20379 ( .A1(n28922), .A2(n1914), .B1(ram[7217]), .B2(n1915), 
        .ZN(n11458) );
  MOAI22 U20380 ( .A1(n28687), .A2(n1914), .B1(ram[7218]), .B2(n1915), 
        .ZN(n11459) );
  MOAI22 U20381 ( .A1(n28452), .A2(n1914), .B1(ram[7219]), .B2(n1915), 
        .ZN(n11460) );
  MOAI22 U20382 ( .A1(n28217), .A2(n1914), .B1(ram[7220]), .B2(n1915), 
        .ZN(n11461) );
  MOAI22 U20383 ( .A1(n27982), .A2(n1914), .B1(ram[7221]), .B2(n1915), 
        .ZN(n11462) );
  MOAI22 U20384 ( .A1(n27747), .A2(n1914), .B1(ram[7222]), .B2(n1915), 
        .ZN(n11463) );
  MOAI22 U20385 ( .A1(n27512), .A2(n1914), .B1(ram[7223]), .B2(n1915), 
        .ZN(n11464) );
  MOAI22 U20386 ( .A1(n29157), .A2(n1916), .B1(ram[7224]), .B2(n1917), 
        .ZN(n11465) );
  MOAI22 U20387 ( .A1(n28922), .A2(n1916), .B1(ram[7225]), .B2(n1917), 
        .ZN(n11466) );
  MOAI22 U20388 ( .A1(n28687), .A2(n1916), .B1(ram[7226]), .B2(n1917), 
        .ZN(n11467) );
  MOAI22 U20389 ( .A1(n28452), .A2(n1916), .B1(ram[7227]), .B2(n1917), 
        .ZN(n11468) );
  MOAI22 U20390 ( .A1(n28217), .A2(n1916), .B1(ram[7228]), .B2(n1917), 
        .ZN(n11469) );
  MOAI22 U20391 ( .A1(n27982), .A2(n1916), .B1(ram[7229]), .B2(n1917), 
        .ZN(n11470) );
  MOAI22 U20392 ( .A1(n27747), .A2(n1916), .B1(ram[7230]), .B2(n1917), 
        .ZN(n11471) );
  MOAI22 U20393 ( .A1(n27512), .A2(n1916), .B1(ram[7231]), .B2(n1917), 
        .ZN(n11472) );
  MOAI22 U20394 ( .A1(n29157), .A2(n1918), .B1(ram[7232]), .B2(n1919), 
        .ZN(n11473) );
  MOAI22 U20395 ( .A1(n28922), .A2(n1918), .B1(ram[7233]), .B2(n1919), 
        .ZN(n11474) );
  MOAI22 U20396 ( .A1(n28687), .A2(n1918), .B1(ram[7234]), .B2(n1919), 
        .ZN(n11475) );
  MOAI22 U20397 ( .A1(n28452), .A2(n1918), .B1(ram[7235]), .B2(n1919), 
        .ZN(n11476) );
  MOAI22 U20398 ( .A1(n28217), .A2(n1918), .B1(ram[7236]), .B2(n1919), 
        .ZN(n11477) );
  MOAI22 U20399 ( .A1(n27982), .A2(n1918), .B1(ram[7237]), .B2(n1919), 
        .ZN(n11478) );
  MOAI22 U20400 ( .A1(n27747), .A2(n1918), .B1(ram[7238]), .B2(n1919), 
        .ZN(n11479) );
  MOAI22 U20401 ( .A1(n27512), .A2(n1918), .B1(ram[7239]), .B2(n1919), 
        .ZN(n11480) );
  MOAI22 U20402 ( .A1(n29157), .A2(n1920), .B1(ram[7240]), .B2(n1921), 
        .ZN(n11481) );
  MOAI22 U20403 ( .A1(n28922), .A2(n1920), .B1(ram[7241]), .B2(n1921), 
        .ZN(n11482) );
  MOAI22 U20404 ( .A1(n28687), .A2(n1920), .B1(ram[7242]), .B2(n1921), 
        .ZN(n11483) );
  MOAI22 U20405 ( .A1(n28452), .A2(n1920), .B1(ram[7243]), .B2(n1921), 
        .ZN(n11484) );
  MOAI22 U20406 ( .A1(n28217), .A2(n1920), .B1(ram[7244]), .B2(n1921), 
        .ZN(n11485) );
  MOAI22 U20407 ( .A1(n27982), .A2(n1920), .B1(ram[7245]), .B2(n1921), 
        .ZN(n11486) );
  MOAI22 U20408 ( .A1(n27747), .A2(n1920), .B1(ram[7246]), .B2(n1921), 
        .ZN(n11487) );
  MOAI22 U20409 ( .A1(n27512), .A2(n1920), .B1(ram[7247]), .B2(n1921), 
        .ZN(n11488) );
  MOAI22 U20410 ( .A1(n29157), .A2(n1922), .B1(ram[7248]), .B2(n1923), 
        .ZN(n11489) );
  MOAI22 U20411 ( .A1(n28922), .A2(n1922), .B1(ram[7249]), .B2(n1923), 
        .ZN(n11490) );
  MOAI22 U20412 ( .A1(n28687), .A2(n1922), .B1(ram[7250]), .B2(n1923), 
        .ZN(n11491) );
  MOAI22 U20413 ( .A1(n28452), .A2(n1922), .B1(ram[7251]), .B2(n1923), 
        .ZN(n11492) );
  MOAI22 U20414 ( .A1(n28217), .A2(n1922), .B1(ram[7252]), .B2(n1923), 
        .ZN(n11493) );
  MOAI22 U20415 ( .A1(n27982), .A2(n1922), .B1(ram[7253]), .B2(n1923), 
        .ZN(n11494) );
  MOAI22 U20416 ( .A1(n27747), .A2(n1922), .B1(ram[7254]), .B2(n1923), 
        .ZN(n11495) );
  MOAI22 U20417 ( .A1(n27512), .A2(n1922), .B1(ram[7255]), .B2(n1923), 
        .ZN(n11496) );
  MOAI22 U20418 ( .A1(n29157), .A2(n1924), .B1(ram[7256]), .B2(n1925), 
        .ZN(n11497) );
  MOAI22 U20419 ( .A1(n28922), .A2(n1924), .B1(ram[7257]), .B2(n1925), 
        .ZN(n11498) );
  MOAI22 U20420 ( .A1(n28687), .A2(n1924), .B1(ram[7258]), .B2(n1925), 
        .ZN(n11499) );
  MOAI22 U20421 ( .A1(n28452), .A2(n1924), .B1(ram[7259]), .B2(n1925), 
        .ZN(n11500) );
  MOAI22 U20422 ( .A1(n28217), .A2(n1924), .B1(ram[7260]), .B2(n1925), 
        .ZN(n11501) );
  MOAI22 U20423 ( .A1(n27982), .A2(n1924), .B1(ram[7261]), .B2(n1925), 
        .ZN(n11502) );
  MOAI22 U20424 ( .A1(n27747), .A2(n1924), .B1(ram[7262]), .B2(n1925), 
        .ZN(n11503) );
  MOAI22 U20425 ( .A1(n27512), .A2(n1924), .B1(ram[7263]), .B2(n1925), 
        .ZN(n11504) );
  MOAI22 U20426 ( .A1(n29157), .A2(n1926), .B1(ram[7264]), .B2(n1927), 
        .ZN(n11505) );
  MOAI22 U20427 ( .A1(n28922), .A2(n1926), .B1(ram[7265]), .B2(n1927), 
        .ZN(n11506) );
  MOAI22 U20428 ( .A1(n28687), .A2(n1926), .B1(ram[7266]), .B2(n1927), 
        .ZN(n11507) );
  MOAI22 U20429 ( .A1(n28452), .A2(n1926), .B1(ram[7267]), .B2(n1927), 
        .ZN(n11508) );
  MOAI22 U20430 ( .A1(n28217), .A2(n1926), .B1(ram[7268]), .B2(n1927), 
        .ZN(n11509) );
  MOAI22 U20431 ( .A1(n27982), .A2(n1926), .B1(ram[7269]), .B2(n1927), 
        .ZN(n11510) );
  MOAI22 U20432 ( .A1(n27747), .A2(n1926), .B1(ram[7270]), .B2(n1927), 
        .ZN(n11511) );
  MOAI22 U20433 ( .A1(n27512), .A2(n1926), .B1(ram[7271]), .B2(n1927), 
        .ZN(n11512) );
  MOAI22 U20434 ( .A1(n29157), .A2(n1928), .B1(ram[7272]), .B2(n1929), 
        .ZN(n11513) );
  MOAI22 U20435 ( .A1(n28922), .A2(n1928), .B1(ram[7273]), .B2(n1929), 
        .ZN(n11514) );
  MOAI22 U20436 ( .A1(n28687), .A2(n1928), .B1(ram[7274]), .B2(n1929), 
        .ZN(n11515) );
  MOAI22 U20437 ( .A1(n28452), .A2(n1928), .B1(ram[7275]), .B2(n1929), 
        .ZN(n11516) );
  MOAI22 U20438 ( .A1(n28217), .A2(n1928), .B1(ram[7276]), .B2(n1929), 
        .ZN(n11517) );
  MOAI22 U20439 ( .A1(n27982), .A2(n1928), .B1(ram[7277]), .B2(n1929), 
        .ZN(n11518) );
  MOAI22 U20440 ( .A1(n27747), .A2(n1928), .B1(ram[7278]), .B2(n1929), 
        .ZN(n11519) );
  MOAI22 U20441 ( .A1(n27512), .A2(n1928), .B1(ram[7279]), .B2(n1929), 
        .ZN(n11520) );
  MOAI22 U20442 ( .A1(n29158), .A2(n1930), .B1(ram[7280]), .B2(n1931), 
        .ZN(n11521) );
  MOAI22 U20443 ( .A1(n28923), .A2(n1930), .B1(ram[7281]), .B2(n1931), 
        .ZN(n11522) );
  MOAI22 U20444 ( .A1(n28688), .A2(n1930), .B1(ram[7282]), .B2(n1931), 
        .ZN(n11523) );
  MOAI22 U20445 ( .A1(n28453), .A2(n1930), .B1(ram[7283]), .B2(n1931), 
        .ZN(n11524) );
  MOAI22 U20446 ( .A1(n28218), .A2(n1930), .B1(ram[7284]), .B2(n1931), 
        .ZN(n11525) );
  MOAI22 U20447 ( .A1(n27983), .A2(n1930), .B1(ram[7285]), .B2(n1931), 
        .ZN(n11526) );
  MOAI22 U20448 ( .A1(n27748), .A2(n1930), .B1(ram[7286]), .B2(n1931), 
        .ZN(n11527) );
  MOAI22 U20449 ( .A1(n27513), .A2(n1930), .B1(ram[7287]), .B2(n1931), 
        .ZN(n11528) );
  MOAI22 U20450 ( .A1(n29158), .A2(n1932), .B1(ram[7288]), .B2(n1933), 
        .ZN(n11529) );
  MOAI22 U20451 ( .A1(n28923), .A2(n1932), .B1(ram[7289]), .B2(n1933), 
        .ZN(n11530) );
  MOAI22 U20452 ( .A1(n28688), .A2(n1932), .B1(ram[7290]), .B2(n1933), 
        .ZN(n11531) );
  MOAI22 U20453 ( .A1(n28453), .A2(n1932), .B1(ram[7291]), .B2(n1933), 
        .ZN(n11532) );
  MOAI22 U20454 ( .A1(n28218), .A2(n1932), .B1(ram[7292]), .B2(n1933), 
        .ZN(n11533) );
  MOAI22 U20455 ( .A1(n27983), .A2(n1932), .B1(ram[7293]), .B2(n1933), 
        .ZN(n11534) );
  MOAI22 U20456 ( .A1(n27748), .A2(n1932), .B1(ram[7294]), .B2(n1933), 
        .ZN(n11535) );
  MOAI22 U20457 ( .A1(n27513), .A2(n1932), .B1(ram[7295]), .B2(n1933), 
        .ZN(n11536) );
  MOAI22 U20458 ( .A1(n29158), .A2(n1934), .B1(ram[7296]), .B2(n1935), 
        .ZN(n11537) );
  MOAI22 U20459 ( .A1(n28923), .A2(n1934), .B1(ram[7297]), .B2(n1935), 
        .ZN(n11538) );
  MOAI22 U20460 ( .A1(n28688), .A2(n1934), .B1(ram[7298]), .B2(n1935), 
        .ZN(n11539) );
  MOAI22 U20461 ( .A1(n28453), .A2(n1934), .B1(ram[7299]), .B2(n1935), 
        .ZN(n11540) );
  MOAI22 U20462 ( .A1(n28218), .A2(n1934), .B1(ram[7300]), .B2(n1935), 
        .ZN(n11541) );
  MOAI22 U20463 ( .A1(n27983), .A2(n1934), .B1(ram[7301]), .B2(n1935), 
        .ZN(n11542) );
  MOAI22 U20464 ( .A1(n27748), .A2(n1934), .B1(ram[7302]), .B2(n1935), 
        .ZN(n11543) );
  MOAI22 U20465 ( .A1(n27513), .A2(n1934), .B1(ram[7303]), .B2(n1935), 
        .ZN(n11544) );
  MOAI22 U20466 ( .A1(n29158), .A2(n1936), .B1(ram[7304]), .B2(n1937), 
        .ZN(n11545) );
  MOAI22 U20467 ( .A1(n28923), .A2(n1936), .B1(ram[7305]), .B2(n1937), 
        .ZN(n11546) );
  MOAI22 U20468 ( .A1(n28688), .A2(n1936), .B1(ram[7306]), .B2(n1937), 
        .ZN(n11547) );
  MOAI22 U20469 ( .A1(n28453), .A2(n1936), .B1(ram[7307]), .B2(n1937), 
        .ZN(n11548) );
  MOAI22 U20470 ( .A1(n28218), .A2(n1936), .B1(ram[7308]), .B2(n1937), 
        .ZN(n11549) );
  MOAI22 U20471 ( .A1(n27983), .A2(n1936), .B1(ram[7309]), .B2(n1937), 
        .ZN(n11550) );
  MOAI22 U20472 ( .A1(n27748), .A2(n1936), .B1(ram[7310]), .B2(n1937), 
        .ZN(n11551) );
  MOAI22 U20473 ( .A1(n27513), .A2(n1936), .B1(ram[7311]), .B2(n1937), 
        .ZN(n11552) );
  MOAI22 U20474 ( .A1(n29158), .A2(n1938), .B1(ram[7312]), .B2(n1939), 
        .ZN(n11553) );
  MOAI22 U20475 ( .A1(n28923), .A2(n1938), .B1(ram[7313]), .B2(n1939), 
        .ZN(n11554) );
  MOAI22 U20476 ( .A1(n28688), .A2(n1938), .B1(ram[7314]), .B2(n1939), 
        .ZN(n11555) );
  MOAI22 U20477 ( .A1(n28453), .A2(n1938), .B1(ram[7315]), .B2(n1939), 
        .ZN(n11556) );
  MOAI22 U20478 ( .A1(n28218), .A2(n1938), .B1(ram[7316]), .B2(n1939), 
        .ZN(n11557) );
  MOAI22 U20479 ( .A1(n27983), .A2(n1938), .B1(ram[7317]), .B2(n1939), 
        .ZN(n11558) );
  MOAI22 U20480 ( .A1(n27748), .A2(n1938), .B1(ram[7318]), .B2(n1939), 
        .ZN(n11559) );
  MOAI22 U20481 ( .A1(n27513), .A2(n1938), .B1(ram[7319]), .B2(n1939), 
        .ZN(n11560) );
  MOAI22 U20482 ( .A1(n29158), .A2(n1940), .B1(ram[7320]), .B2(n1941), 
        .ZN(n11561) );
  MOAI22 U20483 ( .A1(n28923), .A2(n1940), .B1(ram[7321]), .B2(n1941), 
        .ZN(n11562) );
  MOAI22 U20484 ( .A1(n28688), .A2(n1940), .B1(ram[7322]), .B2(n1941), 
        .ZN(n11563) );
  MOAI22 U20485 ( .A1(n28453), .A2(n1940), .B1(ram[7323]), .B2(n1941), 
        .ZN(n11564) );
  MOAI22 U20486 ( .A1(n28218), .A2(n1940), .B1(ram[7324]), .B2(n1941), 
        .ZN(n11565) );
  MOAI22 U20487 ( .A1(n27983), .A2(n1940), .B1(ram[7325]), .B2(n1941), 
        .ZN(n11566) );
  MOAI22 U20488 ( .A1(n27748), .A2(n1940), .B1(ram[7326]), .B2(n1941), 
        .ZN(n11567) );
  MOAI22 U20489 ( .A1(n27513), .A2(n1940), .B1(ram[7327]), .B2(n1941), 
        .ZN(n11568) );
  MOAI22 U20490 ( .A1(n29158), .A2(n1942), .B1(ram[7328]), .B2(n1943), 
        .ZN(n11569) );
  MOAI22 U20491 ( .A1(n28923), .A2(n1942), .B1(ram[7329]), .B2(n1943), 
        .ZN(n11570) );
  MOAI22 U20492 ( .A1(n28688), .A2(n1942), .B1(ram[7330]), .B2(n1943), 
        .ZN(n11571) );
  MOAI22 U20493 ( .A1(n28453), .A2(n1942), .B1(ram[7331]), .B2(n1943), 
        .ZN(n11572) );
  MOAI22 U20494 ( .A1(n28218), .A2(n1942), .B1(ram[7332]), .B2(n1943), 
        .ZN(n11573) );
  MOAI22 U20495 ( .A1(n27983), .A2(n1942), .B1(ram[7333]), .B2(n1943), 
        .ZN(n11574) );
  MOAI22 U20496 ( .A1(n27748), .A2(n1942), .B1(ram[7334]), .B2(n1943), 
        .ZN(n11575) );
  MOAI22 U20497 ( .A1(n27513), .A2(n1942), .B1(ram[7335]), .B2(n1943), 
        .ZN(n11576) );
  MOAI22 U20498 ( .A1(n29158), .A2(n1944), .B1(ram[7336]), .B2(n1945), 
        .ZN(n11577) );
  MOAI22 U20499 ( .A1(n28923), .A2(n1944), .B1(ram[7337]), .B2(n1945), 
        .ZN(n11578) );
  MOAI22 U20500 ( .A1(n28688), .A2(n1944), .B1(ram[7338]), .B2(n1945), 
        .ZN(n11579) );
  MOAI22 U20501 ( .A1(n28453), .A2(n1944), .B1(ram[7339]), .B2(n1945), 
        .ZN(n11580) );
  MOAI22 U20502 ( .A1(n28218), .A2(n1944), .B1(ram[7340]), .B2(n1945), 
        .ZN(n11581) );
  MOAI22 U20503 ( .A1(n27983), .A2(n1944), .B1(ram[7341]), .B2(n1945), 
        .ZN(n11582) );
  MOAI22 U20504 ( .A1(n27748), .A2(n1944), .B1(ram[7342]), .B2(n1945), 
        .ZN(n11583) );
  MOAI22 U20505 ( .A1(n27513), .A2(n1944), .B1(ram[7343]), .B2(n1945), 
        .ZN(n11584) );
  MOAI22 U20506 ( .A1(n29158), .A2(n1946), .B1(ram[7344]), .B2(n1947), 
        .ZN(n11585) );
  MOAI22 U20507 ( .A1(n28923), .A2(n1946), .B1(ram[7345]), .B2(n1947), 
        .ZN(n11586) );
  MOAI22 U20508 ( .A1(n28688), .A2(n1946), .B1(ram[7346]), .B2(n1947), 
        .ZN(n11587) );
  MOAI22 U20509 ( .A1(n28453), .A2(n1946), .B1(ram[7347]), .B2(n1947), 
        .ZN(n11588) );
  MOAI22 U20510 ( .A1(n28218), .A2(n1946), .B1(ram[7348]), .B2(n1947), 
        .ZN(n11589) );
  MOAI22 U20511 ( .A1(n27983), .A2(n1946), .B1(ram[7349]), .B2(n1947), 
        .ZN(n11590) );
  MOAI22 U20512 ( .A1(n27748), .A2(n1946), .B1(ram[7350]), .B2(n1947), 
        .ZN(n11591) );
  MOAI22 U20513 ( .A1(n27513), .A2(n1946), .B1(ram[7351]), .B2(n1947), 
        .ZN(n11592) );
  MOAI22 U20514 ( .A1(n29158), .A2(n1948), .B1(ram[7352]), .B2(n1949), 
        .ZN(n11593) );
  MOAI22 U20515 ( .A1(n28923), .A2(n1948), .B1(ram[7353]), .B2(n1949), 
        .ZN(n11594) );
  MOAI22 U20516 ( .A1(n28688), .A2(n1948), .B1(ram[7354]), .B2(n1949), 
        .ZN(n11595) );
  MOAI22 U20517 ( .A1(n28453), .A2(n1948), .B1(ram[7355]), .B2(n1949), 
        .ZN(n11596) );
  MOAI22 U20518 ( .A1(n28218), .A2(n1948), .B1(ram[7356]), .B2(n1949), 
        .ZN(n11597) );
  MOAI22 U20519 ( .A1(n27983), .A2(n1948), .B1(ram[7357]), .B2(n1949), 
        .ZN(n11598) );
  MOAI22 U20520 ( .A1(n27748), .A2(n1948), .B1(ram[7358]), .B2(n1949), 
        .ZN(n11599) );
  MOAI22 U20521 ( .A1(n27513), .A2(n1948), .B1(ram[7359]), .B2(n1949), 
        .ZN(n11600) );
  MOAI22 U20522 ( .A1(n29158), .A2(n1950), .B1(ram[7360]), .B2(n1951), 
        .ZN(n11601) );
  MOAI22 U20523 ( .A1(n28923), .A2(n1950), .B1(ram[7361]), .B2(n1951), 
        .ZN(n11602) );
  MOAI22 U20524 ( .A1(n28688), .A2(n1950), .B1(ram[7362]), .B2(n1951), 
        .ZN(n11603) );
  MOAI22 U20525 ( .A1(n28453), .A2(n1950), .B1(ram[7363]), .B2(n1951), 
        .ZN(n11604) );
  MOAI22 U20526 ( .A1(n28218), .A2(n1950), .B1(ram[7364]), .B2(n1951), 
        .ZN(n11605) );
  MOAI22 U20527 ( .A1(n27983), .A2(n1950), .B1(ram[7365]), .B2(n1951), 
        .ZN(n11606) );
  MOAI22 U20528 ( .A1(n27748), .A2(n1950), .B1(ram[7366]), .B2(n1951), 
        .ZN(n11607) );
  MOAI22 U20529 ( .A1(n27513), .A2(n1950), .B1(ram[7367]), .B2(n1951), 
        .ZN(n11608) );
  MOAI22 U20530 ( .A1(n29158), .A2(n1952), .B1(ram[7368]), .B2(n1953), 
        .ZN(n11609) );
  MOAI22 U20531 ( .A1(n28923), .A2(n1952), .B1(ram[7369]), .B2(n1953), 
        .ZN(n11610) );
  MOAI22 U20532 ( .A1(n28688), .A2(n1952), .B1(ram[7370]), .B2(n1953), 
        .ZN(n11611) );
  MOAI22 U20533 ( .A1(n28453), .A2(n1952), .B1(ram[7371]), .B2(n1953), 
        .ZN(n11612) );
  MOAI22 U20534 ( .A1(n28218), .A2(n1952), .B1(ram[7372]), .B2(n1953), 
        .ZN(n11613) );
  MOAI22 U20535 ( .A1(n27983), .A2(n1952), .B1(ram[7373]), .B2(n1953), 
        .ZN(n11614) );
  MOAI22 U20536 ( .A1(n27748), .A2(n1952), .B1(ram[7374]), .B2(n1953), 
        .ZN(n11615) );
  MOAI22 U20537 ( .A1(n27513), .A2(n1952), .B1(ram[7375]), .B2(n1953), 
        .ZN(n11616) );
  MOAI22 U20538 ( .A1(n29158), .A2(n1954), .B1(ram[7376]), .B2(n1955), 
        .ZN(n11617) );
  MOAI22 U20539 ( .A1(n28923), .A2(n1954), .B1(ram[7377]), .B2(n1955), 
        .ZN(n11618) );
  MOAI22 U20540 ( .A1(n28688), .A2(n1954), .B1(ram[7378]), .B2(n1955), 
        .ZN(n11619) );
  MOAI22 U20541 ( .A1(n28453), .A2(n1954), .B1(ram[7379]), .B2(n1955), 
        .ZN(n11620) );
  MOAI22 U20542 ( .A1(n28218), .A2(n1954), .B1(ram[7380]), .B2(n1955), 
        .ZN(n11621) );
  MOAI22 U20543 ( .A1(n27983), .A2(n1954), .B1(ram[7381]), .B2(n1955), 
        .ZN(n11622) );
  MOAI22 U20544 ( .A1(n27748), .A2(n1954), .B1(ram[7382]), .B2(n1955), 
        .ZN(n11623) );
  MOAI22 U20545 ( .A1(n27513), .A2(n1954), .B1(ram[7383]), .B2(n1955), 
        .ZN(n11624) );
  MOAI22 U20546 ( .A1(n29159), .A2(n1956), .B1(ram[7384]), .B2(n1957), 
        .ZN(n11625) );
  MOAI22 U20547 ( .A1(n28924), .A2(n1956), .B1(ram[7385]), .B2(n1957), 
        .ZN(n11626) );
  MOAI22 U20548 ( .A1(n28689), .A2(n1956), .B1(ram[7386]), .B2(n1957), 
        .ZN(n11627) );
  MOAI22 U20549 ( .A1(n28454), .A2(n1956), .B1(ram[7387]), .B2(n1957), 
        .ZN(n11628) );
  MOAI22 U20550 ( .A1(n28219), .A2(n1956), .B1(ram[7388]), .B2(n1957), 
        .ZN(n11629) );
  MOAI22 U20551 ( .A1(n27984), .A2(n1956), .B1(ram[7389]), .B2(n1957), 
        .ZN(n11630) );
  MOAI22 U20552 ( .A1(n27749), .A2(n1956), .B1(ram[7390]), .B2(n1957), 
        .ZN(n11631) );
  MOAI22 U20553 ( .A1(n27514), .A2(n1956), .B1(ram[7391]), .B2(n1957), 
        .ZN(n11632) );
  MOAI22 U20554 ( .A1(n29159), .A2(n1958), .B1(ram[7392]), .B2(n1959), 
        .ZN(n11633) );
  MOAI22 U20555 ( .A1(n28924), .A2(n1958), .B1(ram[7393]), .B2(n1959), 
        .ZN(n11634) );
  MOAI22 U20556 ( .A1(n28689), .A2(n1958), .B1(ram[7394]), .B2(n1959), 
        .ZN(n11635) );
  MOAI22 U20557 ( .A1(n28454), .A2(n1958), .B1(ram[7395]), .B2(n1959), 
        .ZN(n11636) );
  MOAI22 U20558 ( .A1(n28219), .A2(n1958), .B1(ram[7396]), .B2(n1959), 
        .ZN(n11637) );
  MOAI22 U20559 ( .A1(n27984), .A2(n1958), .B1(ram[7397]), .B2(n1959), 
        .ZN(n11638) );
  MOAI22 U20560 ( .A1(n27749), .A2(n1958), .B1(ram[7398]), .B2(n1959), 
        .ZN(n11639) );
  MOAI22 U20561 ( .A1(n27514), .A2(n1958), .B1(ram[7399]), .B2(n1959), 
        .ZN(n11640) );
  MOAI22 U20562 ( .A1(n29159), .A2(n1960), .B1(ram[7400]), .B2(n1961), 
        .ZN(n11641) );
  MOAI22 U20563 ( .A1(n28924), .A2(n1960), .B1(ram[7401]), .B2(n1961), 
        .ZN(n11642) );
  MOAI22 U20564 ( .A1(n28689), .A2(n1960), .B1(ram[7402]), .B2(n1961), 
        .ZN(n11643) );
  MOAI22 U20565 ( .A1(n28454), .A2(n1960), .B1(ram[7403]), .B2(n1961), 
        .ZN(n11644) );
  MOAI22 U20566 ( .A1(n28219), .A2(n1960), .B1(ram[7404]), .B2(n1961), 
        .ZN(n11645) );
  MOAI22 U20567 ( .A1(n27984), .A2(n1960), .B1(ram[7405]), .B2(n1961), 
        .ZN(n11646) );
  MOAI22 U20568 ( .A1(n27749), .A2(n1960), .B1(ram[7406]), .B2(n1961), 
        .ZN(n11647) );
  MOAI22 U20569 ( .A1(n27514), .A2(n1960), .B1(ram[7407]), .B2(n1961), 
        .ZN(n11648) );
  MOAI22 U20570 ( .A1(n29159), .A2(n1962), .B1(ram[7408]), .B2(n1963), 
        .ZN(n11649) );
  MOAI22 U20571 ( .A1(n28924), .A2(n1962), .B1(ram[7409]), .B2(n1963), 
        .ZN(n11650) );
  MOAI22 U20572 ( .A1(n28689), .A2(n1962), .B1(ram[7410]), .B2(n1963), 
        .ZN(n11651) );
  MOAI22 U20573 ( .A1(n28454), .A2(n1962), .B1(ram[7411]), .B2(n1963), 
        .ZN(n11652) );
  MOAI22 U20574 ( .A1(n28219), .A2(n1962), .B1(ram[7412]), .B2(n1963), 
        .ZN(n11653) );
  MOAI22 U20575 ( .A1(n27984), .A2(n1962), .B1(ram[7413]), .B2(n1963), 
        .ZN(n11654) );
  MOAI22 U20576 ( .A1(n27749), .A2(n1962), .B1(ram[7414]), .B2(n1963), 
        .ZN(n11655) );
  MOAI22 U20577 ( .A1(n27514), .A2(n1962), .B1(ram[7415]), .B2(n1963), 
        .ZN(n11656) );
  MOAI22 U20578 ( .A1(n29159), .A2(n1964), .B1(ram[7416]), .B2(n1965), 
        .ZN(n11657) );
  MOAI22 U20579 ( .A1(n28924), .A2(n1964), .B1(ram[7417]), .B2(n1965), 
        .ZN(n11658) );
  MOAI22 U20580 ( .A1(n28689), .A2(n1964), .B1(ram[7418]), .B2(n1965), 
        .ZN(n11659) );
  MOAI22 U20581 ( .A1(n28454), .A2(n1964), .B1(ram[7419]), .B2(n1965), 
        .ZN(n11660) );
  MOAI22 U20582 ( .A1(n28219), .A2(n1964), .B1(ram[7420]), .B2(n1965), 
        .ZN(n11661) );
  MOAI22 U20583 ( .A1(n27984), .A2(n1964), .B1(ram[7421]), .B2(n1965), 
        .ZN(n11662) );
  MOAI22 U20584 ( .A1(n27749), .A2(n1964), .B1(ram[7422]), .B2(n1965), 
        .ZN(n11663) );
  MOAI22 U20585 ( .A1(n27514), .A2(n1964), .B1(ram[7423]), .B2(n1965), 
        .ZN(n11664) );
  MOAI22 U20586 ( .A1(n29159), .A2(n1966), .B1(ram[7424]), .B2(n1967), 
        .ZN(n11665) );
  MOAI22 U20587 ( .A1(n28924), .A2(n1966), .B1(ram[7425]), .B2(n1967), 
        .ZN(n11666) );
  MOAI22 U20588 ( .A1(n28689), .A2(n1966), .B1(ram[7426]), .B2(n1967), 
        .ZN(n11667) );
  MOAI22 U20589 ( .A1(n28454), .A2(n1966), .B1(ram[7427]), .B2(n1967), 
        .ZN(n11668) );
  MOAI22 U20590 ( .A1(n28219), .A2(n1966), .B1(ram[7428]), .B2(n1967), 
        .ZN(n11669) );
  MOAI22 U20591 ( .A1(n27984), .A2(n1966), .B1(ram[7429]), .B2(n1967), 
        .ZN(n11670) );
  MOAI22 U20592 ( .A1(n27749), .A2(n1966), .B1(ram[7430]), .B2(n1967), 
        .ZN(n11671) );
  MOAI22 U20593 ( .A1(n27514), .A2(n1966), .B1(ram[7431]), .B2(n1967), 
        .ZN(n11672) );
  MOAI22 U20594 ( .A1(n29159), .A2(n1968), .B1(ram[7432]), .B2(n1969), 
        .ZN(n11673) );
  MOAI22 U20595 ( .A1(n28924), .A2(n1968), .B1(ram[7433]), .B2(n1969), 
        .ZN(n11674) );
  MOAI22 U20596 ( .A1(n28689), .A2(n1968), .B1(ram[7434]), .B2(n1969), 
        .ZN(n11675) );
  MOAI22 U20597 ( .A1(n28454), .A2(n1968), .B1(ram[7435]), .B2(n1969), 
        .ZN(n11676) );
  MOAI22 U20598 ( .A1(n28219), .A2(n1968), .B1(ram[7436]), .B2(n1969), 
        .ZN(n11677) );
  MOAI22 U20599 ( .A1(n27984), .A2(n1968), .B1(ram[7437]), .B2(n1969), 
        .ZN(n11678) );
  MOAI22 U20600 ( .A1(n27749), .A2(n1968), .B1(ram[7438]), .B2(n1969), 
        .ZN(n11679) );
  MOAI22 U20601 ( .A1(n27514), .A2(n1968), .B1(ram[7439]), .B2(n1969), 
        .ZN(n11680) );
  MOAI22 U20602 ( .A1(n29159), .A2(n1970), .B1(ram[7440]), .B2(n1971), 
        .ZN(n11681) );
  MOAI22 U20603 ( .A1(n28924), .A2(n1970), .B1(ram[7441]), .B2(n1971), 
        .ZN(n11682) );
  MOAI22 U20604 ( .A1(n28689), .A2(n1970), .B1(ram[7442]), .B2(n1971), 
        .ZN(n11683) );
  MOAI22 U20605 ( .A1(n28454), .A2(n1970), .B1(ram[7443]), .B2(n1971), 
        .ZN(n11684) );
  MOAI22 U20606 ( .A1(n28219), .A2(n1970), .B1(ram[7444]), .B2(n1971), 
        .ZN(n11685) );
  MOAI22 U20607 ( .A1(n27984), .A2(n1970), .B1(ram[7445]), .B2(n1971), 
        .ZN(n11686) );
  MOAI22 U20608 ( .A1(n27749), .A2(n1970), .B1(ram[7446]), .B2(n1971), 
        .ZN(n11687) );
  MOAI22 U20609 ( .A1(n27514), .A2(n1970), .B1(ram[7447]), .B2(n1971), 
        .ZN(n11688) );
  MOAI22 U20610 ( .A1(n29159), .A2(n1972), .B1(ram[7448]), .B2(n1973), 
        .ZN(n11689) );
  MOAI22 U20611 ( .A1(n28924), .A2(n1972), .B1(ram[7449]), .B2(n1973), 
        .ZN(n11690) );
  MOAI22 U20612 ( .A1(n28689), .A2(n1972), .B1(ram[7450]), .B2(n1973), 
        .ZN(n11691) );
  MOAI22 U20613 ( .A1(n28454), .A2(n1972), .B1(ram[7451]), .B2(n1973), 
        .ZN(n11692) );
  MOAI22 U20614 ( .A1(n28219), .A2(n1972), .B1(ram[7452]), .B2(n1973), 
        .ZN(n11693) );
  MOAI22 U20615 ( .A1(n27984), .A2(n1972), .B1(ram[7453]), .B2(n1973), 
        .ZN(n11694) );
  MOAI22 U20616 ( .A1(n27749), .A2(n1972), .B1(ram[7454]), .B2(n1973), 
        .ZN(n11695) );
  MOAI22 U20617 ( .A1(n27514), .A2(n1972), .B1(ram[7455]), .B2(n1973), 
        .ZN(n11696) );
  MOAI22 U20618 ( .A1(n29159), .A2(n1974), .B1(ram[7456]), .B2(n1975), 
        .ZN(n11697) );
  MOAI22 U20619 ( .A1(n28924), .A2(n1974), .B1(ram[7457]), .B2(n1975), 
        .ZN(n11698) );
  MOAI22 U20620 ( .A1(n28689), .A2(n1974), .B1(ram[7458]), .B2(n1975), 
        .ZN(n11699) );
  MOAI22 U20621 ( .A1(n28454), .A2(n1974), .B1(ram[7459]), .B2(n1975), 
        .ZN(n11700) );
  MOAI22 U20622 ( .A1(n28219), .A2(n1974), .B1(ram[7460]), .B2(n1975), 
        .ZN(n11701) );
  MOAI22 U20623 ( .A1(n27984), .A2(n1974), .B1(ram[7461]), .B2(n1975), 
        .ZN(n11702) );
  MOAI22 U20624 ( .A1(n27749), .A2(n1974), .B1(ram[7462]), .B2(n1975), 
        .ZN(n11703) );
  MOAI22 U20625 ( .A1(n27514), .A2(n1974), .B1(ram[7463]), .B2(n1975), 
        .ZN(n11704) );
  MOAI22 U20626 ( .A1(n29159), .A2(n1976), .B1(ram[7464]), .B2(n1977), 
        .ZN(n11705) );
  MOAI22 U20627 ( .A1(n28924), .A2(n1976), .B1(ram[7465]), .B2(n1977), 
        .ZN(n11706) );
  MOAI22 U20628 ( .A1(n28689), .A2(n1976), .B1(ram[7466]), .B2(n1977), 
        .ZN(n11707) );
  MOAI22 U20629 ( .A1(n28454), .A2(n1976), .B1(ram[7467]), .B2(n1977), 
        .ZN(n11708) );
  MOAI22 U20630 ( .A1(n28219), .A2(n1976), .B1(ram[7468]), .B2(n1977), 
        .ZN(n11709) );
  MOAI22 U20631 ( .A1(n27984), .A2(n1976), .B1(ram[7469]), .B2(n1977), 
        .ZN(n11710) );
  MOAI22 U20632 ( .A1(n27749), .A2(n1976), .B1(ram[7470]), .B2(n1977), 
        .ZN(n11711) );
  MOAI22 U20633 ( .A1(n27514), .A2(n1976), .B1(ram[7471]), .B2(n1977), 
        .ZN(n11712) );
  MOAI22 U20634 ( .A1(n29159), .A2(n1978), .B1(ram[7472]), .B2(n1979), 
        .ZN(n11713) );
  MOAI22 U20635 ( .A1(n28924), .A2(n1978), .B1(ram[7473]), .B2(n1979), 
        .ZN(n11714) );
  MOAI22 U20636 ( .A1(n28689), .A2(n1978), .B1(ram[7474]), .B2(n1979), 
        .ZN(n11715) );
  MOAI22 U20637 ( .A1(n28454), .A2(n1978), .B1(ram[7475]), .B2(n1979), 
        .ZN(n11716) );
  MOAI22 U20638 ( .A1(n28219), .A2(n1978), .B1(ram[7476]), .B2(n1979), 
        .ZN(n11717) );
  MOAI22 U20639 ( .A1(n27984), .A2(n1978), .B1(ram[7477]), .B2(n1979), 
        .ZN(n11718) );
  MOAI22 U20640 ( .A1(n27749), .A2(n1978), .B1(ram[7478]), .B2(n1979), 
        .ZN(n11719) );
  MOAI22 U20641 ( .A1(n27514), .A2(n1978), .B1(ram[7479]), .B2(n1979), 
        .ZN(n11720) );
  MOAI22 U20642 ( .A1(n29159), .A2(n1980), .B1(ram[7480]), .B2(n1981), 
        .ZN(n11721) );
  MOAI22 U20643 ( .A1(n28924), .A2(n1980), .B1(ram[7481]), .B2(n1981), 
        .ZN(n11722) );
  MOAI22 U20644 ( .A1(n28689), .A2(n1980), .B1(ram[7482]), .B2(n1981), 
        .ZN(n11723) );
  MOAI22 U20645 ( .A1(n28454), .A2(n1980), .B1(ram[7483]), .B2(n1981), 
        .ZN(n11724) );
  MOAI22 U20646 ( .A1(n28219), .A2(n1980), .B1(ram[7484]), .B2(n1981), 
        .ZN(n11725) );
  MOAI22 U20647 ( .A1(n27984), .A2(n1980), .B1(ram[7485]), .B2(n1981), 
        .ZN(n11726) );
  MOAI22 U20648 ( .A1(n27749), .A2(n1980), .B1(ram[7486]), .B2(n1981), 
        .ZN(n11727) );
  MOAI22 U20649 ( .A1(n27514), .A2(n1980), .B1(ram[7487]), .B2(n1981), 
        .ZN(n11728) );
  MOAI22 U20650 ( .A1(n29160), .A2(n1982), .B1(ram[7488]), .B2(n1983), 
        .ZN(n11729) );
  MOAI22 U20651 ( .A1(n28925), .A2(n1982), .B1(ram[7489]), .B2(n1983), 
        .ZN(n11730) );
  MOAI22 U20652 ( .A1(n28690), .A2(n1982), .B1(ram[7490]), .B2(n1983), 
        .ZN(n11731) );
  MOAI22 U20653 ( .A1(n28455), .A2(n1982), .B1(ram[7491]), .B2(n1983), 
        .ZN(n11732) );
  MOAI22 U20654 ( .A1(n28220), .A2(n1982), .B1(ram[7492]), .B2(n1983), 
        .ZN(n11733) );
  MOAI22 U20655 ( .A1(n27985), .A2(n1982), .B1(ram[7493]), .B2(n1983), 
        .ZN(n11734) );
  MOAI22 U20656 ( .A1(n27750), .A2(n1982), .B1(ram[7494]), .B2(n1983), 
        .ZN(n11735) );
  MOAI22 U20657 ( .A1(n27515), .A2(n1982), .B1(ram[7495]), .B2(n1983), 
        .ZN(n11736) );
  MOAI22 U20658 ( .A1(n29160), .A2(n1984), .B1(ram[7496]), .B2(n1985), 
        .ZN(n11737) );
  MOAI22 U20659 ( .A1(n28925), .A2(n1984), .B1(ram[7497]), .B2(n1985), 
        .ZN(n11738) );
  MOAI22 U20660 ( .A1(n28690), .A2(n1984), .B1(ram[7498]), .B2(n1985), 
        .ZN(n11739) );
  MOAI22 U20661 ( .A1(n28455), .A2(n1984), .B1(ram[7499]), .B2(n1985), 
        .ZN(n11740) );
  MOAI22 U20662 ( .A1(n28220), .A2(n1984), .B1(ram[7500]), .B2(n1985), 
        .ZN(n11741) );
  MOAI22 U20663 ( .A1(n27985), .A2(n1984), .B1(ram[7501]), .B2(n1985), 
        .ZN(n11742) );
  MOAI22 U20664 ( .A1(n27750), .A2(n1984), .B1(ram[7502]), .B2(n1985), 
        .ZN(n11743) );
  MOAI22 U20665 ( .A1(n27515), .A2(n1984), .B1(ram[7503]), .B2(n1985), 
        .ZN(n11744) );
  MOAI22 U20666 ( .A1(n29160), .A2(n1986), .B1(ram[7504]), .B2(n1987), 
        .ZN(n11745) );
  MOAI22 U20667 ( .A1(n28925), .A2(n1986), .B1(ram[7505]), .B2(n1987), 
        .ZN(n11746) );
  MOAI22 U20668 ( .A1(n28690), .A2(n1986), .B1(ram[7506]), .B2(n1987), 
        .ZN(n11747) );
  MOAI22 U20669 ( .A1(n28455), .A2(n1986), .B1(ram[7507]), .B2(n1987), 
        .ZN(n11748) );
  MOAI22 U20670 ( .A1(n28220), .A2(n1986), .B1(ram[7508]), .B2(n1987), 
        .ZN(n11749) );
  MOAI22 U20671 ( .A1(n27985), .A2(n1986), .B1(ram[7509]), .B2(n1987), 
        .ZN(n11750) );
  MOAI22 U20672 ( .A1(n27750), .A2(n1986), .B1(ram[7510]), .B2(n1987), 
        .ZN(n11751) );
  MOAI22 U20673 ( .A1(n27515), .A2(n1986), .B1(ram[7511]), .B2(n1987), 
        .ZN(n11752) );
  MOAI22 U20674 ( .A1(n29160), .A2(n1988), .B1(ram[7512]), .B2(n1989), 
        .ZN(n11753) );
  MOAI22 U20675 ( .A1(n28925), .A2(n1988), .B1(ram[7513]), .B2(n1989), 
        .ZN(n11754) );
  MOAI22 U20676 ( .A1(n28690), .A2(n1988), .B1(ram[7514]), .B2(n1989), 
        .ZN(n11755) );
  MOAI22 U20677 ( .A1(n28455), .A2(n1988), .B1(ram[7515]), .B2(n1989), 
        .ZN(n11756) );
  MOAI22 U20678 ( .A1(n28220), .A2(n1988), .B1(ram[7516]), .B2(n1989), 
        .ZN(n11757) );
  MOAI22 U20679 ( .A1(n27985), .A2(n1988), .B1(ram[7517]), .B2(n1989), 
        .ZN(n11758) );
  MOAI22 U20680 ( .A1(n27750), .A2(n1988), .B1(ram[7518]), .B2(n1989), 
        .ZN(n11759) );
  MOAI22 U20681 ( .A1(n27515), .A2(n1988), .B1(ram[7519]), .B2(n1989), 
        .ZN(n11760) );
  MOAI22 U20682 ( .A1(n29160), .A2(n1990), .B1(ram[7520]), .B2(n1991), 
        .ZN(n11761) );
  MOAI22 U20683 ( .A1(n28925), .A2(n1990), .B1(ram[7521]), .B2(n1991), 
        .ZN(n11762) );
  MOAI22 U20684 ( .A1(n28690), .A2(n1990), .B1(ram[7522]), .B2(n1991), 
        .ZN(n11763) );
  MOAI22 U20685 ( .A1(n28455), .A2(n1990), .B1(ram[7523]), .B2(n1991), 
        .ZN(n11764) );
  MOAI22 U20686 ( .A1(n28220), .A2(n1990), .B1(ram[7524]), .B2(n1991), 
        .ZN(n11765) );
  MOAI22 U20687 ( .A1(n27985), .A2(n1990), .B1(ram[7525]), .B2(n1991), 
        .ZN(n11766) );
  MOAI22 U20688 ( .A1(n27750), .A2(n1990), .B1(ram[7526]), .B2(n1991), 
        .ZN(n11767) );
  MOAI22 U20689 ( .A1(n27515), .A2(n1990), .B1(ram[7527]), .B2(n1991), 
        .ZN(n11768) );
  MOAI22 U20690 ( .A1(n29160), .A2(n1992), .B1(ram[7528]), .B2(n1993), 
        .ZN(n11769) );
  MOAI22 U20691 ( .A1(n28925), .A2(n1992), .B1(ram[7529]), .B2(n1993), 
        .ZN(n11770) );
  MOAI22 U20692 ( .A1(n28690), .A2(n1992), .B1(ram[7530]), .B2(n1993), 
        .ZN(n11771) );
  MOAI22 U20693 ( .A1(n28455), .A2(n1992), .B1(ram[7531]), .B2(n1993), 
        .ZN(n11772) );
  MOAI22 U20694 ( .A1(n28220), .A2(n1992), .B1(ram[7532]), .B2(n1993), 
        .ZN(n11773) );
  MOAI22 U20695 ( .A1(n27985), .A2(n1992), .B1(ram[7533]), .B2(n1993), 
        .ZN(n11774) );
  MOAI22 U20696 ( .A1(n27750), .A2(n1992), .B1(ram[7534]), .B2(n1993), 
        .ZN(n11775) );
  MOAI22 U20697 ( .A1(n27515), .A2(n1992), .B1(ram[7535]), .B2(n1993), 
        .ZN(n11776) );
  MOAI22 U20698 ( .A1(n29160), .A2(n1994), .B1(ram[7536]), .B2(n1995), 
        .ZN(n11777) );
  MOAI22 U20699 ( .A1(n28925), .A2(n1994), .B1(ram[7537]), .B2(n1995), 
        .ZN(n11778) );
  MOAI22 U20700 ( .A1(n28690), .A2(n1994), .B1(ram[7538]), .B2(n1995), 
        .ZN(n11779) );
  MOAI22 U20701 ( .A1(n28455), .A2(n1994), .B1(ram[7539]), .B2(n1995), 
        .ZN(n11780) );
  MOAI22 U20702 ( .A1(n28220), .A2(n1994), .B1(ram[7540]), .B2(n1995), 
        .ZN(n11781) );
  MOAI22 U20703 ( .A1(n27985), .A2(n1994), .B1(ram[7541]), .B2(n1995), 
        .ZN(n11782) );
  MOAI22 U20704 ( .A1(n27750), .A2(n1994), .B1(ram[7542]), .B2(n1995), 
        .ZN(n11783) );
  MOAI22 U20705 ( .A1(n27515), .A2(n1994), .B1(ram[7543]), .B2(n1995), 
        .ZN(n11784) );
  MOAI22 U20706 ( .A1(n29160), .A2(n1996), .B1(ram[7544]), .B2(n1997), 
        .ZN(n11785) );
  MOAI22 U20707 ( .A1(n28925), .A2(n1996), .B1(ram[7545]), .B2(n1997), 
        .ZN(n11786) );
  MOAI22 U20708 ( .A1(n28690), .A2(n1996), .B1(ram[7546]), .B2(n1997), 
        .ZN(n11787) );
  MOAI22 U20709 ( .A1(n28455), .A2(n1996), .B1(ram[7547]), .B2(n1997), 
        .ZN(n11788) );
  MOAI22 U20710 ( .A1(n28220), .A2(n1996), .B1(ram[7548]), .B2(n1997), 
        .ZN(n11789) );
  MOAI22 U20711 ( .A1(n27985), .A2(n1996), .B1(ram[7549]), .B2(n1997), 
        .ZN(n11790) );
  MOAI22 U20712 ( .A1(n27750), .A2(n1996), .B1(ram[7550]), .B2(n1997), 
        .ZN(n11791) );
  MOAI22 U20713 ( .A1(n27515), .A2(n1996), .B1(ram[7551]), .B2(n1997), 
        .ZN(n11792) );
  MOAI22 U20714 ( .A1(n29160), .A2(n1998), .B1(ram[7552]), .B2(n1999), 
        .ZN(n11793) );
  MOAI22 U20715 ( .A1(n28925), .A2(n1998), .B1(ram[7553]), .B2(n1999), 
        .ZN(n11794) );
  MOAI22 U20716 ( .A1(n28690), .A2(n1998), .B1(ram[7554]), .B2(n1999), 
        .ZN(n11795) );
  MOAI22 U20717 ( .A1(n28455), .A2(n1998), .B1(ram[7555]), .B2(n1999), 
        .ZN(n11796) );
  MOAI22 U20718 ( .A1(n28220), .A2(n1998), .B1(ram[7556]), .B2(n1999), 
        .ZN(n11797) );
  MOAI22 U20719 ( .A1(n27985), .A2(n1998), .B1(ram[7557]), .B2(n1999), 
        .ZN(n11798) );
  MOAI22 U20720 ( .A1(n27750), .A2(n1998), .B1(ram[7558]), .B2(n1999), 
        .ZN(n11799) );
  MOAI22 U20721 ( .A1(n27515), .A2(n1998), .B1(ram[7559]), .B2(n1999), 
        .ZN(n11800) );
  MOAI22 U20722 ( .A1(n29160), .A2(n2000), .B1(ram[7560]), .B2(n2001), 
        .ZN(n11801) );
  MOAI22 U20723 ( .A1(n28925), .A2(n2000), .B1(ram[7561]), .B2(n2001), 
        .ZN(n11802) );
  MOAI22 U20724 ( .A1(n28690), .A2(n2000), .B1(ram[7562]), .B2(n2001), 
        .ZN(n11803) );
  MOAI22 U20725 ( .A1(n28455), .A2(n2000), .B1(ram[7563]), .B2(n2001), 
        .ZN(n11804) );
  MOAI22 U20726 ( .A1(n28220), .A2(n2000), .B1(ram[7564]), .B2(n2001), 
        .ZN(n11805) );
  MOAI22 U20727 ( .A1(n27985), .A2(n2000), .B1(ram[7565]), .B2(n2001), 
        .ZN(n11806) );
  MOAI22 U20728 ( .A1(n27750), .A2(n2000), .B1(ram[7566]), .B2(n2001), 
        .ZN(n11807) );
  MOAI22 U20729 ( .A1(n27515), .A2(n2000), .B1(ram[7567]), .B2(n2001), 
        .ZN(n11808) );
  MOAI22 U20730 ( .A1(n29160), .A2(n2002), .B1(ram[7568]), .B2(n2003), 
        .ZN(n11809) );
  MOAI22 U20731 ( .A1(n28925), .A2(n2002), .B1(ram[7569]), .B2(n2003), 
        .ZN(n11810) );
  MOAI22 U20732 ( .A1(n28690), .A2(n2002), .B1(ram[7570]), .B2(n2003), 
        .ZN(n11811) );
  MOAI22 U20733 ( .A1(n28455), .A2(n2002), .B1(ram[7571]), .B2(n2003), 
        .ZN(n11812) );
  MOAI22 U20734 ( .A1(n28220), .A2(n2002), .B1(ram[7572]), .B2(n2003), 
        .ZN(n11813) );
  MOAI22 U20735 ( .A1(n27985), .A2(n2002), .B1(ram[7573]), .B2(n2003), 
        .ZN(n11814) );
  MOAI22 U20736 ( .A1(n27750), .A2(n2002), .B1(ram[7574]), .B2(n2003), 
        .ZN(n11815) );
  MOAI22 U20737 ( .A1(n27515), .A2(n2002), .B1(ram[7575]), .B2(n2003), 
        .ZN(n11816) );
  MOAI22 U20738 ( .A1(n29160), .A2(n2004), .B1(ram[7576]), .B2(n2005), 
        .ZN(n11817) );
  MOAI22 U20739 ( .A1(n28925), .A2(n2004), .B1(ram[7577]), .B2(n2005), 
        .ZN(n11818) );
  MOAI22 U20740 ( .A1(n28690), .A2(n2004), .B1(ram[7578]), .B2(n2005), 
        .ZN(n11819) );
  MOAI22 U20741 ( .A1(n28455), .A2(n2004), .B1(ram[7579]), .B2(n2005), 
        .ZN(n11820) );
  MOAI22 U20742 ( .A1(n28220), .A2(n2004), .B1(ram[7580]), .B2(n2005), 
        .ZN(n11821) );
  MOAI22 U20743 ( .A1(n27985), .A2(n2004), .B1(ram[7581]), .B2(n2005), 
        .ZN(n11822) );
  MOAI22 U20744 ( .A1(n27750), .A2(n2004), .B1(ram[7582]), .B2(n2005), 
        .ZN(n11823) );
  MOAI22 U20745 ( .A1(n27515), .A2(n2004), .B1(ram[7583]), .B2(n2005), 
        .ZN(n11824) );
  MOAI22 U20746 ( .A1(n29160), .A2(n2006), .B1(ram[7584]), .B2(n2007), 
        .ZN(n11825) );
  MOAI22 U20747 ( .A1(n28925), .A2(n2006), .B1(ram[7585]), .B2(n2007), 
        .ZN(n11826) );
  MOAI22 U20748 ( .A1(n28690), .A2(n2006), .B1(ram[7586]), .B2(n2007), 
        .ZN(n11827) );
  MOAI22 U20749 ( .A1(n28455), .A2(n2006), .B1(ram[7587]), .B2(n2007), 
        .ZN(n11828) );
  MOAI22 U20750 ( .A1(n28220), .A2(n2006), .B1(ram[7588]), .B2(n2007), 
        .ZN(n11829) );
  MOAI22 U20751 ( .A1(n27985), .A2(n2006), .B1(ram[7589]), .B2(n2007), 
        .ZN(n11830) );
  MOAI22 U20752 ( .A1(n27750), .A2(n2006), .B1(ram[7590]), .B2(n2007), 
        .ZN(n11831) );
  MOAI22 U20753 ( .A1(n27515), .A2(n2006), .B1(ram[7591]), .B2(n2007), 
        .ZN(n11832) );
  MOAI22 U20754 ( .A1(n29161), .A2(n2008), .B1(ram[7592]), .B2(n2009), 
        .ZN(n11833) );
  MOAI22 U20755 ( .A1(n28926), .A2(n2008), .B1(ram[7593]), .B2(n2009), 
        .ZN(n11834) );
  MOAI22 U20756 ( .A1(n28691), .A2(n2008), .B1(ram[7594]), .B2(n2009), 
        .ZN(n11835) );
  MOAI22 U20757 ( .A1(n28456), .A2(n2008), .B1(ram[7595]), .B2(n2009), 
        .ZN(n11836) );
  MOAI22 U20758 ( .A1(n28221), .A2(n2008), .B1(ram[7596]), .B2(n2009), 
        .ZN(n11837) );
  MOAI22 U20759 ( .A1(n27986), .A2(n2008), .B1(ram[7597]), .B2(n2009), 
        .ZN(n11838) );
  MOAI22 U20760 ( .A1(n27751), .A2(n2008), .B1(ram[7598]), .B2(n2009), 
        .ZN(n11839) );
  MOAI22 U20761 ( .A1(n27516), .A2(n2008), .B1(ram[7599]), .B2(n2009), 
        .ZN(n11840) );
  MOAI22 U20762 ( .A1(n29161), .A2(n2010), .B1(ram[7600]), .B2(n2011), 
        .ZN(n11841) );
  MOAI22 U20763 ( .A1(n28926), .A2(n2010), .B1(ram[7601]), .B2(n2011), 
        .ZN(n11842) );
  MOAI22 U20764 ( .A1(n28691), .A2(n2010), .B1(ram[7602]), .B2(n2011), 
        .ZN(n11843) );
  MOAI22 U20765 ( .A1(n28456), .A2(n2010), .B1(ram[7603]), .B2(n2011), 
        .ZN(n11844) );
  MOAI22 U20766 ( .A1(n28221), .A2(n2010), .B1(ram[7604]), .B2(n2011), 
        .ZN(n11845) );
  MOAI22 U20767 ( .A1(n27986), .A2(n2010), .B1(ram[7605]), .B2(n2011), 
        .ZN(n11846) );
  MOAI22 U20768 ( .A1(n27751), .A2(n2010), .B1(ram[7606]), .B2(n2011), 
        .ZN(n11847) );
  MOAI22 U20769 ( .A1(n27516), .A2(n2010), .B1(ram[7607]), .B2(n2011), 
        .ZN(n11848) );
  MOAI22 U20770 ( .A1(n29161), .A2(n2012), .B1(ram[7608]), .B2(n2013), 
        .ZN(n11849) );
  MOAI22 U20771 ( .A1(n28926), .A2(n2012), .B1(ram[7609]), .B2(n2013), 
        .ZN(n11850) );
  MOAI22 U20772 ( .A1(n28691), .A2(n2012), .B1(ram[7610]), .B2(n2013), 
        .ZN(n11851) );
  MOAI22 U20773 ( .A1(n28456), .A2(n2012), .B1(ram[7611]), .B2(n2013), 
        .ZN(n11852) );
  MOAI22 U20774 ( .A1(n28221), .A2(n2012), .B1(ram[7612]), .B2(n2013), 
        .ZN(n11853) );
  MOAI22 U20775 ( .A1(n27986), .A2(n2012), .B1(ram[7613]), .B2(n2013), 
        .ZN(n11854) );
  MOAI22 U20776 ( .A1(n27751), .A2(n2012), .B1(ram[7614]), .B2(n2013), 
        .ZN(n11855) );
  MOAI22 U20777 ( .A1(n27516), .A2(n2012), .B1(ram[7615]), .B2(n2013), 
        .ZN(n11856) );
  MOAI22 U20778 ( .A1(n29161), .A2(n2014), .B1(ram[7616]), .B2(n2015), 
        .ZN(n11857) );
  MOAI22 U20779 ( .A1(n28926), .A2(n2014), .B1(ram[7617]), .B2(n2015), 
        .ZN(n11858) );
  MOAI22 U20780 ( .A1(n28691), .A2(n2014), .B1(ram[7618]), .B2(n2015), 
        .ZN(n11859) );
  MOAI22 U20781 ( .A1(n28456), .A2(n2014), .B1(ram[7619]), .B2(n2015), 
        .ZN(n11860) );
  MOAI22 U20782 ( .A1(n28221), .A2(n2014), .B1(ram[7620]), .B2(n2015), 
        .ZN(n11861) );
  MOAI22 U20783 ( .A1(n27986), .A2(n2014), .B1(ram[7621]), .B2(n2015), 
        .ZN(n11862) );
  MOAI22 U20784 ( .A1(n27751), .A2(n2014), .B1(ram[7622]), .B2(n2015), 
        .ZN(n11863) );
  MOAI22 U20785 ( .A1(n27516), .A2(n2014), .B1(ram[7623]), .B2(n2015), 
        .ZN(n11864) );
  MOAI22 U20786 ( .A1(n29161), .A2(n2016), .B1(ram[7624]), .B2(n2017), 
        .ZN(n11865) );
  MOAI22 U20787 ( .A1(n28926), .A2(n2016), .B1(ram[7625]), .B2(n2017), 
        .ZN(n11866) );
  MOAI22 U20788 ( .A1(n28691), .A2(n2016), .B1(ram[7626]), .B2(n2017), 
        .ZN(n11867) );
  MOAI22 U20789 ( .A1(n28456), .A2(n2016), .B1(ram[7627]), .B2(n2017), 
        .ZN(n11868) );
  MOAI22 U20790 ( .A1(n28221), .A2(n2016), .B1(ram[7628]), .B2(n2017), 
        .ZN(n11869) );
  MOAI22 U20791 ( .A1(n27986), .A2(n2016), .B1(ram[7629]), .B2(n2017), 
        .ZN(n11870) );
  MOAI22 U20792 ( .A1(n27751), .A2(n2016), .B1(ram[7630]), .B2(n2017), 
        .ZN(n11871) );
  MOAI22 U20793 ( .A1(n27516), .A2(n2016), .B1(ram[7631]), .B2(n2017), 
        .ZN(n11872) );
  MOAI22 U20794 ( .A1(n29161), .A2(n2018), .B1(ram[7632]), .B2(n2019), 
        .ZN(n11873) );
  MOAI22 U20795 ( .A1(n28926), .A2(n2018), .B1(ram[7633]), .B2(n2019), 
        .ZN(n11874) );
  MOAI22 U20796 ( .A1(n28691), .A2(n2018), .B1(ram[7634]), .B2(n2019), 
        .ZN(n11875) );
  MOAI22 U20797 ( .A1(n28456), .A2(n2018), .B1(ram[7635]), .B2(n2019), 
        .ZN(n11876) );
  MOAI22 U20798 ( .A1(n28221), .A2(n2018), .B1(ram[7636]), .B2(n2019), 
        .ZN(n11877) );
  MOAI22 U20799 ( .A1(n27986), .A2(n2018), .B1(ram[7637]), .B2(n2019), 
        .ZN(n11878) );
  MOAI22 U20800 ( .A1(n27751), .A2(n2018), .B1(ram[7638]), .B2(n2019), 
        .ZN(n11879) );
  MOAI22 U20801 ( .A1(n27516), .A2(n2018), .B1(ram[7639]), .B2(n2019), 
        .ZN(n11880) );
  MOAI22 U20802 ( .A1(n29161), .A2(n2020), .B1(ram[7640]), .B2(n2021), 
        .ZN(n11881) );
  MOAI22 U20803 ( .A1(n28926), .A2(n2020), .B1(ram[7641]), .B2(n2021), 
        .ZN(n11882) );
  MOAI22 U20804 ( .A1(n28691), .A2(n2020), .B1(ram[7642]), .B2(n2021), 
        .ZN(n11883) );
  MOAI22 U20805 ( .A1(n28456), .A2(n2020), .B1(ram[7643]), .B2(n2021), 
        .ZN(n11884) );
  MOAI22 U20806 ( .A1(n28221), .A2(n2020), .B1(ram[7644]), .B2(n2021), 
        .ZN(n11885) );
  MOAI22 U20807 ( .A1(n27986), .A2(n2020), .B1(ram[7645]), .B2(n2021), 
        .ZN(n11886) );
  MOAI22 U20808 ( .A1(n27751), .A2(n2020), .B1(ram[7646]), .B2(n2021), 
        .ZN(n11887) );
  MOAI22 U20809 ( .A1(n27516), .A2(n2020), .B1(ram[7647]), .B2(n2021), 
        .ZN(n11888) );
  MOAI22 U20810 ( .A1(n29161), .A2(n2022), .B1(ram[7648]), .B2(n2023), 
        .ZN(n11889) );
  MOAI22 U20811 ( .A1(n28926), .A2(n2022), .B1(ram[7649]), .B2(n2023), 
        .ZN(n11890) );
  MOAI22 U20812 ( .A1(n28691), .A2(n2022), .B1(ram[7650]), .B2(n2023), 
        .ZN(n11891) );
  MOAI22 U20813 ( .A1(n28456), .A2(n2022), .B1(ram[7651]), .B2(n2023), 
        .ZN(n11892) );
  MOAI22 U20814 ( .A1(n28221), .A2(n2022), .B1(ram[7652]), .B2(n2023), 
        .ZN(n11893) );
  MOAI22 U20815 ( .A1(n27986), .A2(n2022), .B1(ram[7653]), .B2(n2023), 
        .ZN(n11894) );
  MOAI22 U20816 ( .A1(n27751), .A2(n2022), .B1(ram[7654]), .B2(n2023), 
        .ZN(n11895) );
  MOAI22 U20817 ( .A1(n27516), .A2(n2022), .B1(ram[7655]), .B2(n2023), 
        .ZN(n11896) );
  MOAI22 U20818 ( .A1(n29161), .A2(n2024), .B1(ram[7656]), .B2(n2025), 
        .ZN(n11897) );
  MOAI22 U20819 ( .A1(n28926), .A2(n2024), .B1(ram[7657]), .B2(n2025), 
        .ZN(n11898) );
  MOAI22 U20820 ( .A1(n28691), .A2(n2024), .B1(ram[7658]), .B2(n2025), 
        .ZN(n11899) );
  MOAI22 U20821 ( .A1(n28456), .A2(n2024), .B1(ram[7659]), .B2(n2025), 
        .ZN(n11900) );
  MOAI22 U20822 ( .A1(n28221), .A2(n2024), .B1(ram[7660]), .B2(n2025), 
        .ZN(n11901) );
  MOAI22 U20823 ( .A1(n27986), .A2(n2024), .B1(ram[7661]), .B2(n2025), 
        .ZN(n11902) );
  MOAI22 U20824 ( .A1(n27751), .A2(n2024), .B1(ram[7662]), .B2(n2025), 
        .ZN(n11903) );
  MOAI22 U20825 ( .A1(n27516), .A2(n2024), .B1(ram[7663]), .B2(n2025), 
        .ZN(n11904) );
  MOAI22 U20826 ( .A1(n29161), .A2(n2026), .B1(ram[7664]), .B2(n2027), 
        .ZN(n11905) );
  MOAI22 U20827 ( .A1(n28926), .A2(n2026), .B1(ram[7665]), .B2(n2027), 
        .ZN(n11906) );
  MOAI22 U20828 ( .A1(n28691), .A2(n2026), .B1(ram[7666]), .B2(n2027), 
        .ZN(n11907) );
  MOAI22 U20829 ( .A1(n28456), .A2(n2026), .B1(ram[7667]), .B2(n2027), 
        .ZN(n11908) );
  MOAI22 U20830 ( .A1(n28221), .A2(n2026), .B1(ram[7668]), .B2(n2027), 
        .ZN(n11909) );
  MOAI22 U20831 ( .A1(n27986), .A2(n2026), .B1(ram[7669]), .B2(n2027), 
        .ZN(n11910) );
  MOAI22 U20832 ( .A1(n27751), .A2(n2026), .B1(ram[7670]), .B2(n2027), 
        .ZN(n11911) );
  MOAI22 U20833 ( .A1(n27516), .A2(n2026), .B1(ram[7671]), .B2(n2027), 
        .ZN(n11912) );
  MOAI22 U20834 ( .A1(n29161), .A2(n2028), .B1(ram[7672]), .B2(n2029), 
        .ZN(n11913) );
  MOAI22 U20835 ( .A1(n28926), .A2(n2028), .B1(ram[7673]), .B2(n2029), 
        .ZN(n11914) );
  MOAI22 U20836 ( .A1(n28691), .A2(n2028), .B1(ram[7674]), .B2(n2029), 
        .ZN(n11915) );
  MOAI22 U20837 ( .A1(n28456), .A2(n2028), .B1(ram[7675]), .B2(n2029), 
        .ZN(n11916) );
  MOAI22 U20838 ( .A1(n28221), .A2(n2028), .B1(ram[7676]), .B2(n2029), 
        .ZN(n11917) );
  MOAI22 U20839 ( .A1(n27986), .A2(n2028), .B1(ram[7677]), .B2(n2029), 
        .ZN(n11918) );
  MOAI22 U20840 ( .A1(n27751), .A2(n2028), .B1(ram[7678]), .B2(n2029), 
        .ZN(n11919) );
  MOAI22 U20841 ( .A1(n27516), .A2(n2028), .B1(ram[7679]), .B2(n2029), 
        .ZN(n11920) );
  MOAI22 U20842 ( .A1(n29161), .A2(n2030), .B1(ram[7680]), .B2(n2031), 
        .ZN(n11921) );
  MOAI22 U20843 ( .A1(n28926), .A2(n2030), .B1(ram[7681]), .B2(n2031), 
        .ZN(n11922) );
  MOAI22 U20844 ( .A1(n28691), .A2(n2030), .B1(ram[7682]), .B2(n2031), 
        .ZN(n11923) );
  MOAI22 U20845 ( .A1(n28456), .A2(n2030), .B1(ram[7683]), .B2(n2031), 
        .ZN(n11924) );
  MOAI22 U20846 ( .A1(n28221), .A2(n2030), .B1(ram[7684]), .B2(n2031), 
        .ZN(n11925) );
  MOAI22 U20847 ( .A1(n27986), .A2(n2030), .B1(ram[7685]), .B2(n2031), 
        .ZN(n11926) );
  MOAI22 U20848 ( .A1(n27751), .A2(n2030), .B1(ram[7686]), .B2(n2031), 
        .ZN(n11927) );
  MOAI22 U20849 ( .A1(n27516), .A2(n2030), .B1(ram[7687]), .B2(n2031), 
        .ZN(n11928) );
  MOAI22 U20850 ( .A1(n29161), .A2(n2033), .B1(ram[7688]), .B2(n2034), 
        .ZN(n11929) );
  MOAI22 U20851 ( .A1(n28926), .A2(n2033), .B1(ram[7689]), .B2(n2034), 
        .ZN(n11930) );
  MOAI22 U20852 ( .A1(n28691), .A2(n2033), .B1(ram[7690]), .B2(n2034), 
        .ZN(n11931) );
  MOAI22 U20853 ( .A1(n28456), .A2(n2033), .B1(ram[7691]), .B2(n2034), 
        .ZN(n11932) );
  MOAI22 U20854 ( .A1(n28221), .A2(n2033), .B1(ram[7692]), .B2(n2034), 
        .ZN(n11933) );
  MOAI22 U20855 ( .A1(n27986), .A2(n2033), .B1(ram[7693]), .B2(n2034), 
        .ZN(n11934) );
  MOAI22 U20856 ( .A1(n27751), .A2(n2033), .B1(ram[7694]), .B2(n2034), 
        .ZN(n11935) );
  MOAI22 U20857 ( .A1(n27516), .A2(n2033), .B1(ram[7695]), .B2(n2034), 
        .ZN(n11936) );
  MOAI22 U20858 ( .A1(n29162), .A2(n2035), .B1(ram[7696]), .B2(n2036), 
        .ZN(n11937) );
  MOAI22 U20859 ( .A1(n28927), .A2(n2035), .B1(ram[7697]), .B2(n2036), 
        .ZN(n11938) );
  MOAI22 U20860 ( .A1(n28692), .A2(n2035), .B1(ram[7698]), .B2(n2036), 
        .ZN(n11939) );
  MOAI22 U20861 ( .A1(n28457), .A2(n2035), .B1(ram[7699]), .B2(n2036), 
        .ZN(n11940) );
  MOAI22 U20862 ( .A1(n28222), .A2(n2035), .B1(ram[7700]), .B2(n2036), 
        .ZN(n11941) );
  MOAI22 U20863 ( .A1(n27987), .A2(n2035), .B1(ram[7701]), .B2(n2036), 
        .ZN(n11942) );
  MOAI22 U20864 ( .A1(n27752), .A2(n2035), .B1(ram[7702]), .B2(n2036), 
        .ZN(n11943) );
  MOAI22 U20865 ( .A1(n27517), .A2(n2035), .B1(ram[7703]), .B2(n2036), 
        .ZN(n11944) );
  MOAI22 U20866 ( .A1(n29162), .A2(n2037), .B1(ram[7704]), .B2(n2038), 
        .ZN(n11945) );
  MOAI22 U20867 ( .A1(n28927), .A2(n2037), .B1(ram[7705]), .B2(n2038), 
        .ZN(n11946) );
  MOAI22 U20868 ( .A1(n28692), .A2(n2037), .B1(ram[7706]), .B2(n2038), 
        .ZN(n11947) );
  MOAI22 U20869 ( .A1(n28457), .A2(n2037), .B1(ram[7707]), .B2(n2038), 
        .ZN(n11948) );
  MOAI22 U20870 ( .A1(n28222), .A2(n2037), .B1(ram[7708]), .B2(n2038), 
        .ZN(n11949) );
  MOAI22 U20871 ( .A1(n27987), .A2(n2037), .B1(ram[7709]), .B2(n2038), 
        .ZN(n11950) );
  MOAI22 U20872 ( .A1(n27752), .A2(n2037), .B1(ram[7710]), .B2(n2038), 
        .ZN(n11951) );
  MOAI22 U20873 ( .A1(n27517), .A2(n2037), .B1(ram[7711]), .B2(n2038), 
        .ZN(n11952) );
  MOAI22 U20874 ( .A1(n29162), .A2(n2039), .B1(ram[7712]), .B2(n2040), 
        .ZN(n11953) );
  MOAI22 U20875 ( .A1(n28927), .A2(n2039), .B1(ram[7713]), .B2(n2040), 
        .ZN(n11954) );
  MOAI22 U20876 ( .A1(n28692), .A2(n2039), .B1(ram[7714]), .B2(n2040), 
        .ZN(n11955) );
  MOAI22 U20877 ( .A1(n28457), .A2(n2039), .B1(ram[7715]), .B2(n2040), 
        .ZN(n11956) );
  MOAI22 U20878 ( .A1(n28222), .A2(n2039), .B1(ram[7716]), .B2(n2040), 
        .ZN(n11957) );
  MOAI22 U20879 ( .A1(n27987), .A2(n2039), .B1(ram[7717]), .B2(n2040), 
        .ZN(n11958) );
  MOAI22 U20880 ( .A1(n27752), .A2(n2039), .B1(ram[7718]), .B2(n2040), 
        .ZN(n11959) );
  MOAI22 U20881 ( .A1(n27517), .A2(n2039), .B1(ram[7719]), .B2(n2040), 
        .ZN(n11960) );
  MOAI22 U20882 ( .A1(n29162), .A2(n2041), .B1(ram[7720]), .B2(n2042), 
        .ZN(n11961) );
  MOAI22 U20883 ( .A1(n28927), .A2(n2041), .B1(ram[7721]), .B2(n2042), 
        .ZN(n11962) );
  MOAI22 U20884 ( .A1(n28692), .A2(n2041), .B1(ram[7722]), .B2(n2042), 
        .ZN(n11963) );
  MOAI22 U20885 ( .A1(n28457), .A2(n2041), .B1(ram[7723]), .B2(n2042), 
        .ZN(n11964) );
  MOAI22 U20886 ( .A1(n28222), .A2(n2041), .B1(ram[7724]), .B2(n2042), 
        .ZN(n11965) );
  MOAI22 U20887 ( .A1(n27987), .A2(n2041), .B1(ram[7725]), .B2(n2042), 
        .ZN(n11966) );
  MOAI22 U20888 ( .A1(n27752), .A2(n2041), .B1(ram[7726]), .B2(n2042), 
        .ZN(n11967) );
  MOAI22 U20889 ( .A1(n27517), .A2(n2041), .B1(ram[7727]), .B2(n2042), 
        .ZN(n11968) );
  MOAI22 U20890 ( .A1(n29162), .A2(n2043), .B1(ram[7728]), .B2(n2044), 
        .ZN(n11969) );
  MOAI22 U20891 ( .A1(n28927), .A2(n2043), .B1(ram[7729]), .B2(n2044), 
        .ZN(n11970) );
  MOAI22 U20892 ( .A1(n28692), .A2(n2043), .B1(ram[7730]), .B2(n2044), 
        .ZN(n11971) );
  MOAI22 U20893 ( .A1(n28457), .A2(n2043), .B1(ram[7731]), .B2(n2044), 
        .ZN(n11972) );
  MOAI22 U20894 ( .A1(n28222), .A2(n2043), .B1(ram[7732]), .B2(n2044), 
        .ZN(n11973) );
  MOAI22 U20895 ( .A1(n27987), .A2(n2043), .B1(ram[7733]), .B2(n2044), 
        .ZN(n11974) );
  MOAI22 U20896 ( .A1(n27752), .A2(n2043), .B1(ram[7734]), .B2(n2044), 
        .ZN(n11975) );
  MOAI22 U20897 ( .A1(n27517), .A2(n2043), .B1(ram[7735]), .B2(n2044), 
        .ZN(n11976) );
  MOAI22 U20898 ( .A1(n29162), .A2(n2045), .B1(ram[7736]), .B2(n2046), 
        .ZN(n11977) );
  MOAI22 U20899 ( .A1(n28927), .A2(n2045), .B1(ram[7737]), .B2(n2046), 
        .ZN(n11978) );
  MOAI22 U20900 ( .A1(n28692), .A2(n2045), .B1(ram[7738]), .B2(n2046), 
        .ZN(n11979) );
  MOAI22 U20901 ( .A1(n28457), .A2(n2045), .B1(ram[7739]), .B2(n2046), 
        .ZN(n11980) );
  MOAI22 U20902 ( .A1(n28222), .A2(n2045), .B1(ram[7740]), .B2(n2046), 
        .ZN(n11981) );
  MOAI22 U20903 ( .A1(n27987), .A2(n2045), .B1(ram[7741]), .B2(n2046), 
        .ZN(n11982) );
  MOAI22 U20904 ( .A1(n27752), .A2(n2045), .B1(ram[7742]), .B2(n2046), 
        .ZN(n11983) );
  MOAI22 U20905 ( .A1(n27517), .A2(n2045), .B1(ram[7743]), .B2(n2046), 
        .ZN(n11984) );
  MOAI22 U20906 ( .A1(n29162), .A2(n2047), .B1(ram[7744]), .B2(n2048), 
        .ZN(n11985) );
  MOAI22 U20907 ( .A1(n28927), .A2(n2047), .B1(ram[7745]), .B2(n2048), 
        .ZN(n11986) );
  MOAI22 U20908 ( .A1(n28692), .A2(n2047), .B1(ram[7746]), .B2(n2048), 
        .ZN(n11987) );
  MOAI22 U20909 ( .A1(n28457), .A2(n2047), .B1(ram[7747]), .B2(n2048), 
        .ZN(n11988) );
  MOAI22 U20910 ( .A1(n28222), .A2(n2047), .B1(ram[7748]), .B2(n2048), 
        .ZN(n11989) );
  MOAI22 U20911 ( .A1(n27987), .A2(n2047), .B1(ram[7749]), .B2(n2048), 
        .ZN(n11990) );
  MOAI22 U20912 ( .A1(n27752), .A2(n2047), .B1(ram[7750]), .B2(n2048), 
        .ZN(n11991) );
  MOAI22 U20913 ( .A1(n27517), .A2(n2047), .B1(ram[7751]), .B2(n2048), 
        .ZN(n11992) );
  MOAI22 U20914 ( .A1(n29162), .A2(n2049), .B1(ram[7752]), .B2(n2050), 
        .ZN(n11993) );
  MOAI22 U20915 ( .A1(n28927), .A2(n2049), .B1(ram[7753]), .B2(n2050), 
        .ZN(n11994) );
  MOAI22 U20916 ( .A1(n28692), .A2(n2049), .B1(ram[7754]), .B2(n2050), 
        .ZN(n11995) );
  MOAI22 U20917 ( .A1(n28457), .A2(n2049), .B1(ram[7755]), .B2(n2050), 
        .ZN(n11996) );
  MOAI22 U20918 ( .A1(n28222), .A2(n2049), .B1(ram[7756]), .B2(n2050), 
        .ZN(n11997) );
  MOAI22 U20919 ( .A1(n27987), .A2(n2049), .B1(ram[7757]), .B2(n2050), 
        .ZN(n11998) );
  MOAI22 U20920 ( .A1(n27752), .A2(n2049), .B1(ram[7758]), .B2(n2050), 
        .ZN(n11999) );
  MOAI22 U20921 ( .A1(n27517), .A2(n2049), .B1(ram[7759]), .B2(n2050), 
        .ZN(n12000) );
  MOAI22 U20922 ( .A1(n29162), .A2(n2051), .B1(ram[7760]), .B2(n2052), 
        .ZN(n12001) );
  MOAI22 U20923 ( .A1(n28927), .A2(n2051), .B1(ram[7761]), .B2(n2052), 
        .ZN(n12002) );
  MOAI22 U20924 ( .A1(n28692), .A2(n2051), .B1(ram[7762]), .B2(n2052), 
        .ZN(n12003) );
  MOAI22 U20925 ( .A1(n28457), .A2(n2051), .B1(ram[7763]), .B2(n2052), 
        .ZN(n12004) );
  MOAI22 U20926 ( .A1(n28222), .A2(n2051), .B1(ram[7764]), .B2(n2052), 
        .ZN(n12005) );
  MOAI22 U20927 ( .A1(n27987), .A2(n2051), .B1(ram[7765]), .B2(n2052), 
        .ZN(n12006) );
  MOAI22 U20928 ( .A1(n27752), .A2(n2051), .B1(ram[7766]), .B2(n2052), 
        .ZN(n12007) );
  MOAI22 U20929 ( .A1(n27517), .A2(n2051), .B1(ram[7767]), .B2(n2052), 
        .ZN(n12008) );
  MOAI22 U20930 ( .A1(n29162), .A2(n2053), .B1(ram[7768]), .B2(n2054), 
        .ZN(n12009) );
  MOAI22 U20931 ( .A1(n28927), .A2(n2053), .B1(ram[7769]), .B2(n2054), 
        .ZN(n12010) );
  MOAI22 U20932 ( .A1(n28692), .A2(n2053), .B1(ram[7770]), .B2(n2054), 
        .ZN(n12011) );
  MOAI22 U20933 ( .A1(n28457), .A2(n2053), .B1(ram[7771]), .B2(n2054), 
        .ZN(n12012) );
  MOAI22 U20934 ( .A1(n28222), .A2(n2053), .B1(ram[7772]), .B2(n2054), 
        .ZN(n12013) );
  MOAI22 U20935 ( .A1(n27987), .A2(n2053), .B1(ram[7773]), .B2(n2054), 
        .ZN(n12014) );
  MOAI22 U20936 ( .A1(n27752), .A2(n2053), .B1(ram[7774]), .B2(n2054), 
        .ZN(n12015) );
  MOAI22 U20937 ( .A1(n27517), .A2(n2053), .B1(ram[7775]), .B2(n2054), 
        .ZN(n12016) );
  MOAI22 U20938 ( .A1(n29162), .A2(n2055), .B1(ram[7776]), .B2(n2056), 
        .ZN(n12017) );
  MOAI22 U20939 ( .A1(n28927), .A2(n2055), .B1(ram[7777]), .B2(n2056), 
        .ZN(n12018) );
  MOAI22 U20940 ( .A1(n28692), .A2(n2055), .B1(ram[7778]), .B2(n2056), 
        .ZN(n12019) );
  MOAI22 U20941 ( .A1(n28457), .A2(n2055), .B1(ram[7779]), .B2(n2056), 
        .ZN(n12020) );
  MOAI22 U20942 ( .A1(n28222), .A2(n2055), .B1(ram[7780]), .B2(n2056), 
        .ZN(n12021) );
  MOAI22 U20943 ( .A1(n27987), .A2(n2055), .B1(ram[7781]), .B2(n2056), 
        .ZN(n12022) );
  MOAI22 U20944 ( .A1(n27752), .A2(n2055), .B1(ram[7782]), .B2(n2056), 
        .ZN(n12023) );
  MOAI22 U20945 ( .A1(n27517), .A2(n2055), .B1(ram[7783]), .B2(n2056), 
        .ZN(n12024) );
  MOAI22 U20946 ( .A1(n29162), .A2(n2057), .B1(ram[7784]), .B2(n2058), 
        .ZN(n12025) );
  MOAI22 U20947 ( .A1(n28927), .A2(n2057), .B1(ram[7785]), .B2(n2058), 
        .ZN(n12026) );
  MOAI22 U20948 ( .A1(n28692), .A2(n2057), .B1(ram[7786]), .B2(n2058), 
        .ZN(n12027) );
  MOAI22 U20949 ( .A1(n28457), .A2(n2057), .B1(ram[7787]), .B2(n2058), 
        .ZN(n12028) );
  MOAI22 U20950 ( .A1(n28222), .A2(n2057), .B1(ram[7788]), .B2(n2058), 
        .ZN(n12029) );
  MOAI22 U20951 ( .A1(n27987), .A2(n2057), .B1(ram[7789]), .B2(n2058), 
        .ZN(n12030) );
  MOAI22 U20952 ( .A1(n27752), .A2(n2057), .B1(ram[7790]), .B2(n2058), 
        .ZN(n12031) );
  MOAI22 U20953 ( .A1(n27517), .A2(n2057), .B1(ram[7791]), .B2(n2058), 
        .ZN(n12032) );
  MOAI22 U20954 ( .A1(n29162), .A2(n2059), .B1(ram[7792]), .B2(n2060), 
        .ZN(n12033) );
  MOAI22 U20955 ( .A1(n28927), .A2(n2059), .B1(ram[7793]), .B2(n2060), 
        .ZN(n12034) );
  MOAI22 U20956 ( .A1(n28692), .A2(n2059), .B1(ram[7794]), .B2(n2060), 
        .ZN(n12035) );
  MOAI22 U20957 ( .A1(n28457), .A2(n2059), .B1(ram[7795]), .B2(n2060), 
        .ZN(n12036) );
  MOAI22 U20958 ( .A1(n28222), .A2(n2059), .B1(ram[7796]), .B2(n2060), 
        .ZN(n12037) );
  MOAI22 U20959 ( .A1(n27987), .A2(n2059), .B1(ram[7797]), .B2(n2060), 
        .ZN(n12038) );
  MOAI22 U20960 ( .A1(n27752), .A2(n2059), .B1(ram[7798]), .B2(n2060), 
        .ZN(n12039) );
  MOAI22 U20961 ( .A1(n27517), .A2(n2059), .B1(ram[7799]), .B2(n2060), 
        .ZN(n12040) );
  MOAI22 U20962 ( .A1(n29163), .A2(n2061), .B1(ram[7800]), .B2(n2062), 
        .ZN(n12041) );
  MOAI22 U20963 ( .A1(n28928), .A2(n2061), .B1(ram[7801]), .B2(n2062), 
        .ZN(n12042) );
  MOAI22 U20964 ( .A1(n28693), .A2(n2061), .B1(ram[7802]), .B2(n2062), 
        .ZN(n12043) );
  MOAI22 U20965 ( .A1(n28458), .A2(n2061), .B1(ram[7803]), .B2(n2062), 
        .ZN(n12044) );
  MOAI22 U20966 ( .A1(n28223), .A2(n2061), .B1(ram[7804]), .B2(n2062), 
        .ZN(n12045) );
  MOAI22 U20967 ( .A1(n27988), .A2(n2061), .B1(ram[7805]), .B2(n2062), 
        .ZN(n12046) );
  MOAI22 U20968 ( .A1(n27753), .A2(n2061), .B1(ram[7806]), .B2(n2062), 
        .ZN(n12047) );
  MOAI22 U20969 ( .A1(n27518), .A2(n2061), .B1(ram[7807]), .B2(n2062), 
        .ZN(n12048) );
  MOAI22 U20970 ( .A1(n29163), .A2(n2063), .B1(ram[7808]), .B2(n2064), 
        .ZN(n12049) );
  MOAI22 U20971 ( .A1(n28928), .A2(n2063), .B1(ram[7809]), .B2(n2064), 
        .ZN(n12050) );
  MOAI22 U20972 ( .A1(n28693), .A2(n2063), .B1(ram[7810]), .B2(n2064), 
        .ZN(n12051) );
  MOAI22 U20973 ( .A1(n28458), .A2(n2063), .B1(ram[7811]), .B2(n2064), 
        .ZN(n12052) );
  MOAI22 U20974 ( .A1(n28223), .A2(n2063), .B1(ram[7812]), .B2(n2064), 
        .ZN(n12053) );
  MOAI22 U20975 ( .A1(n27988), .A2(n2063), .B1(ram[7813]), .B2(n2064), 
        .ZN(n12054) );
  MOAI22 U20976 ( .A1(n27753), .A2(n2063), .B1(ram[7814]), .B2(n2064), 
        .ZN(n12055) );
  MOAI22 U20977 ( .A1(n27518), .A2(n2063), .B1(ram[7815]), .B2(n2064), 
        .ZN(n12056) );
  MOAI22 U20978 ( .A1(n29163), .A2(n2065), .B1(ram[7816]), .B2(n2066), 
        .ZN(n12057) );
  MOAI22 U20979 ( .A1(n28928), .A2(n2065), .B1(ram[7817]), .B2(n2066), 
        .ZN(n12058) );
  MOAI22 U20980 ( .A1(n28693), .A2(n2065), .B1(ram[7818]), .B2(n2066), 
        .ZN(n12059) );
  MOAI22 U20981 ( .A1(n28458), .A2(n2065), .B1(ram[7819]), .B2(n2066), 
        .ZN(n12060) );
  MOAI22 U20982 ( .A1(n28223), .A2(n2065), .B1(ram[7820]), .B2(n2066), 
        .ZN(n12061) );
  MOAI22 U20983 ( .A1(n27988), .A2(n2065), .B1(ram[7821]), .B2(n2066), 
        .ZN(n12062) );
  MOAI22 U20984 ( .A1(n27753), .A2(n2065), .B1(ram[7822]), .B2(n2066), 
        .ZN(n12063) );
  MOAI22 U20985 ( .A1(n27518), .A2(n2065), .B1(ram[7823]), .B2(n2066), 
        .ZN(n12064) );
  MOAI22 U20986 ( .A1(n29163), .A2(n2067), .B1(ram[7824]), .B2(n2068), 
        .ZN(n12065) );
  MOAI22 U20987 ( .A1(n28928), .A2(n2067), .B1(ram[7825]), .B2(n2068), 
        .ZN(n12066) );
  MOAI22 U20988 ( .A1(n28693), .A2(n2067), .B1(ram[7826]), .B2(n2068), 
        .ZN(n12067) );
  MOAI22 U20989 ( .A1(n28458), .A2(n2067), .B1(ram[7827]), .B2(n2068), 
        .ZN(n12068) );
  MOAI22 U20990 ( .A1(n28223), .A2(n2067), .B1(ram[7828]), .B2(n2068), 
        .ZN(n12069) );
  MOAI22 U20991 ( .A1(n27988), .A2(n2067), .B1(ram[7829]), .B2(n2068), 
        .ZN(n12070) );
  MOAI22 U20992 ( .A1(n27753), .A2(n2067), .B1(ram[7830]), .B2(n2068), 
        .ZN(n12071) );
  MOAI22 U20993 ( .A1(n27518), .A2(n2067), .B1(ram[7831]), .B2(n2068), 
        .ZN(n12072) );
  MOAI22 U20994 ( .A1(n29163), .A2(n2069), .B1(ram[7832]), .B2(n2070), 
        .ZN(n12073) );
  MOAI22 U20995 ( .A1(n28928), .A2(n2069), .B1(ram[7833]), .B2(n2070), 
        .ZN(n12074) );
  MOAI22 U20996 ( .A1(n28693), .A2(n2069), .B1(ram[7834]), .B2(n2070), 
        .ZN(n12075) );
  MOAI22 U20997 ( .A1(n28458), .A2(n2069), .B1(ram[7835]), .B2(n2070), 
        .ZN(n12076) );
  MOAI22 U20998 ( .A1(n28223), .A2(n2069), .B1(ram[7836]), .B2(n2070), 
        .ZN(n12077) );
  MOAI22 U20999 ( .A1(n27988), .A2(n2069), .B1(ram[7837]), .B2(n2070), 
        .ZN(n12078) );
  MOAI22 U21000 ( .A1(n27753), .A2(n2069), .B1(ram[7838]), .B2(n2070), 
        .ZN(n12079) );
  MOAI22 U21001 ( .A1(n27518), .A2(n2069), .B1(ram[7839]), .B2(n2070), 
        .ZN(n12080) );
  MOAI22 U21002 ( .A1(n29163), .A2(n2071), .B1(ram[7840]), .B2(n2072), 
        .ZN(n12081) );
  MOAI22 U21003 ( .A1(n28928), .A2(n2071), .B1(ram[7841]), .B2(n2072), 
        .ZN(n12082) );
  MOAI22 U21004 ( .A1(n28693), .A2(n2071), .B1(ram[7842]), .B2(n2072), 
        .ZN(n12083) );
  MOAI22 U21005 ( .A1(n28458), .A2(n2071), .B1(ram[7843]), .B2(n2072), 
        .ZN(n12084) );
  MOAI22 U21006 ( .A1(n28223), .A2(n2071), .B1(ram[7844]), .B2(n2072), 
        .ZN(n12085) );
  MOAI22 U21007 ( .A1(n27988), .A2(n2071), .B1(ram[7845]), .B2(n2072), 
        .ZN(n12086) );
  MOAI22 U21008 ( .A1(n27753), .A2(n2071), .B1(ram[7846]), .B2(n2072), 
        .ZN(n12087) );
  MOAI22 U21009 ( .A1(n27518), .A2(n2071), .B1(ram[7847]), .B2(n2072), 
        .ZN(n12088) );
  MOAI22 U21010 ( .A1(n29163), .A2(n2073), .B1(ram[7848]), .B2(n2074), 
        .ZN(n12089) );
  MOAI22 U21011 ( .A1(n28928), .A2(n2073), .B1(ram[7849]), .B2(n2074), 
        .ZN(n12090) );
  MOAI22 U21012 ( .A1(n28693), .A2(n2073), .B1(ram[7850]), .B2(n2074), 
        .ZN(n12091) );
  MOAI22 U21013 ( .A1(n28458), .A2(n2073), .B1(ram[7851]), .B2(n2074), 
        .ZN(n12092) );
  MOAI22 U21014 ( .A1(n28223), .A2(n2073), .B1(ram[7852]), .B2(n2074), 
        .ZN(n12093) );
  MOAI22 U21015 ( .A1(n27988), .A2(n2073), .B1(ram[7853]), .B2(n2074), 
        .ZN(n12094) );
  MOAI22 U21016 ( .A1(n27753), .A2(n2073), .B1(ram[7854]), .B2(n2074), 
        .ZN(n12095) );
  MOAI22 U21017 ( .A1(n27518), .A2(n2073), .B1(ram[7855]), .B2(n2074), 
        .ZN(n12096) );
  MOAI22 U21018 ( .A1(n29163), .A2(n2075), .B1(ram[7856]), .B2(n2076), 
        .ZN(n12097) );
  MOAI22 U21019 ( .A1(n28928), .A2(n2075), .B1(ram[7857]), .B2(n2076), 
        .ZN(n12098) );
  MOAI22 U21020 ( .A1(n28693), .A2(n2075), .B1(ram[7858]), .B2(n2076), 
        .ZN(n12099) );
  MOAI22 U21021 ( .A1(n28458), .A2(n2075), .B1(ram[7859]), .B2(n2076), 
        .ZN(n12100) );
  MOAI22 U21022 ( .A1(n28223), .A2(n2075), .B1(ram[7860]), .B2(n2076), 
        .ZN(n12101) );
  MOAI22 U21023 ( .A1(n27988), .A2(n2075), .B1(ram[7861]), .B2(n2076), 
        .ZN(n12102) );
  MOAI22 U21024 ( .A1(n27753), .A2(n2075), .B1(ram[7862]), .B2(n2076), 
        .ZN(n12103) );
  MOAI22 U21025 ( .A1(n27518), .A2(n2075), .B1(ram[7863]), .B2(n2076), 
        .ZN(n12104) );
  MOAI22 U21026 ( .A1(n29163), .A2(n2077), .B1(ram[7864]), .B2(n2078), 
        .ZN(n12105) );
  MOAI22 U21027 ( .A1(n28928), .A2(n2077), .B1(ram[7865]), .B2(n2078), 
        .ZN(n12106) );
  MOAI22 U21028 ( .A1(n28693), .A2(n2077), .B1(ram[7866]), .B2(n2078), 
        .ZN(n12107) );
  MOAI22 U21029 ( .A1(n28458), .A2(n2077), .B1(ram[7867]), .B2(n2078), 
        .ZN(n12108) );
  MOAI22 U21030 ( .A1(n28223), .A2(n2077), .B1(ram[7868]), .B2(n2078), 
        .ZN(n12109) );
  MOAI22 U21031 ( .A1(n27988), .A2(n2077), .B1(ram[7869]), .B2(n2078), 
        .ZN(n12110) );
  MOAI22 U21032 ( .A1(n27753), .A2(n2077), .B1(ram[7870]), .B2(n2078), 
        .ZN(n12111) );
  MOAI22 U21033 ( .A1(n27518), .A2(n2077), .B1(ram[7871]), .B2(n2078), 
        .ZN(n12112) );
  MOAI22 U21034 ( .A1(n29163), .A2(n2079), .B1(ram[7872]), .B2(n2080), 
        .ZN(n12113) );
  MOAI22 U21035 ( .A1(n28928), .A2(n2079), .B1(ram[7873]), .B2(n2080), 
        .ZN(n12114) );
  MOAI22 U21036 ( .A1(n28693), .A2(n2079), .B1(ram[7874]), .B2(n2080), 
        .ZN(n12115) );
  MOAI22 U21037 ( .A1(n28458), .A2(n2079), .B1(ram[7875]), .B2(n2080), 
        .ZN(n12116) );
  MOAI22 U21038 ( .A1(n28223), .A2(n2079), .B1(ram[7876]), .B2(n2080), 
        .ZN(n12117) );
  MOAI22 U21039 ( .A1(n27988), .A2(n2079), .B1(ram[7877]), .B2(n2080), 
        .ZN(n12118) );
  MOAI22 U21040 ( .A1(n27753), .A2(n2079), .B1(ram[7878]), .B2(n2080), 
        .ZN(n12119) );
  MOAI22 U21041 ( .A1(n27518), .A2(n2079), .B1(ram[7879]), .B2(n2080), 
        .ZN(n12120) );
  MOAI22 U21042 ( .A1(n29163), .A2(n2081), .B1(ram[7880]), .B2(n2082), 
        .ZN(n12121) );
  MOAI22 U21043 ( .A1(n28928), .A2(n2081), .B1(ram[7881]), .B2(n2082), 
        .ZN(n12122) );
  MOAI22 U21044 ( .A1(n28693), .A2(n2081), .B1(ram[7882]), .B2(n2082), 
        .ZN(n12123) );
  MOAI22 U21045 ( .A1(n28458), .A2(n2081), .B1(ram[7883]), .B2(n2082), 
        .ZN(n12124) );
  MOAI22 U21046 ( .A1(n28223), .A2(n2081), .B1(ram[7884]), .B2(n2082), 
        .ZN(n12125) );
  MOAI22 U21047 ( .A1(n27988), .A2(n2081), .B1(ram[7885]), .B2(n2082), 
        .ZN(n12126) );
  MOAI22 U21048 ( .A1(n27753), .A2(n2081), .B1(ram[7886]), .B2(n2082), 
        .ZN(n12127) );
  MOAI22 U21049 ( .A1(n27518), .A2(n2081), .B1(ram[7887]), .B2(n2082), 
        .ZN(n12128) );
  MOAI22 U21050 ( .A1(n29163), .A2(n2083), .B1(ram[7888]), .B2(n2084), 
        .ZN(n12129) );
  MOAI22 U21051 ( .A1(n28928), .A2(n2083), .B1(ram[7889]), .B2(n2084), 
        .ZN(n12130) );
  MOAI22 U21052 ( .A1(n28693), .A2(n2083), .B1(ram[7890]), .B2(n2084), 
        .ZN(n12131) );
  MOAI22 U21053 ( .A1(n28458), .A2(n2083), .B1(ram[7891]), .B2(n2084), 
        .ZN(n12132) );
  MOAI22 U21054 ( .A1(n28223), .A2(n2083), .B1(ram[7892]), .B2(n2084), 
        .ZN(n12133) );
  MOAI22 U21055 ( .A1(n27988), .A2(n2083), .B1(ram[7893]), .B2(n2084), 
        .ZN(n12134) );
  MOAI22 U21056 ( .A1(n27753), .A2(n2083), .B1(ram[7894]), .B2(n2084), 
        .ZN(n12135) );
  MOAI22 U21057 ( .A1(n27518), .A2(n2083), .B1(ram[7895]), .B2(n2084), 
        .ZN(n12136) );
  MOAI22 U21058 ( .A1(n29163), .A2(n2085), .B1(ram[7896]), .B2(n2086), 
        .ZN(n12137) );
  MOAI22 U21059 ( .A1(n28928), .A2(n2085), .B1(ram[7897]), .B2(n2086), 
        .ZN(n12138) );
  MOAI22 U21060 ( .A1(n28693), .A2(n2085), .B1(ram[7898]), .B2(n2086), 
        .ZN(n12139) );
  MOAI22 U21061 ( .A1(n28458), .A2(n2085), .B1(ram[7899]), .B2(n2086), 
        .ZN(n12140) );
  MOAI22 U21062 ( .A1(n28223), .A2(n2085), .B1(ram[7900]), .B2(n2086), 
        .ZN(n12141) );
  MOAI22 U21063 ( .A1(n27988), .A2(n2085), .B1(ram[7901]), .B2(n2086), 
        .ZN(n12142) );
  MOAI22 U21064 ( .A1(n27753), .A2(n2085), .B1(ram[7902]), .B2(n2086), 
        .ZN(n12143) );
  MOAI22 U21065 ( .A1(n27518), .A2(n2085), .B1(ram[7903]), .B2(n2086), 
        .ZN(n12144) );
  MOAI22 U21066 ( .A1(n29164), .A2(n2087), .B1(ram[7904]), .B2(n2088), 
        .ZN(n12145) );
  MOAI22 U21067 ( .A1(n28929), .A2(n2087), .B1(ram[7905]), .B2(n2088), 
        .ZN(n12146) );
  MOAI22 U21068 ( .A1(n28694), .A2(n2087), .B1(ram[7906]), .B2(n2088), 
        .ZN(n12147) );
  MOAI22 U21069 ( .A1(n28459), .A2(n2087), .B1(ram[7907]), .B2(n2088), 
        .ZN(n12148) );
  MOAI22 U21070 ( .A1(n28224), .A2(n2087), .B1(ram[7908]), .B2(n2088), 
        .ZN(n12149) );
  MOAI22 U21071 ( .A1(n27989), .A2(n2087), .B1(ram[7909]), .B2(n2088), 
        .ZN(n12150) );
  MOAI22 U21072 ( .A1(n27754), .A2(n2087), .B1(ram[7910]), .B2(n2088), 
        .ZN(n12151) );
  MOAI22 U21073 ( .A1(n27519), .A2(n2087), .B1(ram[7911]), .B2(n2088), 
        .ZN(n12152) );
  MOAI22 U21074 ( .A1(n29164), .A2(n2089), .B1(ram[7912]), .B2(n2090), 
        .ZN(n12153) );
  MOAI22 U21075 ( .A1(n28929), .A2(n2089), .B1(ram[7913]), .B2(n2090), 
        .ZN(n12154) );
  MOAI22 U21076 ( .A1(n28694), .A2(n2089), .B1(ram[7914]), .B2(n2090), 
        .ZN(n12155) );
  MOAI22 U21077 ( .A1(n28459), .A2(n2089), .B1(ram[7915]), .B2(n2090), 
        .ZN(n12156) );
  MOAI22 U21078 ( .A1(n28224), .A2(n2089), .B1(ram[7916]), .B2(n2090), 
        .ZN(n12157) );
  MOAI22 U21079 ( .A1(n27989), .A2(n2089), .B1(ram[7917]), .B2(n2090), 
        .ZN(n12158) );
  MOAI22 U21080 ( .A1(n27754), .A2(n2089), .B1(ram[7918]), .B2(n2090), 
        .ZN(n12159) );
  MOAI22 U21081 ( .A1(n27519), .A2(n2089), .B1(ram[7919]), .B2(n2090), 
        .ZN(n12160) );
  MOAI22 U21082 ( .A1(n29164), .A2(n2091), .B1(ram[7920]), .B2(n2092), 
        .ZN(n12161) );
  MOAI22 U21083 ( .A1(n28929), .A2(n2091), .B1(ram[7921]), .B2(n2092), 
        .ZN(n12162) );
  MOAI22 U21084 ( .A1(n28694), .A2(n2091), .B1(ram[7922]), .B2(n2092), 
        .ZN(n12163) );
  MOAI22 U21085 ( .A1(n28459), .A2(n2091), .B1(ram[7923]), .B2(n2092), 
        .ZN(n12164) );
  MOAI22 U21086 ( .A1(n28224), .A2(n2091), .B1(ram[7924]), .B2(n2092), 
        .ZN(n12165) );
  MOAI22 U21087 ( .A1(n27989), .A2(n2091), .B1(ram[7925]), .B2(n2092), 
        .ZN(n12166) );
  MOAI22 U21088 ( .A1(n27754), .A2(n2091), .B1(ram[7926]), .B2(n2092), 
        .ZN(n12167) );
  MOAI22 U21089 ( .A1(n27519), .A2(n2091), .B1(ram[7927]), .B2(n2092), 
        .ZN(n12168) );
  MOAI22 U21090 ( .A1(n29164), .A2(n2093), .B1(ram[7928]), .B2(n2094), 
        .ZN(n12169) );
  MOAI22 U21091 ( .A1(n28929), .A2(n2093), .B1(ram[7929]), .B2(n2094), 
        .ZN(n12170) );
  MOAI22 U21092 ( .A1(n28694), .A2(n2093), .B1(ram[7930]), .B2(n2094), 
        .ZN(n12171) );
  MOAI22 U21093 ( .A1(n28459), .A2(n2093), .B1(ram[7931]), .B2(n2094), 
        .ZN(n12172) );
  MOAI22 U21094 ( .A1(n28224), .A2(n2093), .B1(ram[7932]), .B2(n2094), 
        .ZN(n12173) );
  MOAI22 U21095 ( .A1(n27989), .A2(n2093), .B1(ram[7933]), .B2(n2094), 
        .ZN(n12174) );
  MOAI22 U21096 ( .A1(n27754), .A2(n2093), .B1(ram[7934]), .B2(n2094), 
        .ZN(n12175) );
  MOAI22 U21097 ( .A1(n27519), .A2(n2093), .B1(ram[7935]), .B2(n2094), 
        .ZN(n12176) );
  MOAI22 U21098 ( .A1(n29164), .A2(n2095), .B1(ram[7936]), .B2(n2096), 
        .ZN(n12177) );
  MOAI22 U21099 ( .A1(n28929), .A2(n2095), .B1(ram[7937]), .B2(n2096), 
        .ZN(n12178) );
  MOAI22 U21100 ( .A1(n28694), .A2(n2095), .B1(ram[7938]), .B2(n2096), 
        .ZN(n12179) );
  MOAI22 U21101 ( .A1(n28459), .A2(n2095), .B1(ram[7939]), .B2(n2096), 
        .ZN(n12180) );
  MOAI22 U21102 ( .A1(n28224), .A2(n2095), .B1(ram[7940]), .B2(n2096), 
        .ZN(n12181) );
  MOAI22 U21103 ( .A1(n27989), .A2(n2095), .B1(ram[7941]), .B2(n2096), 
        .ZN(n12182) );
  MOAI22 U21104 ( .A1(n27754), .A2(n2095), .B1(ram[7942]), .B2(n2096), 
        .ZN(n12183) );
  MOAI22 U21105 ( .A1(n27519), .A2(n2095), .B1(ram[7943]), .B2(n2096), 
        .ZN(n12184) );
  MOAI22 U21106 ( .A1(n29164), .A2(n2097), .B1(ram[7944]), .B2(n2098), 
        .ZN(n12185) );
  MOAI22 U21107 ( .A1(n28929), .A2(n2097), .B1(ram[7945]), .B2(n2098), 
        .ZN(n12186) );
  MOAI22 U21108 ( .A1(n28694), .A2(n2097), .B1(ram[7946]), .B2(n2098), 
        .ZN(n12187) );
  MOAI22 U21109 ( .A1(n28459), .A2(n2097), .B1(ram[7947]), .B2(n2098), 
        .ZN(n12188) );
  MOAI22 U21110 ( .A1(n28224), .A2(n2097), .B1(ram[7948]), .B2(n2098), 
        .ZN(n12189) );
  MOAI22 U21111 ( .A1(n27989), .A2(n2097), .B1(ram[7949]), .B2(n2098), 
        .ZN(n12190) );
  MOAI22 U21112 ( .A1(n27754), .A2(n2097), .B1(ram[7950]), .B2(n2098), 
        .ZN(n12191) );
  MOAI22 U21113 ( .A1(n27519), .A2(n2097), .B1(ram[7951]), .B2(n2098), 
        .ZN(n12192) );
  MOAI22 U21114 ( .A1(n29164), .A2(n2099), .B1(ram[7952]), .B2(n2100), 
        .ZN(n12193) );
  MOAI22 U21115 ( .A1(n28929), .A2(n2099), .B1(ram[7953]), .B2(n2100), 
        .ZN(n12194) );
  MOAI22 U21116 ( .A1(n28694), .A2(n2099), .B1(ram[7954]), .B2(n2100), 
        .ZN(n12195) );
  MOAI22 U21117 ( .A1(n28459), .A2(n2099), .B1(ram[7955]), .B2(n2100), 
        .ZN(n12196) );
  MOAI22 U21118 ( .A1(n28224), .A2(n2099), .B1(ram[7956]), .B2(n2100), 
        .ZN(n12197) );
  MOAI22 U21119 ( .A1(n27989), .A2(n2099), .B1(ram[7957]), .B2(n2100), 
        .ZN(n12198) );
  MOAI22 U21120 ( .A1(n27754), .A2(n2099), .B1(ram[7958]), .B2(n2100), 
        .ZN(n12199) );
  MOAI22 U21121 ( .A1(n27519), .A2(n2099), .B1(ram[7959]), .B2(n2100), 
        .ZN(n12200) );
  MOAI22 U21122 ( .A1(n29164), .A2(n2101), .B1(ram[7960]), .B2(n2102), 
        .ZN(n12201) );
  MOAI22 U21123 ( .A1(n28929), .A2(n2101), .B1(ram[7961]), .B2(n2102), 
        .ZN(n12202) );
  MOAI22 U21124 ( .A1(n28694), .A2(n2101), .B1(ram[7962]), .B2(n2102), 
        .ZN(n12203) );
  MOAI22 U21125 ( .A1(n28459), .A2(n2101), .B1(ram[7963]), .B2(n2102), 
        .ZN(n12204) );
  MOAI22 U21126 ( .A1(n28224), .A2(n2101), .B1(ram[7964]), .B2(n2102), 
        .ZN(n12205) );
  MOAI22 U21127 ( .A1(n27989), .A2(n2101), .B1(ram[7965]), .B2(n2102), 
        .ZN(n12206) );
  MOAI22 U21128 ( .A1(n27754), .A2(n2101), .B1(ram[7966]), .B2(n2102), 
        .ZN(n12207) );
  MOAI22 U21129 ( .A1(n27519), .A2(n2101), .B1(ram[7967]), .B2(n2102), 
        .ZN(n12208) );
  MOAI22 U21130 ( .A1(n29164), .A2(n2103), .B1(ram[7968]), .B2(n2104), 
        .ZN(n12209) );
  MOAI22 U21131 ( .A1(n28929), .A2(n2103), .B1(ram[7969]), .B2(n2104), 
        .ZN(n12210) );
  MOAI22 U21132 ( .A1(n28694), .A2(n2103), .B1(ram[7970]), .B2(n2104), 
        .ZN(n12211) );
  MOAI22 U21133 ( .A1(n28459), .A2(n2103), .B1(ram[7971]), .B2(n2104), 
        .ZN(n12212) );
  MOAI22 U21134 ( .A1(n28224), .A2(n2103), .B1(ram[7972]), .B2(n2104), 
        .ZN(n12213) );
  MOAI22 U21135 ( .A1(n27989), .A2(n2103), .B1(ram[7973]), .B2(n2104), 
        .ZN(n12214) );
  MOAI22 U21136 ( .A1(n27754), .A2(n2103), .B1(ram[7974]), .B2(n2104), 
        .ZN(n12215) );
  MOAI22 U21137 ( .A1(n27519), .A2(n2103), .B1(ram[7975]), .B2(n2104), 
        .ZN(n12216) );
  MOAI22 U21138 ( .A1(n29164), .A2(n2105), .B1(ram[7976]), .B2(n2106), 
        .ZN(n12217) );
  MOAI22 U21139 ( .A1(n28929), .A2(n2105), .B1(ram[7977]), .B2(n2106), 
        .ZN(n12218) );
  MOAI22 U21140 ( .A1(n28694), .A2(n2105), .B1(ram[7978]), .B2(n2106), 
        .ZN(n12219) );
  MOAI22 U21141 ( .A1(n28459), .A2(n2105), .B1(ram[7979]), .B2(n2106), 
        .ZN(n12220) );
  MOAI22 U21142 ( .A1(n28224), .A2(n2105), .B1(ram[7980]), .B2(n2106), 
        .ZN(n12221) );
  MOAI22 U21143 ( .A1(n27989), .A2(n2105), .B1(ram[7981]), .B2(n2106), 
        .ZN(n12222) );
  MOAI22 U21144 ( .A1(n27754), .A2(n2105), .B1(ram[7982]), .B2(n2106), 
        .ZN(n12223) );
  MOAI22 U21145 ( .A1(n27519), .A2(n2105), .B1(ram[7983]), .B2(n2106), 
        .ZN(n12224) );
  MOAI22 U21146 ( .A1(n29164), .A2(n2107), .B1(ram[7984]), .B2(n2108), 
        .ZN(n12225) );
  MOAI22 U21147 ( .A1(n28929), .A2(n2107), .B1(ram[7985]), .B2(n2108), 
        .ZN(n12226) );
  MOAI22 U21148 ( .A1(n28694), .A2(n2107), .B1(ram[7986]), .B2(n2108), 
        .ZN(n12227) );
  MOAI22 U21149 ( .A1(n28459), .A2(n2107), .B1(ram[7987]), .B2(n2108), 
        .ZN(n12228) );
  MOAI22 U21150 ( .A1(n28224), .A2(n2107), .B1(ram[7988]), .B2(n2108), 
        .ZN(n12229) );
  MOAI22 U21151 ( .A1(n27989), .A2(n2107), .B1(ram[7989]), .B2(n2108), 
        .ZN(n12230) );
  MOAI22 U21152 ( .A1(n27754), .A2(n2107), .B1(ram[7990]), .B2(n2108), 
        .ZN(n12231) );
  MOAI22 U21153 ( .A1(n27519), .A2(n2107), .B1(ram[7991]), .B2(n2108), 
        .ZN(n12232) );
  MOAI22 U21154 ( .A1(n29164), .A2(n2109), .B1(ram[7992]), .B2(n2110), 
        .ZN(n12233) );
  MOAI22 U21155 ( .A1(n28929), .A2(n2109), .B1(ram[7993]), .B2(n2110), 
        .ZN(n12234) );
  MOAI22 U21156 ( .A1(n28694), .A2(n2109), .B1(ram[7994]), .B2(n2110), 
        .ZN(n12235) );
  MOAI22 U21157 ( .A1(n28459), .A2(n2109), .B1(ram[7995]), .B2(n2110), 
        .ZN(n12236) );
  MOAI22 U21158 ( .A1(n28224), .A2(n2109), .B1(ram[7996]), .B2(n2110), 
        .ZN(n12237) );
  MOAI22 U21159 ( .A1(n27989), .A2(n2109), .B1(ram[7997]), .B2(n2110), 
        .ZN(n12238) );
  MOAI22 U21160 ( .A1(n27754), .A2(n2109), .B1(ram[7998]), .B2(n2110), 
        .ZN(n12239) );
  MOAI22 U21161 ( .A1(n27519), .A2(n2109), .B1(ram[7999]), .B2(n2110), 
        .ZN(n12240) );
  MOAI22 U21162 ( .A1(n29164), .A2(n2111), .B1(ram[8000]), .B2(n2112), 
        .ZN(n12241) );
  MOAI22 U21163 ( .A1(n28929), .A2(n2111), .B1(ram[8001]), .B2(n2112), 
        .ZN(n12242) );
  MOAI22 U21164 ( .A1(n28694), .A2(n2111), .B1(ram[8002]), .B2(n2112), 
        .ZN(n12243) );
  MOAI22 U21165 ( .A1(n28459), .A2(n2111), .B1(ram[8003]), .B2(n2112), 
        .ZN(n12244) );
  MOAI22 U21166 ( .A1(n28224), .A2(n2111), .B1(ram[8004]), .B2(n2112), 
        .ZN(n12245) );
  MOAI22 U21167 ( .A1(n27989), .A2(n2111), .B1(ram[8005]), .B2(n2112), 
        .ZN(n12246) );
  MOAI22 U21168 ( .A1(n27754), .A2(n2111), .B1(ram[8006]), .B2(n2112), 
        .ZN(n12247) );
  MOAI22 U21169 ( .A1(n27519), .A2(n2111), .B1(ram[8007]), .B2(n2112), 
        .ZN(n12248) );
  MOAI22 U21170 ( .A1(n29165), .A2(n2113), .B1(ram[8008]), .B2(n2114), 
        .ZN(n12249) );
  MOAI22 U21171 ( .A1(n28930), .A2(n2113), .B1(ram[8009]), .B2(n2114), 
        .ZN(n12250) );
  MOAI22 U21172 ( .A1(n28695), .A2(n2113), .B1(ram[8010]), .B2(n2114), 
        .ZN(n12251) );
  MOAI22 U21173 ( .A1(n28460), .A2(n2113), .B1(ram[8011]), .B2(n2114), 
        .ZN(n12252) );
  MOAI22 U21174 ( .A1(n28225), .A2(n2113), .B1(ram[8012]), .B2(n2114), 
        .ZN(n12253) );
  MOAI22 U21175 ( .A1(n27990), .A2(n2113), .B1(ram[8013]), .B2(n2114), 
        .ZN(n12254) );
  MOAI22 U21176 ( .A1(n27755), .A2(n2113), .B1(ram[8014]), .B2(n2114), 
        .ZN(n12255) );
  MOAI22 U21177 ( .A1(n27520), .A2(n2113), .B1(ram[8015]), .B2(n2114), 
        .ZN(n12256) );
  MOAI22 U21178 ( .A1(n29165), .A2(n2115), .B1(ram[8016]), .B2(n2116), 
        .ZN(n12257) );
  MOAI22 U21179 ( .A1(n28930), .A2(n2115), .B1(ram[8017]), .B2(n2116), 
        .ZN(n12258) );
  MOAI22 U21180 ( .A1(n28695), .A2(n2115), .B1(ram[8018]), .B2(n2116), 
        .ZN(n12259) );
  MOAI22 U21181 ( .A1(n28460), .A2(n2115), .B1(ram[8019]), .B2(n2116), 
        .ZN(n12260) );
  MOAI22 U21182 ( .A1(n28225), .A2(n2115), .B1(ram[8020]), .B2(n2116), 
        .ZN(n12261) );
  MOAI22 U21183 ( .A1(n27990), .A2(n2115), .B1(ram[8021]), .B2(n2116), 
        .ZN(n12262) );
  MOAI22 U21184 ( .A1(n27755), .A2(n2115), .B1(ram[8022]), .B2(n2116), 
        .ZN(n12263) );
  MOAI22 U21185 ( .A1(n27520), .A2(n2115), .B1(ram[8023]), .B2(n2116), 
        .ZN(n12264) );
  MOAI22 U21186 ( .A1(n29165), .A2(n2117), .B1(ram[8024]), .B2(n2118), 
        .ZN(n12265) );
  MOAI22 U21187 ( .A1(n28930), .A2(n2117), .B1(ram[8025]), .B2(n2118), 
        .ZN(n12266) );
  MOAI22 U21188 ( .A1(n28695), .A2(n2117), .B1(ram[8026]), .B2(n2118), 
        .ZN(n12267) );
  MOAI22 U21189 ( .A1(n28460), .A2(n2117), .B1(ram[8027]), .B2(n2118), 
        .ZN(n12268) );
  MOAI22 U21190 ( .A1(n28225), .A2(n2117), .B1(ram[8028]), .B2(n2118), 
        .ZN(n12269) );
  MOAI22 U21191 ( .A1(n27990), .A2(n2117), .B1(ram[8029]), .B2(n2118), 
        .ZN(n12270) );
  MOAI22 U21192 ( .A1(n27755), .A2(n2117), .B1(ram[8030]), .B2(n2118), 
        .ZN(n12271) );
  MOAI22 U21193 ( .A1(n27520), .A2(n2117), .B1(ram[8031]), .B2(n2118), 
        .ZN(n12272) );
  MOAI22 U21194 ( .A1(n29165), .A2(n2119), .B1(ram[8032]), .B2(n2120), 
        .ZN(n12273) );
  MOAI22 U21195 ( .A1(n28930), .A2(n2119), .B1(ram[8033]), .B2(n2120), 
        .ZN(n12274) );
  MOAI22 U21196 ( .A1(n28695), .A2(n2119), .B1(ram[8034]), .B2(n2120), 
        .ZN(n12275) );
  MOAI22 U21197 ( .A1(n28460), .A2(n2119), .B1(ram[8035]), .B2(n2120), 
        .ZN(n12276) );
  MOAI22 U21198 ( .A1(n28225), .A2(n2119), .B1(ram[8036]), .B2(n2120), 
        .ZN(n12277) );
  MOAI22 U21199 ( .A1(n27990), .A2(n2119), .B1(ram[8037]), .B2(n2120), 
        .ZN(n12278) );
  MOAI22 U21200 ( .A1(n27755), .A2(n2119), .B1(ram[8038]), .B2(n2120), 
        .ZN(n12279) );
  MOAI22 U21201 ( .A1(n27520), .A2(n2119), .B1(ram[8039]), .B2(n2120), 
        .ZN(n12280) );
  MOAI22 U21202 ( .A1(n29165), .A2(n2121), .B1(ram[8040]), .B2(n2122), 
        .ZN(n12281) );
  MOAI22 U21203 ( .A1(n28930), .A2(n2121), .B1(ram[8041]), .B2(n2122), 
        .ZN(n12282) );
  MOAI22 U21204 ( .A1(n28695), .A2(n2121), .B1(ram[8042]), .B2(n2122), 
        .ZN(n12283) );
  MOAI22 U21205 ( .A1(n28460), .A2(n2121), .B1(ram[8043]), .B2(n2122), 
        .ZN(n12284) );
  MOAI22 U21206 ( .A1(n28225), .A2(n2121), .B1(ram[8044]), .B2(n2122), 
        .ZN(n12285) );
  MOAI22 U21207 ( .A1(n27990), .A2(n2121), .B1(ram[8045]), .B2(n2122), 
        .ZN(n12286) );
  MOAI22 U21208 ( .A1(n27755), .A2(n2121), .B1(ram[8046]), .B2(n2122), 
        .ZN(n12287) );
  MOAI22 U21209 ( .A1(n27520), .A2(n2121), .B1(ram[8047]), .B2(n2122), 
        .ZN(n12288) );
  MOAI22 U21210 ( .A1(n29165), .A2(n2123), .B1(ram[8048]), .B2(n2124), 
        .ZN(n12289) );
  MOAI22 U21211 ( .A1(n28930), .A2(n2123), .B1(ram[8049]), .B2(n2124), 
        .ZN(n12290) );
  MOAI22 U21212 ( .A1(n28695), .A2(n2123), .B1(ram[8050]), .B2(n2124), 
        .ZN(n12291) );
  MOAI22 U21213 ( .A1(n28460), .A2(n2123), .B1(ram[8051]), .B2(n2124), 
        .ZN(n12292) );
  MOAI22 U21214 ( .A1(n28225), .A2(n2123), .B1(ram[8052]), .B2(n2124), 
        .ZN(n12293) );
  MOAI22 U21215 ( .A1(n27990), .A2(n2123), .B1(ram[8053]), .B2(n2124), 
        .ZN(n12294) );
  MOAI22 U21216 ( .A1(n27755), .A2(n2123), .B1(ram[8054]), .B2(n2124), 
        .ZN(n12295) );
  MOAI22 U21217 ( .A1(n27520), .A2(n2123), .B1(ram[8055]), .B2(n2124), 
        .ZN(n12296) );
  MOAI22 U21218 ( .A1(n29165), .A2(n2125), .B1(ram[8056]), .B2(n2126), 
        .ZN(n12297) );
  MOAI22 U21219 ( .A1(n28930), .A2(n2125), .B1(ram[8057]), .B2(n2126), 
        .ZN(n12298) );
  MOAI22 U21220 ( .A1(n28695), .A2(n2125), .B1(ram[8058]), .B2(n2126), 
        .ZN(n12299) );
  MOAI22 U21221 ( .A1(n28460), .A2(n2125), .B1(ram[8059]), .B2(n2126), 
        .ZN(n12300) );
  MOAI22 U21222 ( .A1(n28225), .A2(n2125), .B1(ram[8060]), .B2(n2126), 
        .ZN(n12301) );
  MOAI22 U21223 ( .A1(n27990), .A2(n2125), .B1(ram[8061]), .B2(n2126), 
        .ZN(n12302) );
  MOAI22 U21224 ( .A1(n27755), .A2(n2125), .B1(ram[8062]), .B2(n2126), 
        .ZN(n12303) );
  MOAI22 U21225 ( .A1(n27520), .A2(n2125), .B1(ram[8063]), .B2(n2126), 
        .ZN(n12304) );
  MOAI22 U21226 ( .A1(n29165), .A2(n2127), .B1(ram[8064]), .B2(n2128), 
        .ZN(n12305) );
  MOAI22 U21227 ( .A1(n28930), .A2(n2127), .B1(ram[8065]), .B2(n2128), 
        .ZN(n12306) );
  MOAI22 U21228 ( .A1(n28695), .A2(n2127), .B1(ram[8066]), .B2(n2128), 
        .ZN(n12307) );
  MOAI22 U21229 ( .A1(n28460), .A2(n2127), .B1(ram[8067]), .B2(n2128), 
        .ZN(n12308) );
  MOAI22 U21230 ( .A1(n28225), .A2(n2127), .B1(ram[8068]), .B2(n2128), 
        .ZN(n12309) );
  MOAI22 U21231 ( .A1(n27990), .A2(n2127), .B1(ram[8069]), .B2(n2128), 
        .ZN(n12310) );
  MOAI22 U21232 ( .A1(n27755), .A2(n2127), .B1(ram[8070]), .B2(n2128), 
        .ZN(n12311) );
  MOAI22 U21233 ( .A1(n27520), .A2(n2127), .B1(ram[8071]), .B2(n2128), 
        .ZN(n12312) );
  MOAI22 U21234 ( .A1(n29165), .A2(n2129), .B1(ram[8072]), .B2(n2130), 
        .ZN(n12313) );
  MOAI22 U21235 ( .A1(n28930), .A2(n2129), .B1(ram[8073]), .B2(n2130), 
        .ZN(n12314) );
  MOAI22 U21236 ( .A1(n28695), .A2(n2129), .B1(ram[8074]), .B2(n2130), 
        .ZN(n12315) );
  MOAI22 U21237 ( .A1(n28460), .A2(n2129), .B1(ram[8075]), .B2(n2130), 
        .ZN(n12316) );
  MOAI22 U21238 ( .A1(n28225), .A2(n2129), .B1(ram[8076]), .B2(n2130), 
        .ZN(n12317) );
  MOAI22 U21239 ( .A1(n27990), .A2(n2129), .B1(ram[8077]), .B2(n2130), 
        .ZN(n12318) );
  MOAI22 U21240 ( .A1(n27755), .A2(n2129), .B1(ram[8078]), .B2(n2130), 
        .ZN(n12319) );
  MOAI22 U21241 ( .A1(n27520), .A2(n2129), .B1(ram[8079]), .B2(n2130), 
        .ZN(n12320) );
  MOAI22 U21242 ( .A1(n29165), .A2(n2131), .B1(ram[8080]), .B2(n2132), 
        .ZN(n12321) );
  MOAI22 U21243 ( .A1(n28930), .A2(n2131), .B1(ram[8081]), .B2(n2132), 
        .ZN(n12322) );
  MOAI22 U21244 ( .A1(n28695), .A2(n2131), .B1(ram[8082]), .B2(n2132), 
        .ZN(n12323) );
  MOAI22 U21245 ( .A1(n28460), .A2(n2131), .B1(ram[8083]), .B2(n2132), 
        .ZN(n12324) );
  MOAI22 U21246 ( .A1(n28225), .A2(n2131), .B1(ram[8084]), .B2(n2132), 
        .ZN(n12325) );
  MOAI22 U21247 ( .A1(n27990), .A2(n2131), .B1(ram[8085]), .B2(n2132), 
        .ZN(n12326) );
  MOAI22 U21248 ( .A1(n27755), .A2(n2131), .B1(ram[8086]), .B2(n2132), 
        .ZN(n12327) );
  MOAI22 U21249 ( .A1(n27520), .A2(n2131), .B1(ram[8087]), .B2(n2132), 
        .ZN(n12328) );
  MOAI22 U21250 ( .A1(n29165), .A2(n2133), .B1(ram[8088]), .B2(n2134), 
        .ZN(n12329) );
  MOAI22 U21251 ( .A1(n28930), .A2(n2133), .B1(ram[8089]), .B2(n2134), 
        .ZN(n12330) );
  MOAI22 U21252 ( .A1(n28695), .A2(n2133), .B1(ram[8090]), .B2(n2134), 
        .ZN(n12331) );
  MOAI22 U21253 ( .A1(n28460), .A2(n2133), .B1(ram[8091]), .B2(n2134), 
        .ZN(n12332) );
  MOAI22 U21254 ( .A1(n28225), .A2(n2133), .B1(ram[8092]), .B2(n2134), 
        .ZN(n12333) );
  MOAI22 U21255 ( .A1(n27990), .A2(n2133), .B1(ram[8093]), .B2(n2134), 
        .ZN(n12334) );
  MOAI22 U21256 ( .A1(n27755), .A2(n2133), .B1(ram[8094]), .B2(n2134), 
        .ZN(n12335) );
  MOAI22 U21257 ( .A1(n27520), .A2(n2133), .B1(ram[8095]), .B2(n2134), 
        .ZN(n12336) );
  MOAI22 U21258 ( .A1(n29165), .A2(n2135), .B1(ram[8096]), .B2(n2136), 
        .ZN(n12337) );
  MOAI22 U21259 ( .A1(n28930), .A2(n2135), .B1(ram[8097]), .B2(n2136), 
        .ZN(n12338) );
  MOAI22 U21260 ( .A1(n28695), .A2(n2135), .B1(ram[8098]), .B2(n2136), 
        .ZN(n12339) );
  MOAI22 U21261 ( .A1(n28460), .A2(n2135), .B1(ram[8099]), .B2(n2136), 
        .ZN(n12340) );
  MOAI22 U21262 ( .A1(n28225), .A2(n2135), .B1(ram[8100]), .B2(n2136), 
        .ZN(n12341) );
  MOAI22 U21263 ( .A1(n27990), .A2(n2135), .B1(ram[8101]), .B2(n2136), 
        .ZN(n12342) );
  MOAI22 U21264 ( .A1(n27755), .A2(n2135), .B1(ram[8102]), .B2(n2136), 
        .ZN(n12343) );
  MOAI22 U21265 ( .A1(n27520), .A2(n2135), .B1(ram[8103]), .B2(n2136), 
        .ZN(n12344) );
  MOAI22 U21266 ( .A1(n29165), .A2(n2137), .B1(ram[8104]), .B2(n2138), 
        .ZN(n12345) );
  MOAI22 U21267 ( .A1(n28930), .A2(n2137), .B1(ram[8105]), .B2(n2138), 
        .ZN(n12346) );
  MOAI22 U21268 ( .A1(n28695), .A2(n2137), .B1(ram[8106]), .B2(n2138), 
        .ZN(n12347) );
  MOAI22 U21269 ( .A1(n28460), .A2(n2137), .B1(ram[8107]), .B2(n2138), 
        .ZN(n12348) );
  MOAI22 U21270 ( .A1(n28225), .A2(n2137), .B1(ram[8108]), .B2(n2138), 
        .ZN(n12349) );
  MOAI22 U21271 ( .A1(n27990), .A2(n2137), .B1(ram[8109]), .B2(n2138), 
        .ZN(n12350) );
  MOAI22 U21272 ( .A1(n27755), .A2(n2137), .B1(ram[8110]), .B2(n2138), 
        .ZN(n12351) );
  MOAI22 U21273 ( .A1(n27520), .A2(n2137), .B1(ram[8111]), .B2(n2138), 
        .ZN(n12352) );
  MOAI22 U21274 ( .A1(n29166), .A2(n2139), .B1(ram[8112]), .B2(n2140), 
        .ZN(n12353) );
  MOAI22 U21275 ( .A1(n28931), .A2(n2139), .B1(ram[8113]), .B2(n2140), 
        .ZN(n12354) );
  MOAI22 U21276 ( .A1(n28696), .A2(n2139), .B1(ram[8114]), .B2(n2140), 
        .ZN(n12355) );
  MOAI22 U21277 ( .A1(n28461), .A2(n2139), .B1(ram[8115]), .B2(n2140), 
        .ZN(n12356) );
  MOAI22 U21278 ( .A1(n28226), .A2(n2139), .B1(ram[8116]), .B2(n2140), 
        .ZN(n12357) );
  MOAI22 U21279 ( .A1(n27991), .A2(n2139), .B1(ram[8117]), .B2(n2140), 
        .ZN(n12358) );
  MOAI22 U21280 ( .A1(n27756), .A2(n2139), .B1(ram[8118]), .B2(n2140), 
        .ZN(n12359) );
  MOAI22 U21281 ( .A1(n27521), .A2(n2139), .B1(ram[8119]), .B2(n2140), 
        .ZN(n12360) );
  MOAI22 U21282 ( .A1(n29166), .A2(n2141), .B1(ram[8120]), .B2(n2142), 
        .ZN(n12361) );
  MOAI22 U21283 ( .A1(n28931), .A2(n2141), .B1(ram[8121]), .B2(n2142), 
        .ZN(n12362) );
  MOAI22 U21284 ( .A1(n28696), .A2(n2141), .B1(ram[8122]), .B2(n2142), 
        .ZN(n12363) );
  MOAI22 U21285 ( .A1(n28461), .A2(n2141), .B1(ram[8123]), .B2(n2142), 
        .ZN(n12364) );
  MOAI22 U21286 ( .A1(n28226), .A2(n2141), .B1(ram[8124]), .B2(n2142), 
        .ZN(n12365) );
  MOAI22 U21287 ( .A1(n27991), .A2(n2141), .B1(ram[8125]), .B2(n2142), 
        .ZN(n12366) );
  MOAI22 U21288 ( .A1(n27756), .A2(n2141), .B1(ram[8126]), .B2(n2142), 
        .ZN(n12367) );
  MOAI22 U21289 ( .A1(n27521), .A2(n2141), .B1(ram[8127]), .B2(n2142), 
        .ZN(n12368) );
  MOAI22 U21290 ( .A1(n29166), .A2(n2143), .B1(ram[8128]), .B2(n2144), 
        .ZN(n12369) );
  MOAI22 U21291 ( .A1(n28931), .A2(n2143), .B1(ram[8129]), .B2(n2144), 
        .ZN(n12370) );
  MOAI22 U21292 ( .A1(n28696), .A2(n2143), .B1(ram[8130]), .B2(n2144), 
        .ZN(n12371) );
  MOAI22 U21293 ( .A1(n28461), .A2(n2143), .B1(ram[8131]), .B2(n2144), 
        .ZN(n12372) );
  MOAI22 U21294 ( .A1(n28226), .A2(n2143), .B1(ram[8132]), .B2(n2144), 
        .ZN(n12373) );
  MOAI22 U21295 ( .A1(n27991), .A2(n2143), .B1(ram[8133]), .B2(n2144), 
        .ZN(n12374) );
  MOAI22 U21296 ( .A1(n27756), .A2(n2143), .B1(ram[8134]), .B2(n2144), 
        .ZN(n12375) );
  MOAI22 U21297 ( .A1(n27521), .A2(n2143), .B1(ram[8135]), .B2(n2144), 
        .ZN(n12376) );
  MOAI22 U21298 ( .A1(n29166), .A2(n2145), .B1(ram[8136]), .B2(n2146), 
        .ZN(n12377) );
  MOAI22 U21299 ( .A1(n28931), .A2(n2145), .B1(ram[8137]), .B2(n2146), 
        .ZN(n12378) );
  MOAI22 U21300 ( .A1(n28696), .A2(n2145), .B1(ram[8138]), .B2(n2146), 
        .ZN(n12379) );
  MOAI22 U21301 ( .A1(n28461), .A2(n2145), .B1(ram[8139]), .B2(n2146), 
        .ZN(n12380) );
  MOAI22 U21302 ( .A1(n28226), .A2(n2145), .B1(ram[8140]), .B2(n2146), 
        .ZN(n12381) );
  MOAI22 U21303 ( .A1(n27991), .A2(n2145), .B1(ram[8141]), .B2(n2146), 
        .ZN(n12382) );
  MOAI22 U21304 ( .A1(n27756), .A2(n2145), .B1(ram[8142]), .B2(n2146), 
        .ZN(n12383) );
  MOAI22 U21305 ( .A1(n27521), .A2(n2145), .B1(ram[8143]), .B2(n2146), 
        .ZN(n12384) );
  MOAI22 U21306 ( .A1(n29166), .A2(n2147), .B1(ram[8144]), .B2(n2148), 
        .ZN(n12385) );
  MOAI22 U21307 ( .A1(n28931), .A2(n2147), .B1(ram[8145]), .B2(n2148), 
        .ZN(n12386) );
  MOAI22 U21308 ( .A1(n28696), .A2(n2147), .B1(ram[8146]), .B2(n2148), 
        .ZN(n12387) );
  MOAI22 U21309 ( .A1(n28461), .A2(n2147), .B1(ram[8147]), .B2(n2148), 
        .ZN(n12388) );
  MOAI22 U21310 ( .A1(n28226), .A2(n2147), .B1(ram[8148]), .B2(n2148), 
        .ZN(n12389) );
  MOAI22 U21311 ( .A1(n27991), .A2(n2147), .B1(ram[8149]), .B2(n2148), 
        .ZN(n12390) );
  MOAI22 U21312 ( .A1(n27756), .A2(n2147), .B1(ram[8150]), .B2(n2148), 
        .ZN(n12391) );
  MOAI22 U21313 ( .A1(n27521), .A2(n2147), .B1(ram[8151]), .B2(n2148), 
        .ZN(n12392) );
  MOAI22 U21314 ( .A1(n29166), .A2(n2149), .B1(ram[8152]), .B2(n2150), 
        .ZN(n12393) );
  MOAI22 U21315 ( .A1(n28931), .A2(n2149), .B1(ram[8153]), .B2(n2150), 
        .ZN(n12394) );
  MOAI22 U21316 ( .A1(n28696), .A2(n2149), .B1(ram[8154]), .B2(n2150), 
        .ZN(n12395) );
  MOAI22 U21317 ( .A1(n28461), .A2(n2149), .B1(ram[8155]), .B2(n2150), 
        .ZN(n12396) );
  MOAI22 U21318 ( .A1(n28226), .A2(n2149), .B1(ram[8156]), .B2(n2150), 
        .ZN(n12397) );
  MOAI22 U21319 ( .A1(n27991), .A2(n2149), .B1(ram[8157]), .B2(n2150), 
        .ZN(n12398) );
  MOAI22 U21320 ( .A1(n27756), .A2(n2149), .B1(ram[8158]), .B2(n2150), 
        .ZN(n12399) );
  MOAI22 U21321 ( .A1(n27521), .A2(n2149), .B1(ram[8159]), .B2(n2150), 
        .ZN(n12400) );
  MOAI22 U21322 ( .A1(n29166), .A2(n2151), .B1(ram[8160]), .B2(n2152), 
        .ZN(n12401) );
  MOAI22 U21323 ( .A1(n28931), .A2(n2151), .B1(ram[8161]), .B2(n2152), 
        .ZN(n12402) );
  MOAI22 U21324 ( .A1(n28696), .A2(n2151), .B1(ram[8162]), .B2(n2152), 
        .ZN(n12403) );
  MOAI22 U21325 ( .A1(n28461), .A2(n2151), .B1(ram[8163]), .B2(n2152), 
        .ZN(n12404) );
  MOAI22 U21326 ( .A1(n28226), .A2(n2151), .B1(ram[8164]), .B2(n2152), 
        .ZN(n12405) );
  MOAI22 U21327 ( .A1(n27991), .A2(n2151), .B1(ram[8165]), .B2(n2152), 
        .ZN(n12406) );
  MOAI22 U21328 ( .A1(n27756), .A2(n2151), .B1(ram[8166]), .B2(n2152), 
        .ZN(n12407) );
  MOAI22 U21329 ( .A1(n27521), .A2(n2151), .B1(ram[8167]), .B2(n2152), 
        .ZN(n12408) );
  MOAI22 U21330 ( .A1(n29166), .A2(n2153), .B1(ram[8168]), .B2(n2154), 
        .ZN(n12409) );
  MOAI22 U21331 ( .A1(n28931), .A2(n2153), .B1(ram[8169]), .B2(n2154), 
        .ZN(n12410) );
  MOAI22 U21332 ( .A1(n28696), .A2(n2153), .B1(ram[8170]), .B2(n2154), 
        .ZN(n12411) );
  MOAI22 U21333 ( .A1(n28461), .A2(n2153), .B1(ram[8171]), .B2(n2154), 
        .ZN(n12412) );
  MOAI22 U21334 ( .A1(n28226), .A2(n2153), .B1(ram[8172]), .B2(n2154), 
        .ZN(n12413) );
  MOAI22 U21335 ( .A1(n27991), .A2(n2153), .B1(ram[8173]), .B2(n2154), 
        .ZN(n12414) );
  MOAI22 U21336 ( .A1(n27756), .A2(n2153), .B1(ram[8174]), .B2(n2154), 
        .ZN(n12415) );
  MOAI22 U21337 ( .A1(n27521), .A2(n2153), .B1(ram[8175]), .B2(n2154), 
        .ZN(n12416) );
  MOAI22 U21338 ( .A1(n29166), .A2(n2155), .B1(ram[8176]), .B2(n2156), 
        .ZN(n12417) );
  MOAI22 U21339 ( .A1(n28931), .A2(n2155), .B1(ram[8177]), .B2(n2156), 
        .ZN(n12418) );
  MOAI22 U21340 ( .A1(n28696), .A2(n2155), .B1(ram[8178]), .B2(n2156), 
        .ZN(n12419) );
  MOAI22 U21341 ( .A1(n28461), .A2(n2155), .B1(ram[8179]), .B2(n2156), 
        .ZN(n12420) );
  MOAI22 U21342 ( .A1(n28226), .A2(n2155), .B1(ram[8180]), .B2(n2156), 
        .ZN(n12421) );
  MOAI22 U21343 ( .A1(n27991), .A2(n2155), .B1(ram[8181]), .B2(n2156), 
        .ZN(n12422) );
  MOAI22 U21344 ( .A1(n27756), .A2(n2155), .B1(ram[8182]), .B2(n2156), 
        .ZN(n12423) );
  MOAI22 U21345 ( .A1(n27521), .A2(n2155), .B1(ram[8183]), .B2(n2156), 
        .ZN(n12424) );
  MOAI22 U21346 ( .A1(n29166), .A2(n2159), .B1(ram[8192]), .B2(n2160), 
        .ZN(n12433) );
  MOAI22 U21347 ( .A1(n28931), .A2(n2159), .B1(ram[8193]), .B2(n2160), 
        .ZN(n12434) );
  MOAI22 U21348 ( .A1(n28696), .A2(n2159), .B1(ram[8194]), .B2(n2160), 
        .ZN(n12435) );
  MOAI22 U21349 ( .A1(n28461), .A2(n2159), .B1(ram[8195]), .B2(n2160), 
        .ZN(n12436) );
  MOAI22 U21350 ( .A1(n28226), .A2(n2159), .B1(ram[8196]), .B2(n2160), 
        .ZN(n12437) );
  MOAI22 U21351 ( .A1(n27991), .A2(n2159), .B1(ram[8197]), .B2(n2160), 
        .ZN(n12438) );
  MOAI22 U21352 ( .A1(n27756), .A2(n2159), .B1(ram[8198]), .B2(n2160), 
        .ZN(n12439) );
  MOAI22 U21353 ( .A1(n27521), .A2(n2159), .B1(ram[8199]), .B2(n2160), 
        .ZN(n12440) );
  MOAI22 U21354 ( .A1(n29166), .A2(n2162), .B1(ram[8200]), .B2(n2163), 
        .ZN(n12441) );
  MOAI22 U21355 ( .A1(n28931), .A2(n2162), .B1(ram[8201]), .B2(n2163), 
        .ZN(n12442) );
  MOAI22 U21356 ( .A1(n28696), .A2(n2162), .B1(ram[8202]), .B2(n2163), 
        .ZN(n12443) );
  MOAI22 U21357 ( .A1(n28461), .A2(n2162), .B1(ram[8203]), .B2(n2163), 
        .ZN(n12444) );
  MOAI22 U21358 ( .A1(n28226), .A2(n2162), .B1(ram[8204]), .B2(n2163), 
        .ZN(n12445) );
  MOAI22 U21359 ( .A1(n27991), .A2(n2162), .B1(ram[8205]), .B2(n2163), 
        .ZN(n12446) );
  MOAI22 U21360 ( .A1(n27756), .A2(n2162), .B1(ram[8206]), .B2(n2163), 
        .ZN(n12447) );
  MOAI22 U21361 ( .A1(n27521), .A2(n2162), .B1(ram[8207]), .B2(n2163), 
        .ZN(n12448) );
  MOAI22 U21362 ( .A1(n29166), .A2(n2164), .B1(ram[8208]), .B2(n2165), 
        .ZN(n12449) );
  MOAI22 U21363 ( .A1(n28931), .A2(n2164), .B1(ram[8209]), .B2(n2165), 
        .ZN(n12450) );
  MOAI22 U21364 ( .A1(n28696), .A2(n2164), .B1(ram[8210]), .B2(n2165), 
        .ZN(n12451) );
  MOAI22 U21365 ( .A1(n28461), .A2(n2164), .B1(ram[8211]), .B2(n2165), 
        .ZN(n12452) );
  MOAI22 U21366 ( .A1(n28226), .A2(n2164), .B1(ram[8212]), .B2(n2165), 
        .ZN(n12453) );
  MOAI22 U21367 ( .A1(n27991), .A2(n2164), .B1(ram[8213]), .B2(n2165), 
        .ZN(n12454) );
  MOAI22 U21368 ( .A1(n27756), .A2(n2164), .B1(ram[8214]), .B2(n2165), 
        .ZN(n12455) );
  MOAI22 U21369 ( .A1(n27521), .A2(n2164), .B1(ram[8215]), .B2(n2165), 
        .ZN(n12456) );
  MOAI22 U21370 ( .A1(n29167), .A2(n2166), .B1(ram[8216]), .B2(n2167), 
        .ZN(n12457) );
  MOAI22 U21371 ( .A1(n28932), .A2(n2166), .B1(ram[8217]), .B2(n2167), 
        .ZN(n12458) );
  MOAI22 U21372 ( .A1(n28697), .A2(n2166), .B1(ram[8218]), .B2(n2167), 
        .ZN(n12459) );
  MOAI22 U21373 ( .A1(n28462), .A2(n2166), .B1(ram[8219]), .B2(n2167), 
        .ZN(n12460) );
  MOAI22 U21374 ( .A1(n28227), .A2(n2166), .B1(ram[8220]), .B2(n2167), 
        .ZN(n12461) );
  MOAI22 U21375 ( .A1(n27992), .A2(n2166), .B1(ram[8221]), .B2(n2167), 
        .ZN(n12462) );
  MOAI22 U21376 ( .A1(n27757), .A2(n2166), .B1(ram[8222]), .B2(n2167), 
        .ZN(n12463) );
  MOAI22 U21377 ( .A1(n27522), .A2(n2166), .B1(ram[8223]), .B2(n2167), 
        .ZN(n12464) );
  MOAI22 U21378 ( .A1(n29167), .A2(n2168), .B1(ram[8224]), .B2(n2169), 
        .ZN(n12465) );
  MOAI22 U21379 ( .A1(n28932), .A2(n2168), .B1(ram[8225]), .B2(n2169), 
        .ZN(n12466) );
  MOAI22 U21380 ( .A1(n28697), .A2(n2168), .B1(ram[8226]), .B2(n2169), 
        .ZN(n12467) );
  MOAI22 U21381 ( .A1(n28462), .A2(n2168), .B1(ram[8227]), .B2(n2169), 
        .ZN(n12468) );
  MOAI22 U21382 ( .A1(n28227), .A2(n2168), .B1(ram[8228]), .B2(n2169), 
        .ZN(n12469) );
  MOAI22 U21383 ( .A1(n27992), .A2(n2168), .B1(ram[8229]), .B2(n2169), 
        .ZN(n12470) );
  MOAI22 U21384 ( .A1(n27757), .A2(n2168), .B1(ram[8230]), .B2(n2169), 
        .ZN(n12471) );
  MOAI22 U21385 ( .A1(n27522), .A2(n2168), .B1(ram[8231]), .B2(n2169), 
        .ZN(n12472) );
  MOAI22 U21386 ( .A1(n29167), .A2(n2170), .B1(ram[8232]), .B2(n2171), 
        .ZN(n12473) );
  MOAI22 U21387 ( .A1(n28932), .A2(n2170), .B1(ram[8233]), .B2(n2171), 
        .ZN(n12474) );
  MOAI22 U21388 ( .A1(n28697), .A2(n2170), .B1(ram[8234]), .B2(n2171), 
        .ZN(n12475) );
  MOAI22 U21389 ( .A1(n28462), .A2(n2170), .B1(ram[8235]), .B2(n2171), 
        .ZN(n12476) );
  MOAI22 U21390 ( .A1(n28227), .A2(n2170), .B1(ram[8236]), .B2(n2171), 
        .ZN(n12477) );
  MOAI22 U21391 ( .A1(n27992), .A2(n2170), .B1(ram[8237]), .B2(n2171), 
        .ZN(n12478) );
  MOAI22 U21392 ( .A1(n27757), .A2(n2170), .B1(ram[8238]), .B2(n2171), 
        .ZN(n12479) );
  MOAI22 U21393 ( .A1(n27522), .A2(n2170), .B1(ram[8239]), .B2(n2171), 
        .ZN(n12480) );
  MOAI22 U21394 ( .A1(n29167), .A2(n2172), .B1(ram[8240]), .B2(n2173), 
        .ZN(n12481) );
  MOAI22 U21395 ( .A1(n28932), .A2(n2172), .B1(ram[8241]), .B2(n2173), 
        .ZN(n12482) );
  MOAI22 U21396 ( .A1(n28697), .A2(n2172), .B1(ram[8242]), .B2(n2173), 
        .ZN(n12483) );
  MOAI22 U21397 ( .A1(n28462), .A2(n2172), .B1(ram[8243]), .B2(n2173), 
        .ZN(n12484) );
  MOAI22 U21398 ( .A1(n28227), .A2(n2172), .B1(ram[8244]), .B2(n2173), 
        .ZN(n12485) );
  MOAI22 U21399 ( .A1(n27992), .A2(n2172), .B1(ram[8245]), .B2(n2173), 
        .ZN(n12486) );
  MOAI22 U21400 ( .A1(n27757), .A2(n2172), .B1(ram[8246]), .B2(n2173), 
        .ZN(n12487) );
  MOAI22 U21401 ( .A1(n27522), .A2(n2172), .B1(ram[8247]), .B2(n2173), 
        .ZN(n12488) );
  MOAI22 U21402 ( .A1(n29167), .A2(n2174), .B1(ram[8248]), .B2(n2175), 
        .ZN(n12489) );
  MOAI22 U21403 ( .A1(n28932), .A2(n2174), .B1(ram[8249]), .B2(n2175), 
        .ZN(n12490) );
  MOAI22 U21404 ( .A1(n28697), .A2(n2174), .B1(ram[8250]), .B2(n2175), 
        .ZN(n12491) );
  MOAI22 U21405 ( .A1(n28462), .A2(n2174), .B1(ram[8251]), .B2(n2175), 
        .ZN(n12492) );
  MOAI22 U21406 ( .A1(n28227), .A2(n2174), .B1(ram[8252]), .B2(n2175), 
        .ZN(n12493) );
  MOAI22 U21407 ( .A1(n27992), .A2(n2174), .B1(ram[8253]), .B2(n2175), 
        .ZN(n12494) );
  MOAI22 U21408 ( .A1(n27757), .A2(n2174), .B1(ram[8254]), .B2(n2175), 
        .ZN(n12495) );
  MOAI22 U21409 ( .A1(n27522), .A2(n2174), .B1(ram[8255]), .B2(n2175), 
        .ZN(n12496) );
  MOAI22 U21410 ( .A1(n29167), .A2(n2176), .B1(ram[8256]), .B2(n2177), 
        .ZN(n12497) );
  MOAI22 U21411 ( .A1(n28932), .A2(n2176), .B1(ram[8257]), .B2(n2177), 
        .ZN(n12498) );
  MOAI22 U21412 ( .A1(n28697), .A2(n2176), .B1(ram[8258]), .B2(n2177), 
        .ZN(n12499) );
  MOAI22 U21413 ( .A1(n28462), .A2(n2176), .B1(ram[8259]), .B2(n2177), 
        .ZN(n12500) );
  MOAI22 U21414 ( .A1(n28227), .A2(n2176), .B1(ram[8260]), .B2(n2177), 
        .ZN(n12501) );
  MOAI22 U21415 ( .A1(n27992), .A2(n2176), .B1(ram[8261]), .B2(n2177), 
        .ZN(n12502) );
  MOAI22 U21416 ( .A1(n27757), .A2(n2176), .B1(ram[8262]), .B2(n2177), 
        .ZN(n12503) );
  MOAI22 U21417 ( .A1(n27522), .A2(n2176), .B1(ram[8263]), .B2(n2177), 
        .ZN(n12504) );
  MOAI22 U21418 ( .A1(n29167), .A2(n2178), .B1(ram[8264]), .B2(n2179), 
        .ZN(n12505) );
  MOAI22 U21419 ( .A1(n28932), .A2(n2178), .B1(ram[8265]), .B2(n2179), 
        .ZN(n12506) );
  MOAI22 U21420 ( .A1(n28697), .A2(n2178), .B1(ram[8266]), .B2(n2179), 
        .ZN(n12507) );
  MOAI22 U21421 ( .A1(n28462), .A2(n2178), .B1(ram[8267]), .B2(n2179), 
        .ZN(n12508) );
  MOAI22 U21422 ( .A1(n28227), .A2(n2178), .B1(ram[8268]), .B2(n2179), 
        .ZN(n12509) );
  MOAI22 U21423 ( .A1(n27992), .A2(n2178), .B1(ram[8269]), .B2(n2179), 
        .ZN(n12510) );
  MOAI22 U21424 ( .A1(n27757), .A2(n2178), .B1(ram[8270]), .B2(n2179), 
        .ZN(n12511) );
  MOAI22 U21425 ( .A1(n27522), .A2(n2178), .B1(ram[8271]), .B2(n2179), 
        .ZN(n12512) );
  MOAI22 U21426 ( .A1(n29167), .A2(n2180), .B1(ram[8272]), .B2(n2181), 
        .ZN(n12513) );
  MOAI22 U21427 ( .A1(n28932), .A2(n2180), .B1(ram[8273]), .B2(n2181), 
        .ZN(n12514) );
  MOAI22 U21428 ( .A1(n28697), .A2(n2180), .B1(ram[8274]), .B2(n2181), 
        .ZN(n12515) );
  MOAI22 U21429 ( .A1(n28462), .A2(n2180), .B1(ram[8275]), .B2(n2181), 
        .ZN(n12516) );
  MOAI22 U21430 ( .A1(n28227), .A2(n2180), .B1(ram[8276]), .B2(n2181), 
        .ZN(n12517) );
  MOAI22 U21431 ( .A1(n27992), .A2(n2180), .B1(ram[8277]), .B2(n2181), 
        .ZN(n12518) );
  MOAI22 U21432 ( .A1(n27757), .A2(n2180), .B1(ram[8278]), .B2(n2181), 
        .ZN(n12519) );
  MOAI22 U21433 ( .A1(n27522), .A2(n2180), .B1(ram[8279]), .B2(n2181), 
        .ZN(n12520) );
  MOAI22 U21434 ( .A1(n29167), .A2(n2182), .B1(ram[8280]), .B2(n2183), 
        .ZN(n12521) );
  MOAI22 U21435 ( .A1(n28932), .A2(n2182), .B1(ram[8281]), .B2(n2183), 
        .ZN(n12522) );
  MOAI22 U21436 ( .A1(n28697), .A2(n2182), .B1(ram[8282]), .B2(n2183), 
        .ZN(n12523) );
  MOAI22 U21437 ( .A1(n28462), .A2(n2182), .B1(ram[8283]), .B2(n2183), 
        .ZN(n12524) );
  MOAI22 U21438 ( .A1(n28227), .A2(n2182), .B1(ram[8284]), .B2(n2183), 
        .ZN(n12525) );
  MOAI22 U21439 ( .A1(n27992), .A2(n2182), .B1(ram[8285]), .B2(n2183), 
        .ZN(n12526) );
  MOAI22 U21440 ( .A1(n27757), .A2(n2182), .B1(ram[8286]), .B2(n2183), 
        .ZN(n12527) );
  MOAI22 U21441 ( .A1(n27522), .A2(n2182), .B1(ram[8287]), .B2(n2183), 
        .ZN(n12528) );
  MOAI22 U21442 ( .A1(n29167), .A2(n2184), .B1(ram[8288]), .B2(n2185), 
        .ZN(n12529) );
  MOAI22 U21443 ( .A1(n28932), .A2(n2184), .B1(ram[8289]), .B2(n2185), 
        .ZN(n12530) );
  MOAI22 U21444 ( .A1(n28697), .A2(n2184), .B1(ram[8290]), .B2(n2185), 
        .ZN(n12531) );
  MOAI22 U21445 ( .A1(n28462), .A2(n2184), .B1(ram[8291]), .B2(n2185), 
        .ZN(n12532) );
  MOAI22 U21446 ( .A1(n28227), .A2(n2184), .B1(ram[8292]), .B2(n2185), 
        .ZN(n12533) );
  MOAI22 U21447 ( .A1(n27992), .A2(n2184), .B1(ram[8293]), .B2(n2185), 
        .ZN(n12534) );
  MOAI22 U21448 ( .A1(n27757), .A2(n2184), .B1(ram[8294]), .B2(n2185), 
        .ZN(n12535) );
  MOAI22 U21449 ( .A1(n27522), .A2(n2184), .B1(ram[8295]), .B2(n2185), 
        .ZN(n12536) );
  MOAI22 U21450 ( .A1(n29167), .A2(n2186), .B1(ram[8296]), .B2(n2187), 
        .ZN(n12537) );
  MOAI22 U21451 ( .A1(n28932), .A2(n2186), .B1(ram[8297]), .B2(n2187), 
        .ZN(n12538) );
  MOAI22 U21452 ( .A1(n28697), .A2(n2186), .B1(ram[8298]), .B2(n2187), 
        .ZN(n12539) );
  MOAI22 U21453 ( .A1(n28462), .A2(n2186), .B1(ram[8299]), .B2(n2187), 
        .ZN(n12540) );
  MOAI22 U21454 ( .A1(n28227), .A2(n2186), .B1(ram[8300]), .B2(n2187), 
        .ZN(n12541) );
  MOAI22 U21455 ( .A1(n27992), .A2(n2186), .B1(ram[8301]), .B2(n2187), 
        .ZN(n12542) );
  MOAI22 U21456 ( .A1(n27757), .A2(n2186), .B1(ram[8302]), .B2(n2187), 
        .ZN(n12543) );
  MOAI22 U21457 ( .A1(n27522), .A2(n2186), .B1(ram[8303]), .B2(n2187), 
        .ZN(n12544) );
  MOAI22 U21458 ( .A1(n29167), .A2(n2188), .B1(ram[8304]), .B2(n2189), 
        .ZN(n12545) );
  MOAI22 U21459 ( .A1(n28932), .A2(n2188), .B1(ram[8305]), .B2(n2189), 
        .ZN(n12546) );
  MOAI22 U21460 ( .A1(n28697), .A2(n2188), .B1(ram[8306]), .B2(n2189), 
        .ZN(n12547) );
  MOAI22 U21461 ( .A1(n28462), .A2(n2188), .B1(ram[8307]), .B2(n2189), 
        .ZN(n12548) );
  MOAI22 U21462 ( .A1(n28227), .A2(n2188), .B1(ram[8308]), .B2(n2189), 
        .ZN(n12549) );
  MOAI22 U21463 ( .A1(n27992), .A2(n2188), .B1(ram[8309]), .B2(n2189), 
        .ZN(n12550) );
  MOAI22 U21464 ( .A1(n27757), .A2(n2188), .B1(ram[8310]), .B2(n2189), 
        .ZN(n12551) );
  MOAI22 U21465 ( .A1(n27522), .A2(n2188), .B1(ram[8311]), .B2(n2189), 
        .ZN(n12552) );
  MOAI22 U21466 ( .A1(n29167), .A2(n2190), .B1(ram[8312]), .B2(n2191), 
        .ZN(n12553) );
  MOAI22 U21467 ( .A1(n28932), .A2(n2190), .B1(ram[8313]), .B2(n2191), 
        .ZN(n12554) );
  MOAI22 U21468 ( .A1(n28697), .A2(n2190), .B1(ram[8314]), .B2(n2191), 
        .ZN(n12555) );
  MOAI22 U21469 ( .A1(n28462), .A2(n2190), .B1(ram[8315]), .B2(n2191), 
        .ZN(n12556) );
  MOAI22 U21470 ( .A1(n28227), .A2(n2190), .B1(ram[8316]), .B2(n2191), 
        .ZN(n12557) );
  MOAI22 U21471 ( .A1(n27992), .A2(n2190), .B1(ram[8317]), .B2(n2191), 
        .ZN(n12558) );
  MOAI22 U21472 ( .A1(n27757), .A2(n2190), .B1(ram[8318]), .B2(n2191), 
        .ZN(n12559) );
  MOAI22 U21473 ( .A1(n27522), .A2(n2190), .B1(ram[8319]), .B2(n2191), 
        .ZN(n12560) );
  MOAI22 U21474 ( .A1(n29168), .A2(n2192), .B1(ram[8320]), .B2(n2193), 
        .ZN(n12561) );
  MOAI22 U21475 ( .A1(n28933), .A2(n2192), .B1(ram[8321]), .B2(n2193), 
        .ZN(n12562) );
  MOAI22 U21476 ( .A1(n28698), .A2(n2192), .B1(ram[8322]), .B2(n2193), 
        .ZN(n12563) );
  MOAI22 U21477 ( .A1(n28463), .A2(n2192), .B1(ram[8323]), .B2(n2193), 
        .ZN(n12564) );
  MOAI22 U21478 ( .A1(n28228), .A2(n2192), .B1(ram[8324]), .B2(n2193), 
        .ZN(n12565) );
  MOAI22 U21479 ( .A1(n27993), .A2(n2192), .B1(ram[8325]), .B2(n2193), 
        .ZN(n12566) );
  MOAI22 U21480 ( .A1(n27758), .A2(n2192), .B1(ram[8326]), .B2(n2193), 
        .ZN(n12567) );
  MOAI22 U21481 ( .A1(n27523), .A2(n2192), .B1(ram[8327]), .B2(n2193), 
        .ZN(n12568) );
  MOAI22 U21482 ( .A1(n29168), .A2(n2194), .B1(ram[8328]), .B2(n2195), 
        .ZN(n12569) );
  MOAI22 U21483 ( .A1(n28933), .A2(n2194), .B1(ram[8329]), .B2(n2195), 
        .ZN(n12570) );
  MOAI22 U21484 ( .A1(n28698), .A2(n2194), .B1(ram[8330]), .B2(n2195), 
        .ZN(n12571) );
  MOAI22 U21485 ( .A1(n28463), .A2(n2194), .B1(ram[8331]), .B2(n2195), 
        .ZN(n12572) );
  MOAI22 U21486 ( .A1(n28228), .A2(n2194), .B1(ram[8332]), .B2(n2195), 
        .ZN(n12573) );
  MOAI22 U21487 ( .A1(n27993), .A2(n2194), .B1(ram[8333]), .B2(n2195), 
        .ZN(n12574) );
  MOAI22 U21488 ( .A1(n27758), .A2(n2194), .B1(ram[8334]), .B2(n2195), 
        .ZN(n12575) );
  MOAI22 U21489 ( .A1(n27523), .A2(n2194), .B1(ram[8335]), .B2(n2195), 
        .ZN(n12576) );
  MOAI22 U21490 ( .A1(n29168), .A2(n2196), .B1(ram[8336]), .B2(n2197), 
        .ZN(n12577) );
  MOAI22 U21491 ( .A1(n28933), .A2(n2196), .B1(ram[8337]), .B2(n2197), 
        .ZN(n12578) );
  MOAI22 U21492 ( .A1(n28698), .A2(n2196), .B1(ram[8338]), .B2(n2197), 
        .ZN(n12579) );
  MOAI22 U21493 ( .A1(n28463), .A2(n2196), .B1(ram[8339]), .B2(n2197), 
        .ZN(n12580) );
  MOAI22 U21494 ( .A1(n28228), .A2(n2196), .B1(ram[8340]), .B2(n2197), 
        .ZN(n12581) );
  MOAI22 U21495 ( .A1(n27993), .A2(n2196), .B1(ram[8341]), .B2(n2197), 
        .ZN(n12582) );
  MOAI22 U21496 ( .A1(n27758), .A2(n2196), .B1(ram[8342]), .B2(n2197), 
        .ZN(n12583) );
  MOAI22 U21497 ( .A1(n27523), .A2(n2196), .B1(ram[8343]), .B2(n2197), 
        .ZN(n12584) );
  MOAI22 U21498 ( .A1(n29168), .A2(n2198), .B1(ram[8344]), .B2(n2199), 
        .ZN(n12585) );
  MOAI22 U21499 ( .A1(n28933), .A2(n2198), .B1(ram[8345]), .B2(n2199), 
        .ZN(n12586) );
  MOAI22 U21500 ( .A1(n28698), .A2(n2198), .B1(ram[8346]), .B2(n2199), 
        .ZN(n12587) );
  MOAI22 U21501 ( .A1(n28463), .A2(n2198), .B1(ram[8347]), .B2(n2199), 
        .ZN(n12588) );
  MOAI22 U21502 ( .A1(n28228), .A2(n2198), .B1(ram[8348]), .B2(n2199), 
        .ZN(n12589) );
  MOAI22 U21503 ( .A1(n27993), .A2(n2198), .B1(ram[8349]), .B2(n2199), 
        .ZN(n12590) );
  MOAI22 U21504 ( .A1(n27758), .A2(n2198), .B1(ram[8350]), .B2(n2199), 
        .ZN(n12591) );
  MOAI22 U21505 ( .A1(n27523), .A2(n2198), .B1(ram[8351]), .B2(n2199), 
        .ZN(n12592) );
  MOAI22 U21506 ( .A1(n29168), .A2(n2200), .B1(ram[8352]), .B2(n2201), 
        .ZN(n12593) );
  MOAI22 U21507 ( .A1(n28933), .A2(n2200), .B1(ram[8353]), .B2(n2201), 
        .ZN(n12594) );
  MOAI22 U21508 ( .A1(n28698), .A2(n2200), .B1(ram[8354]), .B2(n2201), 
        .ZN(n12595) );
  MOAI22 U21509 ( .A1(n28463), .A2(n2200), .B1(ram[8355]), .B2(n2201), 
        .ZN(n12596) );
  MOAI22 U21510 ( .A1(n28228), .A2(n2200), .B1(ram[8356]), .B2(n2201), 
        .ZN(n12597) );
  MOAI22 U21511 ( .A1(n27993), .A2(n2200), .B1(ram[8357]), .B2(n2201), 
        .ZN(n12598) );
  MOAI22 U21512 ( .A1(n27758), .A2(n2200), .B1(ram[8358]), .B2(n2201), 
        .ZN(n12599) );
  MOAI22 U21513 ( .A1(n27523), .A2(n2200), .B1(ram[8359]), .B2(n2201), 
        .ZN(n12600) );
  MOAI22 U21514 ( .A1(n29168), .A2(n2202), .B1(ram[8360]), .B2(n2203), 
        .ZN(n12601) );
  MOAI22 U21515 ( .A1(n28933), .A2(n2202), .B1(ram[8361]), .B2(n2203), 
        .ZN(n12602) );
  MOAI22 U21516 ( .A1(n28698), .A2(n2202), .B1(ram[8362]), .B2(n2203), 
        .ZN(n12603) );
  MOAI22 U21517 ( .A1(n28463), .A2(n2202), .B1(ram[8363]), .B2(n2203), 
        .ZN(n12604) );
  MOAI22 U21518 ( .A1(n28228), .A2(n2202), .B1(ram[8364]), .B2(n2203), 
        .ZN(n12605) );
  MOAI22 U21519 ( .A1(n27993), .A2(n2202), .B1(ram[8365]), .B2(n2203), 
        .ZN(n12606) );
  MOAI22 U21520 ( .A1(n27758), .A2(n2202), .B1(ram[8366]), .B2(n2203), 
        .ZN(n12607) );
  MOAI22 U21521 ( .A1(n27523), .A2(n2202), .B1(ram[8367]), .B2(n2203), 
        .ZN(n12608) );
  MOAI22 U21522 ( .A1(n29168), .A2(n2204), .B1(ram[8368]), .B2(n2205), 
        .ZN(n12609) );
  MOAI22 U21523 ( .A1(n28933), .A2(n2204), .B1(ram[8369]), .B2(n2205), 
        .ZN(n12610) );
  MOAI22 U21524 ( .A1(n28698), .A2(n2204), .B1(ram[8370]), .B2(n2205), 
        .ZN(n12611) );
  MOAI22 U21525 ( .A1(n28463), .A2(n2204), .B1(ram[8371]), .B2(n2205), 
        .ZN(n12612) );
  MOAI22 U21526 ( .A1(n28228), .A2(n2204), .B1(ram[8372]), .B2(n2205), 
        .ZN(n12613) );
  MOAI22 U21527 ( .A1(n27993), .A2(n2204), .B1(ram[8373]), .B2(n2205), 
        .ZN(n12614) );
  MOAI22 U21528 ( .A1(n27758), .A2(n2204), .B1(ram[8374]), .B2(n2205), 
        .ZN(n12615) );
  MOAI22 U21529 ( .A1(n27523), .A2(n2204), .B1(ram[8375]), .B2(n2205), 
        .ZN(n12616) );
  MOAI22 U21530 ( .A1(n29168), .A2(n2206), .B1(ram[8376]), .B2(n2207), 
        .ZN(n12617) );
  MOAI22 U21531 ( .A1(n28933), .A2(n2206), .B1(ram[8377]), .B2(n2207), 
        .ZN(n12618) );
  MOAI22 U21532 ( .A1(n28698), .A2(n2206), .B1(ram[8378]), .B2(n2207), 
        .ZN(n12619) );
  MOAI22 U21533 ( .A1(n28463), .A2(n2206), .B1(ram[8379]), .B2(n2207), 
        .ZN(n12620) );
  MOAI22 U21534 ( .A1(n28228), .A2(n2206), .B1(ram[8380]), .B2(n2207), 
        .ZN(n12621) );
  MOAI22 U21535 ( .A1(n27993), .A2(n2206), .B1(ram[8381]), .B2(n2207), 
        .ZN(n12622) );
  MOAI22 U21536 ( .A1(n27758), .A2(n2206), .B1(ram[8382]), .B2(n2207), 
        .ZN(n12623) );
  MOAI22 U21537 ( .A1(n27523), .A2(n2206), .B1(ram[8383]), .B2(n2207), 
        .ZN(n12624) );
  MOAI22 U21538 ( .A1(n29168), .A2(n2208), .B1(ram[8384]), .B2(n2209), 
        .ZN(n12625) );
  MOAI22 U21539 ( .A1(n28933), .A2(n2208), .B1(ram[8385]), .B2(n2209), 
        .ZN(n12626) );
  MOAI22 U21540 ( .A1(n28698), .A2(n2208), .B1(ram[8386]), .B2(n2209), 
        .ZN(n12627) );
  MOAI22 U21541 ( .A1(n28463), .A2(n2208), .B1(ram[8387]), .B2(n2209), 
        .ZN(n12628) );
  MOAI22 U21542 ( .A1(n28228), .A2(n2208), .B1(ram[8388]), .B2(n2209), 
        .ZN(n12629) );
  MOAI22 U21543 ( .A1(n27993), .A2(n2208), .B1(ram[8389]), .B2(n2209), 
        .ZN(n12630) );
  MOAI22 U21544 ( .A1(n27758), .A2(n2208), .B1(ram[8390]), .B2(n2209), 
        .ZN(n12631) );
  MOAI22 U21545 ( .A1(n27523), .A2(n2208), .B1(ram[8391]), .B2(n2209), 
        .ZN(n12632) );
  MOAI22 U21546 ( .A1(n29168), .A2(n2210), .B1(ram[8392]), .B2(n2211), 
        .ZN(n12633) );
  MOAI22 U21547 ( .A1(n28933), .A2(n2210), .B1(ram[8393]), .B2(n2211), 
        .ZN(n12634) );
  MOAI22 U21548 ( .A1(n28698), .A2(n2210), .B1(ram[8394]), .B2(n2211), 
        .ZN(n12635) );
  MOAI22 U21549 ( .A1(n28463), .A2(n2210), .B1(ram[8395]), .B2(n2211), 
        .ZN(n12636) );
  MOAI22 U21550 ( .A1(n28228), .A2(n2210), .B1(ram[8396]), .B2(n2211), 
        .ZN(n12637) );
  MOAI22 U21551 ( .A1(n27993), .A2(n2210), .B1(ram[8397]), .B2(n2211), 
        .ZN(n12638) );
  MOAI22 U21552 ( .A1(n27758), .A2(n2210), .B1(ram[8398]), .B2(n2211), 
        .ZN(n12639) );
  MOAI22 U21553 ( .A1(n27523), .A2(n2210), .B1(ram[8399]), .B2(n2211), 
        .ZN(n12640) );
  MOAI22 U21554 ( .A1(n29168), .A2(n2212), .B1(ram[8400]), .B2(n2213), 
        .ZN(n12641) );
  MOAI22 U21555 ( .A1(n28933), .A2(n2212), .B1(ram[8401]), .B2(n2213), 
        .ZN(n12642) );
  MOAI22 U21556 ( .A1(n28698), .A2(n2212), .B1(ram[8402]), .B2(n2213), 
        .ZN(n12643) );
  MOAI22 U21557 ( .A1(n28463), .A2(n2212), .B1(ram[8403]), .B2(n2213), 
        .ZN(n12644) );
  MOAI22 U21558 ( .A1(n28228), .A2(n2212), .B1(ram[8404]), .B2(n2213), 
        .ZN(n12645) );
  MOAI22 U21559 ( .A1(n27993), .A2(n2212), .B1(ram[8405]), .B2(n2213), 
        .ZN(n12646) );
  MOAI22 U21560 ( .A1(n27758), .A2(n2212), .B1(ram[8406]), .B2(n2213), 
        .ZN(n12647) );
  MOAI22 U21561 ( .A1(n27523), .A2(n2212), .B1(ram[8407]), .B2(n2213), 
        .ZN(n12648) );
  MOAI22 U21562 ( .A1(n29168), .A2(n2214), .B1(ram[8408]), .B2(n2215), 
        .ZN(n12649) );
  MOAI22 U21563 ( .A1(n28933), .A2(n2214), .B1(ram[8409]), .B2(n2215), 
        .ZN(n12650) );
  MOAI22 U21564 ( .A1(n28698), .A2(n2214), .B1(ram[8410]), .B2(n2215), 
        .ZN(n12651) );
  MOAI22 U21565 ( .A1(n28463), .A2(n2214), .B1(ram[8411]), .B2(n2215), 
        .ZN(n12652) );
  MOAI22 U21566 ( .A1(n28228), .A2(n2214), .B1(ram[8412]), .B2(n2215), 
        .ZN(n12653) );
  MOAI22 U21567 ( .A1(n27993), .A2(n2214), .B1(ram[8413]), .B2(n2215), 
        .ZN(n12654) );
  MOAI22 U21568 ( .A1(n27758), .A2(n2214), .B1(ram[8414]), .B2(n2215), 
        .ZN(n12655) );
  MOAI22 U21569 ( .A1(n27523), .A2(n2214), .B1(ram[8415]), .B2(n2215), 
        .ZN(n12656) );
  MOAI22 U21570 ( .A1(n29168), .A2(n2216), .B1(ram[8416]), .B2(n2217), 
        .ZN(n12657) );
  MOAI22 U21571 ( .A1(n28933), .A2(n2216), .B1(ram[8417]), .B2(n2217), 
        .ZN(n12658) );
  MOAI22 U21572 ( .A1(n28698), .A2(n2216), .B1(ram[8418]), .B2(n2217), 
        .ZN(n12659) );
  MOAI22 U21573 ( .A1(n28463), .A2(n2216), .B1(ram[8419]), .B2(n2217), 
        .ZN(n12660) );
  MOAI22 U21574 ( .A1(n28228), .A2(n2216), .B1(ram[8420]), .B2(n2217), 
        .ZN(n12661) );
  MOAI22 U21575 ( .A1(n27993), .A2(n2216), .B1(ram[8421]), .B2(n2217), 
        .ZN(n12662) );
  MOAI22 U21576 ( .A1(n27758), .A2(n2216), .B1(ram[8422]), .B2(n2217), 
        .ZN(n12663) );
  MOAI22 U21577 ( .A1(n27523), .A2(n2216), .B1(ram[8423]), .B2(n2217), 
        .ZN(n12664) );
  MOAI22 U21578 ( .A1(n29169), .A2(n2218), .B1(ram[8424]), .B2(n2219), 
        .ZN(n12665) );
  MOAI22 U21579 ( .A1(n28934), .A2(n2218), .B1(ram[8425]), .B2(n2219), 
        .ZN(n12666) );
  MOAI22 U21580 ( .A1(n28699), .A2(n2218), .B1(ram[8426]), .B2(n2219), 
        .ZN(n12667) );
  MOAI22 U21581 ( .A1(n28464), .A2(n2218), .B1(ram[8427]), .B2(n2219), 
        .ZN(n12668) );
  MOAI22 U21582 ( .A1(n28229), .A2(n2218), .B1(ram[8428]), .B2(n2219), 
        .ZN(n12669) );
  MOAI22 U21583 ( .A1(n27994), .A2(n2218), .B1(ram[8429]), .B2(n2219), 
        .ZN(n12670) );
  MOAI22 U21584 ( .A1(n27759), .A2(n2218), .B1(ram[8430]), .B2(n2219), 
        .ZN(n12671) );
  MOAI22 U21585 ( .A1(n27524), .A2(n2218), .B1(ram[8431]), .B2(n2219), 
        .ZN(n12672) );
  MOAI22 U21586 ( .A1(n29169), .A2(n2220), .B1(ram[8432]), .B2(n2221), 
        .ZN(n12673) );
  MOAI22 U21587 ( .A1(n28934), .A2(n2220), .B1(ram[8433]), .B2(n2221), 
        .ZN(n12674) );
  MOAI22 U21588 ( .A1(n28699), .A2(n2220), .B1(ram[8434]), .B2(n2221), 
        .ZN(n12675) );
  MOAI22 U21589 ( .A1(n28464), .A2(n2220), .B1(ram[8435]), .B2(n2221), 
        .ZN(n12676) );
  MOAI22 U21590 ( .A1(n28229), .A2(n2220), .B1(ram[8436]), .B2(n2221), 
        .ZN(n12677) );
  MOAI22 U21591 ( .A1(n27994), .A2(n2220), .B1(ram[8437]), .B2(n2221), 
        .ZN(n12678) );
  MOAI22 U21592 ( .A1(n27759), .A2(n2220), .B1(ram[8438]), .B2(n2221), 
        .ZN(n12679) );
  MOAI22 U21593 ( .A1(n27524), .A2(n2220), .B1(ram[8439]), .B2(n2221), 
        .ZN(n12680) );
  MOAI22 U21594 ( .A1(n29169), .A2(n2222), .B1(ram[8440]), .B2(n2223), 
        .ZN(n12681) );
  MOAI22 U21595 ( .A1(n28934), .A2(n2222), .B1(ram[8441]), .B2(n2223), 
        .ZN(n12682) );
  MOAI22 U21596 ( .A1(n28699), .A2(n2222), .B1(ram[8442]), .B2(n2223), 
        .ZN(n12683) );
  MOAI22 U21597 ( .A1(n28464), .A2(n2222), .B1(ram[8443]), .B2(n2223), 
        .ZN(n12684) );
  MOAI22 U21598 ( .A1(n28229), .A2(n2222), .B1(ram[8444]), .B2(n2223), 
        .ZN(n12685) );
  MOAI22 U21599 ( .A1(n27994), .A2(n2222), .B1(ram[8445]), .B2(n2223), 
        .ZN(n12686) );
  MOAI22 U21600 ( .A1(n27759), .A2(n2222), .B1(ram[8446]), .B2(n2223), 
        .ZN(n12687) );
  MOAI22 U21601 ( .A1(n27524), .A2(n2222), .B1(ram[8447]), .B2(n2223), 
        .ZN(n12688) );
  MOAI22 U21602 ( .A1(n29169), .A2(n2224), .B1(ram[8448]), .B2(n2225), 
        .ZN(n12689) );
  MOAI22 U21603 ( .A1(n28934), .A2(n2224), .B1(ram[8449]), .B2(n2225), 
        .ZN(n12690) );
  MOAI22 U21604 ( .A1(n28699), .A2(n2224), .B1(ram[8450]), .B2(n2225), 
        .ZN(n12691) );
  MOAI22 U21605 ( .A1(n28464), .A2(n2224), .B1(ram[8451]), .B2(n2225), 
        .ZN(n12692) );
  MOAI22 U21606 ( .A1(n28229), .A2(n2224), .B1(ram[8452]), .B2(n2225), 
        .ZN(n12693) );
  MOAI22 U21607 ( .A1(n27994), .A2(n2224), .B1(ram[8453]), .B2(n2225), 
        .ZN(n12694) );
  MOAI22 U21608 ( .A1(n27759), .A2(n2224), .B1(ram[8454]), .B2(n2225), 
        .ZN(n12695) );
  MOAI22 U21609 ( .A1(n27524), .A2(n2224), .B1(ram[8455]), .B2(n2225), 
        .ZN(n12696) );
  MOAI22 U21610 ( .A1(n29169), .A2(n2226), .B1(ram[8456]), .B2(n2227), 
        .ZN(n12697) );
  MOAI22 U21611 ( .A1(n28934), .A2(n2226), .B1(ram[8457]), .B2(n2227), 
        .ZN(n12698) );
  MOAI22 U21612 ( .A1(n28699), .A2(n2226), .B1(ram[8458]), .B2(n2227), 
        .ZN(n12699) );
  MOAI22 U21613 ( .A1(n28464), .A2(n2226), .B1(ram[8459]), .B2(n2227), 
        .ZN(n12700) );
  MOAI22 U21614 ( .A1(n28229), .A2(n2226), .B1(ram[8460]), .B2(n2227), 
        .ZN(n12701) );
  MOAI22 U21615 ( .A1(n27994), .A2(n2226), .B1(ram[8461]), .B2(n2227), 
        .ZN(n12702) );
  MOAI22 U21616 ( .A1(n27759), .A2(n2226), .B1(ram[8462]), .B2(n2227), 
        .ZN(n12703) );
  MOAI22 U21617 ( .A1(n27524), .A2(n2226), .B1(ram[8463]), .B2(n2227), 
        .ZN(n12704) );
  MOAI22 U21618 ( .A1(n29169), .A2(n2228), .B1(ram[8464]), .B2(n2229), 
        .ZN(n12705) );
  MOAI22 U21619 ( .A1(n28934), .A2(n2228), .B1(ram[8465]), .B2(n2229), 
        .ZN(n12706) );
  MOAI22 U21620 ( .A1(n28699), .A2(n2228), .B1(ram[8466]), .B2(n2229), 
        .ZN(n12707) );
  MOAI22 U21621 ( .A1(n28464), .A2(n2228), .B1(ram[8467]), .B2(n2229), 
        .ZN(n12708) );
  MOAI22 U21622 ( .A1(n28229), .A2(n2228), .B1(ram[8468]), .B2(n2229), 
        .ZN(n12709) );
  MOAI22 U21623 ( .A1(n27994), .A2(n2228), .B1(ram[8469]), .B2(n2229), 
        .ZN(n12710) );
  MOAI22 U21624 ( .A1(n27759), .A2(n2228), .B1(ram[8470]), .B2(n2229), 
        .ZN(n12711) );
  MOAI22 U21625 ( .A1(n27524), .A2(n2228), .B1(ram[8471]), .B2(n2229), 
        .ZN(n12712) );
  MOAI22 U21626 ( .A1(n29169), .A2(n2230), .B1(ram[8472]), .B2(n2231), 
        .ZN(n12713) );
  MOAI22 U21627 ( .A1(n28934), .A2(n2230), .B1(ram[8473]), .B2(n2231), 
        .ZN(n12714) );
  MOAI22 U21628 ( .A1(n28699), .A2(n2230), .B1(ram[8474]), .B2(n2231), 
        .ZN(n12715) );
  MOAI22 U21629 ( .A1(n28464), .A2(n2230), .B1(ram[8475]), .B2(n2231), 
        .ZN(n12716) );
  MOAI22 U21630 ( .A1(n28229), .A2(n2230), .B1(ram[8476]), .B2(n2231), 
        .ZN(n12717) );
  MOAI22 U21631 ( .A1(n27994), .A2(n2230), .B1(ram[8477]), .B2(n2231), 
        .ZN(n12718) );
  MOAI22 U21632 ( .A1(n27759), .A2(n2230), .B1(ram[8478]), .B2(n2231), 
        .ZN(n12719) );
  MOAI22 U21633 ( .A1(n27524), .A2(n2230), .B1(ram[8479]), .B2(n2231), 
        .ZN(n12720) );
  MOAI22 U21634 ( .A1(n29169), .A2(n2232), .B1(ram[8480]), .B2(n2233), 
        .ZN(n12721) );
  MOAI22 U21635 ( .A1(n28934), .A2(n2232), .B1(ram[8481]), .B2(n2233), 
        .ZN(n12722) );
  MOAI22 U21636 ( .A1(n28699), .A2(n2232), .B1(ram[8482]), .B2(n2233), 
        .ZN(n12723) );
  MOAI22 U21637 ( .A1(n28464), .A2(n2232), .B1(ram[8483]), .B2(n2233), 
        .ZN(n12724) );
  MOAI22 U21638 ( .A1(n28229), .A2(n2232), .B1(ram[8484]), .B2(n2233), 
        .ZN(n12725) );
  MOAI22 U21639 ( .A1(n27994), .A2(n2232), .B1(ram[8485]), .B2(n2233), 
        .ZN(n12726) );
  MOAI22 U21640 ( .A1(n27759), .A2(n2232), .B1(ram[8486]), .B2(n2233), 
        .ZN(n12727) );
  MOAI22 U21641 ( .A1(n27524), .A2(n2232), .B1(ram[8487]), .B2(n2233), 
        .ZN(n12728) );
  MOAI22 U21642 ( .A1(n29169), .A2(n2234), .B1(ram[8488]), .B2(n2235), 
        .ZN(n12729) );
  MOAI22 U21643 ( .A1(n28934), .A2(n2234), .B1(ram[8489]), .B2(n2235), 
        .ZN(n12730) );
  MOAI22 U21644 ( .A1(n28699), .A2(n2234), .B1(ram[8490]), .B2(n2235), 
        .ZN(n12731) );
  MOAI22 U21645 ( .A1(n28464), .A2(n2234), .B1(ram[8491]), .B2(n2235), 
        .ZN(n12732) );
  MOAI22 U21646 ( .A1(n28229), .A2(n2234), .B1(ram[8492]), .B2(n2235), 
        .ZN(n12733) );
  MOAI22 U21647 ( .A1(n27994), .A2(n2234), .B1(ram[8493]), .B2(n2235), 
        .ZN(n12734) );
  MOAI22 U21648 ( .A1(n27759), .A2(n2234), .B1(ram[8494]), .B2(n2235), 
        .ZN(n12735) );
  MOAI22 U21649 ( .A1(n27524), .A2(n2234), .B1(ram[8495]), .B2(n2235), 
        .ZN(n12736) );
  MOAI22 U21650 ( .A1(n29169), .A2(n2236), .B1(ram[8496]), .B2(n2237), 
        .ZN(n12737) );
  MOAI22 U21651 ( .A1(n28934), .A2(n2236), .B1(ram[8497]), .B2(n2237), 
        .ZN(n12738) );
  MOAI22 U21652 ( .A1(n28699), .A2(n2236), .B1(ram[8498]), .B2(n2237), 
        .ZN(n12739) );
  MOAI22 U21653 ( .A1(n28464), .A2(n2236), .B1(ram[8499]), .B2(n2237), 
        .ZN(n12740) );
  MOAI22 U21654 ( .A1(n28229), .A2(n2236), .B1(ram[8500]), .B2(n2237), 
        .ZN(n12741) );
  MOAI22 U21655 ( .A1(n27994), .A2(n2236), .B1(ram[8501]), .B2(n2237), 
        .ZN(n12742) );
  MOAI22 U21656 ( .A1(n27759), .A2(n2236), .B1(ram[8502]), .B2(n2237), 
        .ZN(n12743) );
  MOAI22 U21657 ( .A1(n27524), .A2(n2236), .B1(ram[8503]), .B2(n2237), 
        .ZN(n12744) );
  MOAI22 U21658 ( .A1(n29169), .A2(n2238), .B1(ram[8504]), .B2(n2239), 
        .ZN(n12745) );
  MOAI22 U21659 ( .A1(n28934), .A2(n2238), .B1(ram[8505]), .B2(n2239), 
        .ZN(n12746) );
  MOAI22 U21660 ( .A1(n28699), .A2(n2238), .B1(ram[8506]), .B2(n2239), 
        .ZN(n12747) );
  MOAI22 U21661 ( .A1(n28464), .A2(n2238), .B1(ram[8507]), .B2(n2239), 
        .ZN(n12748) );
  MOAI22 U21662 ( .A1(n28229), .A2(n2238), .B1(ram[8508]), .B2(n2239), 
        .ZN(n12749) );
  MOAI22 U21663 ( .A1(n27994), .A2(n2238), .B1(ram[8509]), .B2(n2239), 
        .ZN(n12750) );
  MOAI22 U21664 ( .A1(n27759), .A2(n2238), .B1(ram[8510]), .B2(n2239), 
        .ZN(n12751) );
  MOAI22 U21665 ( .A1(n27524), .A2(n2238), .B1(ram[8511]), .B2(n2239), 
        .ZN(n12752) );
  MOAI22 U21666 ( .A1(n29169), .A2(n2240), .B1(ram[8512]), .B2(n2241), 
        .ZN(n12753) );
  MOAI22 U21667 ( .A1(n28934), .A2(n2240), .B1(ram[8513]), .B2(n2241), 
        .ZN(n12754) );
  MOAI22 U21668 ( .A1(n28699), .A2(n2240), .B1(ram[8514]), .B2(n2241), 
        .ZN(n12755) );
  MOAI22 U21669 ( .A1(n28464), .A2(n2240), .B1(ram[8515]), .B2(n2241), 
        .ZN(n12756) );
  MOAI22 U21670 ( .A1(n28229), .A2(n2240), .B1(ram[8516]), .B2(n2241), 
        .ZN(n12757) );
  MOAI22 U21671 ( .A1(n27994), .A2(n2240), .B1(ram[8517]), .B2(n2241), 
        .ZN(n12758) );
  MOAI22 U21672 ( .A1(n27759), .A2(n2240), .B1(ram[8518]), .B2(n2241), 
        .ZN(n12759) );
  MOAI22 U21673 ( .A1(n27524), .A2(n2240), .B1(ram[8519]), .B2(n2241), 
        .ZN(n12760) );
  MOAI22 U21674 ( .A1(n29169), .A2(n2242), .B1(ram[8520]), .B2(n2243), 
        .ZN(n12761) );
  MOAI22 U21675 ( .A1(n28934), .A2(n2242), .B1(ram[8521]), .B2(n2243), 
        .ZN(n12762) );
  MOAI22 U21676 ( .A1(n28699), .A2(n2242), .B1(ram[8522]), .B2(n2243), 
        .ZN(n12763) );
  MOAI22 U21677 ( .A1(n28464), .A2(n2242), .B1(ram[8523]), .B2(n2243), 
        .ZN(n12764) );
  MOAI22 U21678 ( .A1(n28229), .A2(n2242), .B1(ram[8524]), .B2(n2243), 
        .ZN(n12765) );
  MOAI22 U21679 ( .A1(n27994), .A2(n2242), .B1(ram[8525]), .B2(n2243), 
        .ZN(n12766) );
  MOAI22 U21680 ( .A1(n27759), .A2(n2242), .B1(ram[8526]), .B2(n2243), 
        .ZN(n12767) );
  MOAI22 U21681 ( .A1(n27524), .A2(n2242), .B1(ram[8527]), .B2(n2243), 
        .ZN(n12768) );
  MOAI22 U21682 ( .A1(n29170), .A2(n2244), .B1(ram[8528]), .B2(n2245), 
        .ZN(n12769) );
  MOAI22 U21683 ( .A1(n28935), .A2(n2244), .B1(ram[8529]), .B2(n2245), 
        .ZN(n12770) );
  MOAI22 U21684 ( .A1(n28700), .A2(n2244), .B1(ram[8530]), .B2(n2245), 
        .ZN(n12771) );
  MOAI22 U21685 ( .A1(n28465), .A2(n2244), .B1(ram[8531]), .B2(n2245), 
        .ZN(n12772) );
  MOAI22 U21686 ( .A1(n28230), .A2(n2244), .B1(ram[8532]), .B2(n2245), 
        .ZN(n12773) );
  MOAI22 U21687 ( .A1(n27995), .A2(n2244), .B1(ram[8533]), .B2(n2245), 
        .ZN(n12774) );
  MOAI22 U21688 ( .A1(n27760), .A2(n2244), .B1(ram[8534]), .B2(n2245), 
        .ZN(n12775) );
  MOAI22 U21689 ( .A1(n27525), .A2(n2244), .B1(ram[8535]), .B2(n2245), 
        .ZN(n12776) );
  MOAI22 U21690 ( .A1(n29170), .A2(n2246), .B1(ram[8536]), .B2(n2247), 
        .ZN(n12777) );
  MOAI22 U21691 ( .A1(n28935), .A2(n2246), .B1(ram[8537]), .B2(n2247), 
        .ZN(n12778) );
  MOAI22 U21692 ( .A1(n28700), .A2(n2246), .B1(ram[8538]), .B2(n2247), 
        .ZN(n12779) );
  MOAI22 U21693 ( .A1(n28465), .A2(n2246), .B1(ram[8539]), .B2(n2247), 
        .ZN(n12780) );
  MOAI22 U21694 ( .A1(n28230), .A2(n2246), .B1(ram[8540]), .B2(n2247), 
        .ZN(n12781) );
  MOAI22 U21695 ( .A1(n27995), .A2(n2246), .B1(ram[8541]), .B2(n2247), 
        .ZN(n12782) );
  MOAI22 U21696 ( .A1(n27760), .A2(n2246), .B1(ram[8542]), .B2(n2247), 
        .ZN(n12783) );
  MOAI22 U21697 ( .A1(n27525), .A2(n2246), .B1(ram[8543]), .B2(n2247), 
        .ZN(n12784) );
  MOAI22 U21698 ( .A1(n29170), .A2(n2248), .B1(ram[8544]), .B2(n2249), 
        .ZN(n12785) );
  MOAI22 U21699 ( .A1(n28935), .A2(n2248), .B1(ram[8545]), .B2(n2249), 
        .ZN(n12786) );
  MOAI22 U21700 ( .A1(n28700), .A2(n2248), .B1(ram[8546]), .B2(n2249), 
        .ZN(n12787) );
  MOAI22 U21701 ( .A1(n28465), .A2(n2248), .B1(ram[8547]), .B2(n2249), 
        .ZN(n12788) );
  MOAI22 U21702 ( .A1(n28230), .A2(n2248), .B1(ram[8548]), .B2(n2249), 
        .ZN(n12789) );
  MOAI22 U21703 ( .A1(n27995), .A2(n2248), .B1(ram[8549]), .B2(n2249), 
        .ZN(n12790) );
  MOAI22 U21704 ( .A1(n27760), .A2(n2248), .B1(ram[8550]), .B2(n2249), 
        .ZN(n12791) );
  MOAI22 U21705 ( .A1(n27525), .A2(n2248), .B1(ram[8551]), .B2(n2249), 
        .ZN(n12792) );
  MOAI22 U21706 ( .A1(n29170), .A2(n2250), .B1(ram[8552]), .B2(n2251), 
        .ZN(n12793) );
  MOAI22 U21707 ( .A1(n28935), .A2(n2250), .B1(ram[8553]), .B2(n2251), 
        .ZN(n12794) );
  MOAI22 U21708 ( .A1(n28700), .A2(n2250), .B1(ram[8554]), .B2(n2251), 
        .ZN(n12795) );
  MOAI22 U21709 ( .A1(n28465), .A2(n2250), .B1(ram[8555]), .B2(n2251), 
        .ZN(n12796) );
  MOAI22 U21710 ( .A1(n28230), .A2(n2250), .B1(ram[8556]), .B2(n2251), 
        .ZN(n12797) );
  MOAI22 U21711 ( .A1(n27995), .A2(n2250), .B1(ram[8557]), .B2(n2251), 
        .ZN(n12798) );
  MOAI22 U21712 ( .A1(n27760), .A2(n2250), .B1(ram[8558]), .B2(n2251), 
        .ZN(n12799) );
  MOAI22 U21713 ( .A1(n27525), .A2(n2250), .B1(ram[8559]), .B2(n2251), 
        .ZN(n12800) );
  MOAI22 U21714 ( .A1(n29170), .A2(n2252), .B1(ram[8560]), .B2(n2253), 
        .ZN(n12801) );
  MOAI22 U21715 ( .A1(n28935), .A2(n2252), .B1(ram[8561]), .B2(n2253), 
        .ZN(n12802) );
  MOAI22 U21716 ( .A1(n28700), .A2(n2252), .B1(ram[8562]), .B2(n2253), 
        .ZN(n12803) );
  MOAI22 U21717 ( .A1(n28465), .A2(n2252), .B1(ram[8563]), .B2(n2253), 
        .ZN(n12804) );
  MOAI22 U21718 ( .A1(n28230), .A2(n2252), .B1(ram[8564]), .B2(n2253), 
        .ZN(n12805) );
  MOAI22 U21719 ( .A1(n27995), .A2(n2252), .B1(ram[8565]), .B2(n2253), 
        .ZN(n12806) );
  MOAI22 U21720 ( .A1(n27760), .A2(n2252), .B1(ram[8566]), .B2(n2253), 
        .ZN(n12807) );
  MOAI22 U21721 ( .A1(n27525), .A2(n2252), .B1(ram[8567]), .B2(n2253), 
        .ZN(n12808) );
  MOAI22 U21722 ( .A1(n29170), .A2(n2254), .B1(ram[8568]), .B2(n2255), 
        .ZN(n12809) );
  MOAI22 U21723 ( .A1(n28935), .A2(n2254), .B1(ram[8569]), .B2(n2255), 
        .ZN(n12810) );
  MOAI22 U21724 ( .A1(n28700), .A2(n2254), .B1(ram[8570]), .B2(n2255), 
        .ZN(n12811) );
  MOAI22 U21725 ( .A1(n28465), .A2(n2254), .B1(ram[8571]), .B2(n2255), 
        .ZN(n12812) );
  MOAI22 U21726 ( .A1(n28230), .A2(n2254), .B1(ram[8572]), .B2(n2255), 
        .ZN(n12813) );
  MOAI22 U21727 ( .A1(n27995), .A2(n2254), .B1(ram[8573]), .B2(n2255), 
        .ZN(n12814) );
  MOAI22 U21728 ( .A1(n27760), .A2(n2254), .B1(ram[8574]), .B2(n2255), 
        .ZN(n12815) );
  MOAI22 U21729 ( .A1(n27525), .A2(n2254), .B1(ram[8575]), .B2(n2255), 
        .ZN(n12816) );
  MOAI22 U21730 ( .A1(n29170), .A2(n2256), .B1(ram[8576]), .B2(n2257), 
        .ZN(n12817) );
  MOAI22 U21731 ( .A1(n28935), .A2(n2256), .B1(ram[8577]), .B2(n2257), 
        .ZN(n12818) );
  MOAI22 U21732 ( .A1(n28700), .A2(n2256), .B1(ram[8578]), .B2(n2257), 
        .ZN(n12819) );
  MOAI22 U21733 ( .A1(n28465), .A2(n2256), .B1(ram[8579]), .B2(n2257), 
        .ZN(n12820) );
  MOAI22 U21734 ( .A1(n28230), .A2(n2256), .B1(ram[8580]), .B2(n2257), 
        .ZN(n12821) );
  MOAI22 U21735 ( .A1(n27995), .A2(n2256), .B1(ram[8581]), .B2(n2257), 
        .ZN(n12822) );
  MOAI22 U21736 ( .A1(n27760), .A2(n2256), .B1(ram[8582]), .B2(n2257), 
        .ZN(n12823) );
  MOAI22 U21737 ( .A1(n27525), .A2(n2256), .B1(ram[8583]), .B2(n2257), 
        .ZN(n12824) );
  MOAI22 U21738 ( .A1(n29170), .A2(n2258), .B1(ram[8584]), .B2(n2259), 
        .ZN(n12825) );
  MOAI22 U21739 ( .A1(n28935), .A2(n2258), .B1(ram[8585]), .B2(n2259), 
        .ZN(n12826) );
  MOAI22 U21740 ( .A1(n28700), .A2(n2258), .B1(ram[8586]), .B2(n2259), 
        .ZN(n12827) );
  MOAI22 U21741 ( .A1(n28465), .A2(n2258), .B1(ram[8587]), .B2(n2259), 
        .ZN(n12828) );
  MOAI22 U21742 ( .A1(n28230), .A2(n2258), .B1(ram[8588]), .B2(n2259), 
        .ZN(n12829) );
  MOAI22 U21743 ( .A1(n27995), .A2(n2258), .B1(ram[8589]), .B2(n2259), 
        .ZN(n12830) );
  MOAI22 U21744 ( .A1(n27760), .A2(n2258), .B1(ram[8590]), .B2(n2259), 
        .ZN(n12831) );
  MOAI22 U21745 ( .A1(n27525), .A2(n2258), .B1(ram[8591]), .B2(n2259), 
        .ZN(n12832) );
  MOAI22 U21746 ( .A1(n29170), .A2(n2260), .B1(ram[8592]), .B2(n2261), 
        .ZN(n12833) );
  MOAI22 U21747 ( .A1(n28935), .A2(n2260), .B1(ram[8593]), .B2(n2261), 
        .ZN(n12834) );
  MOAI22 U21748 ( .A1(n28700), .A2(n2260), .B1(ram[8594]), .B2(n2261), 
        .ZN(n12835) );
  MOAI22 U21749 ( .A1(n28465), .A2(n2260), .B1(ram[8595]), .B2(n2261), 
        .ZN(n12836) );
  MOAI22 U21750 ( .A1(n28230), .A2(n2260), .B1(ram[8596]), .B2(n2261), 
        .ZN(n12837) );
  MOAI22 U21751 ( .A1(n27995), .A2(n2260), .B1(ram[8597]), .B2(n2261), 
        .ZN(n12838) );
  MOAI22 U21752 ( .A1(n27760), .A2(n2260), .B1(ram[8598]), .B2(n2261), 
        .ZN(n12839) );
  MOAI22 U21753 ( .A1(n27525), .A2(n2260), .B1(ram[8599]), .B2(n2261), 
        .ZN(n12840) );
  MOAI22 U21754 ( .A1(n29170), .A2(n2262), .B1(ram[8600]), .B2(n2263), 
        .ZN(n12841) );
  MOAI22 U21755 ( .A1(n28935), .A2(n2262), .B1(ram[8601]), .B2(n2263), 
        .ZN(n12842) );
  MOAI22 U21756 ( .A1(n28700), .A2(n2262), .B1(ram[8602]), .B2(n2263), 
        .ZN(n12843) );
  MOAI22 U21757 ( .A1(n28465), .A2(n2262), .B1(ram[8603]), .B2(n2263), 
        .ZN(n12844) );
  MOAI22 U21758 ( .A1(n28230), .A2(n2262), .B1(ram[8604]), .B2(n2263), 
        .ZN(n12845) );
  MOAI22 U21759 ( .A1(n27995), .A2(n2262), .B1(ram[8605]), .B2(n2263), 
        .ZN(n12846) );
  MOAI22 U21760 ( .A1(n27760), .A2(n2262), .B1(ram[8606]), .B2(n2263), 
        .ZN(n12847) );
  MOAI22 U21761 ( .A1(n27525), .A2(n2262), .B1(ram[8607]), .B2(n2263), 
        .ZN(n12848) );
  MOAI22 U21762 ( .A1(n29170), .A2(n2264), .B1(ram[8608]), .B2(n2265), 
        .ZN(n12849) );
  MOAI22 U21763 ( .A1(n28935), .A2(n2264), .B1(ram[8609]), .B2(n2265), 
        .ZN(n12850) );
  MOAI22 U21764 ( .A1(n28700), .A2(n2264), .B1(ram[8610]), .B2(n2265), 
        .ZN(n12851) );
  MOAI22 U21765 ( .A1(n28465), .A2(n2264), .B1(ram[8611]), .B2(n2265), 
        .ZN(n12852) );
  MOAI22 U21766 ( .A1(n28230), .A2(n2264), .B1(ram[8612]), .B2(n2265), 
        .ZN(n12853) );
  MOAI22 U21767 ( .A1(n27995), .A2(n2264), .B1(ram[8613]), .B2(n2265), 
        .ZN(n12854) );
  MOAI22 U21768 ( .A1(n27760), .A2(n2264), .B1(ram[8614]), .B2(n2265), 
        .ZN(n12855) );
  MOAI22 U21769 ( .A1(n27525), .A2(n2264), .B1(ram[8615]), .B2(n2265), 
        .ZN(n12856) );
  MOAI22 U21770 ( .A1(n29170), .A2(n2266), .B1(ram[8616]), .B2(n2267), 
        .ZN(n12857) );
  MOAI22 U21771 ( .A1(n28935), .A2(n2266), .B1(ram[8617]), .B2(n2267), 
        .ZN(n12858) );
  MOAI22 U21772 ( .A1(n28700), .A2(n2266), .B1(ram[8618]), .B2(n2267), 
        .ZN(n12859) );
  MOAI22 U21773 ( .A1(n28465), .A2(n2266), .B1(ram[8619]), .B2(n2267), 
        .ZN(n12860) );
  MOAI22 U21774 ( .A1(n28230), .A2(n2266), .B1(ram[8620]), .B2(n2267), 
        .ZN(n12861) );
  MOAI22 U21775 ( .A1(n27995), .A2(n2266), .B1(ram[8621]), .B2(n2267), 
        .ZN(n12862) );
  MOAI22 U21776 ( .A1(n27760), .A2(n2266), .B1(ram[8622]), .B2(n2267), 
        .ZN(n12863) );
  MOAI22 U21777 ( .A1(n27525), .A2(n2266), .B1(ram[8623]), .B2(n2267), 
        .ZN(n12864) );
  MOAI22 U21778 ( .A1(n29170), .A2(n2268), .B1(ram[8624]), .B2(n2269), 
        .ZN(n12865) );
  MOAI22 U21779 ( .A1(n28935), .A2(n2268), .B1(ram[8625]), .B2(n2269), 
        .ZN(n12866) );
  MOAI22 U21780 ( .A1(n28700), .A2(n2268), .B1(ram[8626]), .B2(n2269), 
        .ZN(n12867) );
  MOAI22 U21781 ( .A1(n28465), .A2(n2268), .B1(ram[8627]), .B2(n2269), 
        .ZN(n12868) );
  MOAI22 U21782 ( .A1(n28230), .A2(n2268), .B1(ram[8628]), .B2(n2269), 
        .ZN(n12869) );
  MOAI22 U21783 ( .A1(n27995), .A2(n2268), .B1(ram[8629]), .B2(n2269), 
        .ZN(n12870) );
  MOAI22 U21784 ( .A1(n27760), .A2(n2268), .B1(ram[8630]), .B2(n2269), 
        .ZN(n12871) );
  MOAI22 U21785 ( .A1(n27525), .A2(n2268), .B1(ram[8631]), .B2(n2269), 
        .ZN(n12872) );
  MOAI22 U21786 ( .A1(n29171), .A2(n2270), .B1(ram[8632]), .B2(n2271), 
        .ZN(n12873) );
  MOAI22 U21787 ( .A1(n28936), .A2(n2270), .B1(ram[8633]), .B2(n2271), 
        .ZN(n12874) );
  MOAI22 U21788 ( .A1(n28701), .A2(n2270), .B1(ram[8634]), .B2(n2271), 
        .ZN(n12875) );
  MOAI22 U21789 ( .A1(n28466), .A2(n2270), .B1(ram[8635]), .B2(n2271), 
        .ZN(n12876) );
  MOAI22 U21790 ( .A1(n28231), .A2(n2270), .B1(ram[8636]), .B2(n2271), 
        .ZN(n12877) );
  MOAI22 U21791 ( .A1(n27996), .A2(n2270), .B1(ram[8637]), .B2(n2271), 
        .ZN(n12878) );
  MOAI22 U21792 ( .A1(n27761), .A2(n2270), .B1(ram[8638]), .B2(n2271), 
        .ZN(n12879) );
  MOAI22 U21793 ( .A1(n27526), .A2(n2270), .B1(ram[8639]), .B2(n2271), 
        .ZN(n12880) );
  MOAI22 U21794 ( .A1(n29171), .A2(n2272), .B1(ram[8640]), .B2(n2273), 
        .ZN(n12881) );
  MOAI22 U21795 ( .A1(n28936), .A2(n2272), .B1(ram[8641]), .B2(n2273), 
        .ZN(n12882) );
  MOAI22 U21796 ( .A1(n28701), .A2(n2272), .B1(ram[8642]), .B2(n2273), 
        .ZN(n12883) );
  MOAI22 U21797 ( .A1(n28466), .A2(n2272), .B1(ram[8643]), .B2(n2273), 
        .ZN(n12884) );
  MOAI22 U21798 ( .A1(n28231), .A2(n2272), .B1(ram[8644]), .B2(n2273), 
        .ZN(n12885) );
  MOAI22 U21799 ( .A1(n27996), .A2(n2272), .B1(ram[8645]), .B2(n2273), 
        .ZN(n12886) );
  MOAI22 U21800 ( .A1(n27761), .A2(n2272), .B1(ram[8646]), .B2(n2273), 
        .ZN(n12887) );
  MOAI22 U21801 ( .A1(n27526), .A2(n2272), .B1(ram[8647]), .B2(n2273), 
        .ZN(n12888) );
  MOAI22 U21802 ( .A1(n29171), .A2(n2274), .B1(ram[8648]), .B2(n2275), 
        .ZN(n12889) );
  MOAI22 U21803 ( .A1(n28936), .A2(n2274), .B1(ram[8649]), .B2(n2275), 
        .ZN(n12890) );
  MOAI22 U21804 ( .A1(n28701), .A2(n2274), .B1(ram[8650]), .B2(n2275), 
        .ZN(n12891) );
  MOAI22 U21805 ( .A1(n28466), .A2(n2274), .B1(ram[8651]), .B2(n2275), 
        .ZN(n12892) );
  MOAI22 U21806 ( .A1(n28231), .A2(n2274), .B1(ram[8652]), .B2(n2275), 
        .ZN(n12893) );
  MOAI22 U21807 ( .A1(n27996), .A2(n2274), .B1(ram[8653]), .B2(n2275), 
        .ZN(n12894) );
  MOAI22 U21808 ( .A1(n27761), .A2(n2274), .B1(ram[8654]), .B2(n2275), 
        .ZN(n12895) );
  MOAI22 U21809 ( .A1(n27526), .A2(n2274), .B1(ram[8655]), .B2(n2275), 
        .ZN(n12896) );
  MOAI22 U21810 ( .A1(n29171), .A2(n2276), .B1(ram[8656]), .B2(n2277), 
        .ZN(n12897) );
  MOAI22 U21811 ( .A1(n28936), .A2(n2276), .B1(ram[8657]), .B2(n2277), 
        .ZN(n12898) );
  MOAI22 U21812 ( .A1(n28701), .A2(n2276), .B1(ram[8658]), .B2(n2277), 
        .ZN(n12899) );
  MOAI22 U21813 ( .A1(n28466), .A2(n2276), .B1(ram[8659]), .B2(n2277), 
        .ZN(n12900) );
  MOAI22 U21814 ( .A1(n28231), .A2(n2276), .B1(ram[8660]), .B2(n2277), 
        .ZN(n12901) );
  MOAI22 U21815 ( .A1(n27996), .A2(n2276), .B1(ram[8661]), .B2(n2277), 
        .ZN(n12902) );
  MOAI22 U21816 ( .A1(n27761), .A2(n2276), .B1(ram[8662]), .B2(n2277), 
        .ZN(n12903) );
  MOAI22 U21817 ( .A1(n27526), .A2(n2276), .B1(ram[8663]), .B2(n2277), 
        .ZN(n12904) );
  MOAI22 U21818 ( .A1(n29171), .A2(n2278), .B1(ram[8664]), .B2(n2279), 
        .ZN(n12905) );
  MOAI22 U21819 ( .A1(n28936), .A2(n2278), .B1(ram[8665]), .B2(n2279), 
        .ZN(n12906) );
  MOAI22 U21820 ( .A1(n28701), .A2(n2278), .B1(ram[8666]), .B2(n2279), 
        .ZN(n12907) );
  MOAI22 U21821 ( .A1(n28466), .A2(n2278), .B1(ram[8667]), .B2(n2279), 
        .ZN(n12908) );
  MOAI22 U21822 ( .A1(n28231), .A2(n2278), .B1(ram[8668]), .B2(n2279), 
        .ZN(n12909) );
  MOAI22 U21823 ( .A1(n27996), .A2(n2278), .B1(ram[8669]), .B2(n2279), 
        .ZN(n12910) );
  MOAI22 U21824 ( .A1(n27761), .A2(n2278), .B1(ram[8670]), .B2(n2279), 
        .ZN(n12911) );
  MOAI22 U21825 ( .A1(n27526), .A2(n2278), .B1(ram[8671]), .B2(n2279), 
        .ZN(n12912) );
  MOAI22 U21826 ( .A1(n29171), .A2(n2280), .B1(ram[8672]), .B2(n2281), 
        .ZN(n12913) );
  MOAI22 U21827 ( .A1(n28936), .A2(n2280), .B1(ram[8673]), .B2(n2281), 
        .ZN(n12914) );
  MOAI22 U21828 ( .A1(n28701), .A2(n2280), .B1(ram[8674]), .B2(n2281), 
        .ZN(n12915) );
  MOAI22 U21829 ( .A1(n28466), .A2(n2280), .B1(ram[8675]), .B2(n2281), 
        .ZN(n12916) );
  MOAI22 U21830 ( .A1(n28231), .A2(n2280), .B1(ram[8676]), .B2(n2281), 
        .ZN(n12917) );
  MOAI22 U21831 ( .A1(n27996), .A2(n2280), .B1(ram[8677]), .B2(n2281), 
        .ZN(n12918) );
  MOAI22 U21832 ( .A1(n27761), .A2(n2280), .B1(ram[8678]), .B2(n2281), 
        .ZN(n12919) );
  MOAI22 U21833 ( .A1(n27526), .A2(n2280), .B1(ram[8679]), .B2(n2281), 
        .ZN(n12920) );
  MOAI22 U21834 ( .A1(n29171), .A2(n2282), .B1(ram[8680]), .B2(n2283), 
        .ZN(n12921) );
  MOAI22 U21835 ( .A1(n28936), .A2(n2282), .B1(ram[8681]), .B2(n2283), 
        .ZN(n12922) );
  MOAI22 U21836 ( .A1(n28701), .A2(n2282), .B1(ram[8682]), .B2(n2283), 
        .ZN(n12923) );
  MOAI22 U21837 ( .A1(n28466), .A2(n2282), .B1(ram[8683]), .B2(n2283), 
        .ZN(n12924) );
  MOAI22 U21838 ( .A1(n28231), .A2(n2282), .B1(ram[8684]), .B2(n2283), 
        .ZN(n12925) );
  MOAI22 U21839 ( .A1(n27996), .A2(n2282), .B1(ram[8685]), .B2(n2283), 
        .ZN(n12926) );
  MOAI22 U21840 ( .A1(n27761), .A2(n2282), .B1(ram[8686]), .B2(n2283), 
        .ZN(n12927) );
  MOAI22 U21841 ( .A1(n27526), .A2(n2282), .B1(ram[8687]), .B2(n2283), 
        .ZN(n12928) );
  MOAI22 U21842 ( .A1(n29171), .A2(n2284), .B1(ram[8688]), .B2(n2285), 
        .ZN(n12929) );
  MOAI22 U21843 ( .A1(n28936), .A2(n2284), .B1(ram[8689]), .B2(n2285), 
        .ZN(n12930) );
  MOAI22 U21844 ( .A1(n28701), .A2(n2284), .B1(ram[8690]), .B2(n2285), 
        .ZN(n12931) );
  MOAI22 U21845 ( .A1(n28466), .A2(n2284), .B1(ram[8691]), .B2(n2285), 
        .ZN(n12932) );
  MOAI22 U21846 ( .A1(n28231), .A2(n2284), .B1(ram[8692]), .B2(n2285), 
        .ZN(n12933) );
  MOAI22 U21847 ( .A1(n27996), .A2(n2284), .B1(ram[8693]), .B2(n2285), 
        .ZN(n12934) );
  MOAI22 U21848 ( .A1(n27761), .A2(n2284), .B1(ram[8694]), .B2(n2285), 
        .ZN(n12935) );
  MOAI22 U21849 ( .A1(n27526), .A2(n2284), .B1(ram[8695]), .B2(n2285), 
        .ZN(n12936) );
  MOAI22 U21850 ( .A1(n29171), .A2(n2286), .B1(ram[8696]), .B2(n2287), 
        .ZN(n12937) );
  MOAI22 U21851 ( .A1(n28936), .A2(n2286), .B1(ram[8697]), .B2(n2287), 
        .ZN(n12938) );
  MOAI22 U21852 ( .A1(n28701), .A2(n2286), .B1(ram[8698]), .B2(n2287), 
        .ZN(n12939) );
  MOAI22 U21853 ( .A1(n28466), .A2(n2286), .B1(ram[8699]), .B2(n2287), 
        .ZN(n12940) );
  MOAI22 U21854 ( .A1(n28231), .A2(n2286), .B1(ram[8700]), .B2(n2287), 
        .ZN(n12941) );
  MOAI22 U21855 ( .A1(n27996), .A2(n2286), .B1(ram[8701]), .B2(n2287), 
        .ZN(n12942) );
  MOAI22 U21856 ( .A1(n27761), .A2(n2286), .B1(ram[8702]), .B2(n2287), 
        .ZN(n12943) );
  MOAI22 U21857 ( .A1(n27526), .A2(n2286), .B1(ram[8703]), .B2(n2287), 
        .ZN(n12944) );
  MOAI22 U21858 ( .A1(n29171), .A2(n2289), .B1(ram[8704]), .B2(n2290), 
        .ZN(n12945) );
  MOAI22 U21859 ( .A1(n28936), .A2(n2289), .B1(ram[8705]), .B2(n2290), 
        .ZN(n12946) );
  MOAI22 U21860 ( .A1(n28701), .A2(n2289), .B1(ram[8706]), .B2(n2290), 
        .ZN(n12947) );
  MOAI22 U21861 ( .A1(n28466), .A2(n2289), .B1(ram[8707]), .B2(n2290), 
        .ZN(n12948) );
  MOAI22 U21862 ( .A1(n28231), .A2(n2289), .B1(ram[8708]), .B2(n2290), 
        .ZN(n12949) );
  MOAI22 U21863 ( .A1(n27996), .A2(n2289), .B1(ram[8709]), .B2(n2290), 
        .ZN(n12950) );
  MOAI22 U21864 ( .A1(n27761), .A2(n2289), .B1(ram[8710]), .B2(n2290), 
        .ZN(n12951) );
  MOAI22 U21865 ( .A1(n27526), .A2(n2289), .B1(ram[8711]), .B2(n2290), 
        .ZN(n12952) );
  MOAI22 U21866 ( .A1(n29171), .A2(n2292), .B1(ram[8712]), .B2(n2293), 
        .ZN(n12953) );
  MOAI22 U21867 ( .A1(n28936), .A2(n2292), .B1(ram[8713]), .B2(n2293), 
        .ZN(n12954) );
  MOAI22 U21868 ( .A1(n28701), .A2(n2292), .B1(ram[8714]), .B2(n2293), 
        .ZN(n12955) );
  MOAI22 U21869 ( .A1(n28466), .A2(n2292), .B1(ram[8715]), .B2(n2293), 
        .ZN(n12956) );
  MOAI22 U21870 ( .A1(n28231), .A2(n2292), .B1(ram[8716]), .B2(n2293), 
        .ZN(n12957) );
  MOAI22 U21871 ( .A1(n27996), .A2(n2292), .B1(ram[8717]), .B2(n2293), 
        .ZN(n12958) );
  MOAI22 U21872 ( .A1(n27761), .A2(n2292), .B1(ram[8718]), .B2(n2293), 
        .ZN(n12959) );
  MOAI22 U21873 ( .A1(n27526), .A2(n2292), .B1(ram[8719]), .B2(n2293), 
        .ZN(n12960) );
  MOAI22 U21874 ( .A1(n29171), .A2(n2294), .B1(ram[8720]), .B2(n2295), 
        .ZN(n12961) );
  MOAI22 U21875 ( .A1(n28936), .A2(n2294), .B1(ram[8721]), .B2(n2295), 
        .ZN(n12962) );
  MOAI22 U21876 ( .A1(n28701), .A2(n2294), .B1(ram[8722]), .B2(n2295), 
        .ZN(n12963) );
  MOAI22 U21877 ( .A1(n28466), .A2(n2294), .B1(ram[8723]), .B2(n2295), 
        .ZN(n12964) );
  MOAI22 U21878 ( .A1(n28231), .A2(n2294), .B1(ram[8724]), .B2(n2295), 
        .ZN(n12965) );
  MOAI22 U21879 ( .A1(n27996), .A2(n2294), .B1(ram[8725]), .B2(n2295), 
        .ZN(n12966) );
  MOAI22 U21880 ( .A1(n27761), .A2(n2294), .B1(ram[8726]), .B2(n2295), 
        .ZN(n12967) );
  MOAI22 U21881 ( .A1(n27526), .A2(n2294), .B1(ram[8727]), .B2(n2295), 
        .ZN(n12968) );
  MOAI22 U21882 ( .A1(n29171), .A2(n2296), .B1(ram[8728]), .B2(n2297), 
        .ZN(n12969) );
  MOAI22 U21883 ( .A1(n28936), .A2(n2296), .B1(ram[8729]), .B2(n2297), 
        .ZN(n12970) );
  MOAI22 U21884 ( .A1(n28701), .A2(n2296), .B1(ram[8730]), .B2(n2297), 
        .ZN(n12971) );
  MOAI22 U21885 ( .A1(n28466), .A2(n2296), .B1(ram[8731]), .B2(n2297), 
        .ZN(n12972) );
  MOAI22 U21886 ( .A1(n28231), .A2(n2296), .B1(ram[8732]), .B2(n2297), 
        .ZN(n12973) );
  MOAI22 U21887 ( .A1(n27996), .A2(n2296), .B1(ram[8733]), .B2(n2297), 
        .ZN(n12974) );
  MOAI22 U21888 ( .A1(n27761), .A2(n2296), .B1(ram[8734]), .B2(n2297), 
        .ZN(n12975) );
  MOAI22 U21889 ( .A1(n27526), .A2(n2296), .B1(ram[8735]), .B2(n2297), 
        .ZN(n12976) );
  MOAI22 U21890 ( .A1(n29172), .A2(n2298), .B1(ram[8736]), .B2(n2299), 
        .ZN(n12977) );
  MOAI22 U21891 ( .A1(n28937), .A2(n2298), .B1(ram[8737]), .B2(n2299), 
        .ZN(n12978) );
  MOAI22 U21892 ( .A1(n28702), .A2(n2298), .B1(ram[8738]), .B2(n2299), 
        .ZN(n12979) );
  MOAI22 U21893 ( .A1(n28467), .A2(n2298), .B1(ram[8739]), .B2(n2299), 
        .ZN(n12980) );
  MOAI22 U21894 ( .A1(n28232), .A2(n2298), .B1(ram[8740]), .B2(n2299), 
        .ZN(n12981) );
  MOAI22 U21895 ( .A1(n27997), .A2(n2298), .B1(ram[8741]), .B2(n2299), 
        .ZN(n12982) );
  MOAI22 U21896 ( .A1(n27762), .A2(n2298), .B1(ram[8742]), .B2(n2299), 
        .ZN(n12983) );
  MOAI22 U21897 ( .A1(n27527), .A2(n2298), .B1(ram[8743]), .B2(n2299), 
        .ZN(n12984) );
  MOAI22 U21898 ( .A1(n29172), .A2(n2300), .B1(ram[8744]), .B2(n2301), 
        .ZN(n12985) );
  MOAI22 U21899 ( .A1(n28937), .A2(n2300), .B1(ram[8745]), .B2(n2301), 
        .ZN(n12986) );
  MOAI22 U21900 ( .A1(n28702), .A2(n2300), .B1(ram[8746]), .B2(n2301), 
        .ZN(n12987) );
  MOAI22 U21901 ( .A1(n28467), .A2(n2300), .B1(ram[8747]), .B2(n2301), 
        .ZN(n12988) );
  MOAI22 U21902 ( .A1(n28232), .A2(n2300), .B1(ram[8748]), .B2(n2301), 
        .ZN(n12989) );
  MOAI22 U21903 ( .A1(n27997), .A2(n2300), .B1(ram[8749]), .B2(n2301), 
        .ZN(n12990) );
  MOAI22 U21904 ( .A1(n27762), .A2(n2300), .B1(ram[8750]), .B2(n2301), 
        .ZN(n12991) );
  MOAI22 U21905 ( .A1(n27527), .A2(n2300), .B1(ram[8751]), .B2(n2301), 
        .ZN(n12992) );
  MOAI22 U21906 ( .A1(n29172), .A2(n2302), .B1(ram[8752]), .B2(n2303), 
        .ZN(n12993) );
  MOAI22 U21907 ( .A1(n28937), .A2(n2302), .B1(ram[8753]), .B2(n2303), 
        .ZN(n12994) );
  MOAI22 U21908 ( .A1(n28702), .A2(n2302), .B1(ram[8754]), .B2(n2303), 
        .ZN(n12995) );
  MOAI22 U21909 ( .A1(n28467), .A2(n2302), .B1(ram[8755]), .B2(n2303), 
        .ZN(n12996) );
  MOAI22 U21910 ( .A1(n28232), .A2(n2302), .B1(ram[8756]), .B2(n2303), 
        .ZN(n12997) );
  MOAI22 U21911 ( .A1(n27997), .A2(n2302), .B1(ram[8757]), .B2(n2303), 
        .ZN(n12998) );
  MOAI22 U21912 ( .A1(n27762), .A2(n2302), .B1(ram[8758]), .B2(n2303), 
        .ZN(n12999) );
  MOAI22 U21913 ( .A1(n27527), .A2(n2302), .B1(ram[8759]), .B2(n2303), 
        .ZN(n13000) );
  MOAI22 U21914 ( .A1(n29172), .A2(n2304), .B1(ram[8760]), .B2(n2305), 
        .ZN(n13001) );
  MOAI22 U21915 ( .A1(n28937), .A2(n2304), .B1(ram[8761]), .B2(n2305), 
        .ZN(n13002) );
  MOAI22 U21916 ( .A1(n28702), .A2(n2304), .B1(ram[8762]), .B2(n2305), 
        .ZN(n13003) );
  MOAI22 U21917 ( .A1(n28467), .A2(n2304), .B1(ram[8763]), .B2(n2305), 
        .ZN(n13004) );
  MOAI22 U21918 ( .A1(n28232), .A2(n2304), .B1(ram[8764]), .B2(n2305), 
        .ZN(n13005) );
  MOAI22 U21919 ( .A1(n27997), .A2(n2304), .B1(ram[8765]), .B2(n2305), 
        .ZN(n13006) );
  MOAI22 U21920 ( .A1(n27762), .A2(n2304), .B1(ram[8766]), .B2(n2305), 
        .ZN(n13007) );
  MOAI22 U21921 ( .A1(n27527), .A2(n2304), .B1(ram[8767]), .B2(n2305), 
        .ZN(n13008) );
  MOAI22 U21922 ( .A1(n29172), .A2(n2306), .B1(ram[8768]), .B2(n2307), 
        .ZN(n13009) );
  MOAI22 U21923 ( .A1(n28937), .A2(n2306), .B1(ram[8769]), .B2(n2307), 
        .ZN(n13010) );
  MOAI22 U21924 ( .A1(n28702), .A2(n2306), .B1(ram[8770]), .B2(n2307), 
        .ZN(n13011) );
  MOAI22 U21925 ( .A1(n28467), .A2(n2306), .B1(ram[8771]), .B2(n2307), 
        .ZN(n13012) );
  MOAI22 U21926 ( .A1(n28232), .A2(n2306), .B1(ram[8772]), .B2(n2307), 
        .ZN(n13013) );
  MOAI22 U21927 ( .A1(n27997), .A2(n2306), .B1(ram[8773]), .B2(n2307), 
        .ZN(n13014) );
  MOAI22 U21928 ( .A1(n27762), .A2(n2306), .B1(ram[8774]), .B2(n2307), 
        .ZN(n13015) );
  MOAI22 U21929 ( .A1(n27527), .A2(n2306), .B1(ram[8775]), .B2(n2307), 
        .ZN(n13016) );
  MOAI22 U21930 ( .A1(n29172), .A2(n2308), .B1(ram[8776]), .B2(n2309), 
        .ZN(n13017) );
  MOAI22 U21931 ( .A1(n28937), .A2(n2308), .B1(ram[8777]), .B2(n2309), 
        .ZN(n13018) );
  MOAI22 U21932 ( .A1(n28702), .A2(n2308), .B1(ram[8778]), .B2(n2309), 
        .ZN(n13019) );
  MOAI22 U21933 ( .A1(n28467), .A2(n2308), .B1(ram[8779]), .B2(n2309), 
        .ZN(n13020) );
  MOAI22 U21934 ( .A1(n28232), .A2(n2308), .B1(ram[8780]), .B2(n2309), 
        .ZN(n13021) );
  MOAI22 U21935 ( .A1(n27997), .A2(n2308), .B1(ram[8781]), .B2(n2309), 
        .ZN(n13022) );
  MOAI22 U21936 ( .A1(n27762), .A2(n2308), .B1(ram[8782]), .B2(n2309), 
        .ZN(n13023) );
  MOAI22 U21937 ( .A1(n27527), .A2(n2308), .B1(ram[8783]), .B2(n2309), 
        .ZN(n13024) );
  MOAI22 U21938 ( .A1(n29172), .A2(n2310), .B1(ram[8784]), .B2(n2311), 
        .ZN(n13025) );
  MOAI22 U21939 ( .A1(n28937), .A2(n2310), .B1(ram[8785]), .B2(n2311), 
        .ZN(n13026) );
  MOAI22 U21940 ( .A1(n28702), .A2(n2310), .B1(ram[8786]), .B2(n2311), 
        .ZN(n13027) );
  MOAI22 U21941 ( .A1(n28467), .A2(n2310), .B1(ram[8787]), .B2(n2311), 
        .ZN(n13028) );
  MOAI22 U21942 ( .A1(n28232), .A2(n2310), .B1(ram[8788]), .B2(n2311), 
        .ZN(n13029) );
  MOAI22 U21943 ( .A1(n27997), .A2(n2310), .B1(ram[8789]), .B2(n2311), 
        .ZN(n13030) );
  MOAI22 U21944 ( .A1(n27762), .A2(n2310), .B1(ram[8790]), .B2(n2311), 
        .ZN(n13031) );
  MOAI22 U21945 ( .A1(n27527), .A2(n2310), .B1(ram[8791]), .B2(n2311), 
        .ZN(n13032) );
  MOAI22 U21946 ( .A1(n29172), .A2(n2312), .B1(ram[8792]), .B2(n2313), 
        .ZN(n13033) );
  MOAI22 U21947 ( .A1(n28937), .A2(n2312), .B1(ram[8793]), .B2(n2313), 
        .ZN(n13034) );
  MOAI22 U21948 ( .A1(n28702), .A2(n2312), .B1(ram[8794]), .B2(n2313), 
        .ZN(n13035) );
  MOAI22 U21949 ( .A1(n28467), .A2(n2312), .B1(ram[8795]), .B2(n2313), 
        .ZN(n13036) );
  MOAI22 U21950 ( .A1(n28232), .A2(n2312), .B1(ram[8796]), .B2(n2313), 
        .ZN(n13037) );
  MOAI22 U21951 ( .A1(n27997), .A2(n2312), .B1(ram[8797]), .B2(n2313), 
        .ZN(n13038) );
  MOAI22 U21952 ( .A1(n27762), .A2(n2312), .B1(ram[8798]), .B2(n2313), 
        .ZN(n13039) );
  MOAI22 U21953 ( .A1(n27527), .A2(n2312), .B1(ram[8799]), .B2(n2313), 
        .ZN(n13040) );
  MOAI22 U21954 ( .A1(n29172), .A2(n2314), .B1(ram[8800]), .B2(n2315), 
        .ZN(n13041) );
  MOAI22 U21955 ( .A1(n28937), .A2(n2314), .B1(ram[8801]), .B2(n2315), 
        .ZN(n13042) );
  MOAI22 U21956 ( .A1(n28702), .A2(n2314), .B1(ram[8802]), .B2(n2315), 
        .ZN(n13043) );
  MOAI22 U21957 ( .A1(n28467), .A2(n2314), .B1(ram[8803]), .B2(n2315), 
        .ZN(n13044) );
  MOAI22 U21958 ( .A1(n28232), .A2(n2314), .B1(ram[8804]), .B2(n2315), 
        .ZN(n13045) );
  MOAI22 U21959 ( .A1(n27997), .A2(n2314), .B1(ram[8805]), .B2(n2315), 
        .ZN(n13046) );
  MOAI22 U21960 ( .A1(n27762), .A2(n2314), .B1(ram[8806]), .B2(n2315), 
        .ZN(n13047) );
  MOAI22 U21961 ( .A1(n27527), .A2(n2314), .B1(ram[8807]), .B2(n2315), 
        .ZN(n13048) );
  MOAI22 U21962 ( .A1(n29172), .A2(n2316), .B1(ram[8808]), .B2(n2317), 
        .ZN(n13049) );
  MOAI22 U21963 ( .A1(n28937), .A2(n2316), .B1(ram[8809]), .B2(n2317), 
        .ZN(n13050) );
  MOAI22 U21964 ( .A1(n28702), .A2(n2316), .B1(ram[8810]), .B2(n2317), 
        .ZN(n13051) );
  MOAI22 U21965 ( .A1(n28467), .A2(n2316), .B1(ram[8811]), .B2(n2317), 
        .ZN(n13052) );
  MOAI22 U21966 ( .A1(n28232), .A2(n2316), .B1(ram[8812]), .B2(n2317), 
        .ZN(n13053) );
  MOAI22 U21967 ( .A1(n27997), .A2(n2316), .B1(ram[8813]), .B2(n2317), 
        .ZN(n13054) );
  MOAI22 U21968 ( .A1(n27762), .A2(n2316), .B1(ram[8814]), .B2(n2317), 
        .ZN(n13055) );
  MOAI22 U21969 ( .A1(n27527), .A2(n2316), .B1(ram[8815]), .B2(n2317), 
        .ZN(n13056) );
  MOAI22 U21970 ( .A1(n29172), .A2(n2318), .B1(ram[8816]), .B2(n2319), 
        .ZN(n13057) );
  MOAI22 U21971 ( .A1(n28937), .A2(n2318), .B1(ram[8817]), .B2(n2319), 
        .ZN(n13058) );
  MOAI22 U21972 ( .A1(n28702), .A2(n2318), .B1(ram[8818]), .B2(n2319), 
        .ZN(n13059) );
  MOAI22 U21973 ( .A1(n28467), .A2(n2318), .B1(ram[8819]), .B2(n2319), 
        .ZN(n13060) );
  MOAI22 U21974 ( .A1(n28232), .A2(n2318), .B1(ram[8820]), .B2(n2319), 
        .ZN(n13061) );
  MOAI22 U21975 ( .A1(n27997), .A2(n2318), .B1(ram[8821]), .B2(n2319), 
        .ZN(n13062) );
  MOAI22 U21976 ( .A1(n27762), .A2(n2318), .B1(ram[8822]), .B2(n2319), 
        .ZN(n13063) );
  MOAI22 U21977 ( .A1(n27527), .A2(n2318), .B1(ram[8823]), .B2(n2319), 
        .ZN(n13064) );
  MOAI22 U21978 ( .A1(n29172), .A2(n2320), .B1(ram[8824]), .B2(n2321), 
        .ZN(n13065) );
  MOAI22 U21979 ( .A1(n28937), .A2(n2320), .B1(ram[8825]), .B2(n2321), 
        .ZN(n13066) );
  MOAI22 U21980 ( .A1(n28702), .A2(n2320), .B1(ram[8826]), .B2(n2321), 
        .ZN(n13067) );
  MOAI22 U21981 ( .A1(n28467), .A2(n2320), .B1(ram[8827]), .B2(n2321), 
        .ZN(n13068) );
  MOAI22 U21982 ( .A1(n28232), .A2(n2320), .B1(ram[8828]), .B2(n2321), 
        .ZN(n13069) );
  MOAI22 U21983 ( .A1(n27997), .A2(n2320), .B1(ram[8829]), .B2(n2321), 
        .ZN(n13070) );
  MOAI22 U21984 ( .A1(n27762), .A2(n2320), .B1(ram[8830]), .B2(n2321), 
        .ZN(n13071) );
  MOAI22 U21985 ( .A1(n27527), .A2(n2320), .B1(ram[8831]), .B2(n2321), 
        .ZN(n13072) );
  MOAI22 U21986 ( .A1(n29172), .A2(n2322), .B1(ram[8832]), .B2(n2323), 
        .ZN(n13073) );
  MOAI22 U21987 ( .A1(n28937), .A2(n2322), .B1(ram[8833]), .B2(n2323), 
        .ZN(n13074) );
  MOAI22 U21988 ( .A1(n28702), .A2(n2322), .B1(ram[8834]), .B2(n2323), 
        .ZN(n13075) );
  MOAI22 U21989 ( .A1(n28467), .A2(n2322), .B1(ram[8835]), .B2(n2323), 
        .ZN(n13076) );
  MOAI22 U21990 ( .A1(n28232), .A2(n2322), .B1(ram[8836]), .B2(n2323), 
        .ZN(n13077) );
  MOAI22 U21991 ( .A1(n27997), .A2(n2322), .B1(ram[8837]), .B2(n2323), 
        .ZN(n13078) );
  MOAI22 U21992 ( .A1(n27762), .A2(n2322), .B1(ram[8838]), .B2(n2323), 
        .ZN(n13079) );
  MOAI22 U21993 ( .A1(n27527), .A2(n2322), .B1(ram[8839]), .B2(n2323), 
        .ZN(n13080) );
  MOAI22 U21994 ( .A1(n29173), .A2(n2324), .B1(ram[8840]), .B2(n2325), 
        .ZN(n13081) );
  MOAI22 U21995 ( .A1(n28938), .A2(n2324), .B1(ram[8841]), .B2(n2325), 
        .ZN(n13082) );
  MOAI22 U21996 ( .A1(n28703), .A2(n2324), .B1(ram[8842]), .B2(n2325), 
        .ZN(n13083) );
  MOAI22 U21997 ( .A1(n28468), .A2(n2324), .B1(ram[8843]), .B2(n2325), 
        .ZN(n13084) );
  MOAI22 U21998 ( .A1(n28233), .A2(n2324), .B1(ram[8844]), .B2(n2325), 
        .ZN(n13085) );
  MOAI22 U21999 ( .A1(n27998), .A2(n2324), .B1(ram[8845]), .B2(n2325), 
        .ZN(n13086) );
  MOAI22 U22000 ( .A1(n27763), .A2(n2324), .B1(ram[8846]), .B2(n2325), 
        .ZN(n13087) );
  MOAI22 U22001 ( .A1(n27528), .A2(n2324), .B1(ram[8847]), .B2(n2325), 
        .ZN(n13088) );
  MOAI22 U22002 ( .A1(n29173), .A2(n2326), .B1(ram[8848]), .B2(n2327), 
        .ZN(n13089) );
  MOAI22 U22003 ( .A1(n28938), .A2(n2326), .B1(ram[8849]), .B2(n2327), 
        .ZN(n13090) );
  MOAI22 U22004 ( .A1(n28703), .A2(n2326), .B1(ram[8850]), .B2(n2327), 
        .ZN(n13091) );
  MOAI22 U22005 ( .A1(n28468), .A2(n2326), .B1(ram[8851]), .B2(n2327), 
        .ZN(n13092) );
  MOAI22 U22006 ( .A1(n28233), .A2(n2326), .B1(ram[8852]), .B2(n2327), 
        .ZN(n13093) );
  MOAI22 U22007 ( .A1(n27998), .A2(n2326), .B1(ram[8853]), .B2(n2327), 
        .ZN(n13094) );
  MOAI22 U22008 ( .A1(n27763), .A2(n2326), .B1(ram[8854]), .B2(n2327), 
        .ZN(n13095) );
  MOAI22 U22009 ( .A1(n27528), .A2(n2326), .B1(ram[8855]), .B2(n2327), 
        .ZN(n13096) );
  MOAI22 U22010 ( .A1(n29173), .A2(n2328), .B1(ram[8856]), .B2(n2329), 
        .ZN(n13097) );
  MOAI22 U22011 ( .A1(n28938), .A2(n2328), .B1(ram[8857]), .B2(n2329), 
        .ZN(n13098) );
  MOAI22 U22012 ( .A1(n28703), .A2(n2328), .B1(ram[8858]), .B2(n2329), 
        .ZN(n13099) );
  MOAI22 U22013 ( .A1(n28468), .A2(n2328), .B1(ram[8859]), .B2(n2329), 
        .ZN(n13100) );
  MOAI22 U22014 ( .A1(n28233), .A2(n2328), .B1(ram[8860]), .B2(n2329), 
        .ZN(n13101) );
  MOAI22 U22015 ( .A1(n27998), .A2(n2328), .B1(ram[8861]), .B2(n2329), 
        .ZN(n13102) );
  MOAI22 U22016 ( .A1(n27763), .A2(n2328), .B1(ram[8862]), .B2(n2329), 
        .ZN(n13103) );
  MOAI22 U22017 ( .A1(n27528), .A2(n2328), .B1(ram[8863]), .B2(n2329), 
        .ZN(n13104) );
  MOAI22 U22018 ( .A1(n29173), .A2(n2330), .B1(ram[8864]), .B2(n2331), 
        .ZN(n13105) );
  MOAI22 U22019 ( .A1(n28938), .A2(n2330), .B1(ram[8865]), .B2(n2331), 
        .ZN(n13106) );
  MOAI22 U22020 ( .A1(n28703), .A2(n2330), .B1(ram[8866]), .B2(n2331), 
        .ZN(n13107) );
  MOAI22 U22021 ( .A1(n28468), .A2(n2330), .B1(ram[8867]), .B2(n2331), 
        .ZN(n13108) );
  MOAI22 U22022 ( .A1(n28233), .A2(n2330), .B1(ram[8868]), .B2(n2331), 
        .ZN(n13109) );
  MOAI22 U22023 ( .A1(n27998), .A2(n2330), .B1(ram[8869]), .B2(n2331), 
        .ZN(n13110) );
  MOAI22 U22024 ( .A1(n27763), .A2(n2330), .B1(ram[8870]), .B2(n2331), 
        .ZN(n13111) );
  MOAI22 U22025 ( .A1(n27528), .A2(n2330), .B1(ram[8871]), .B2(n2331), 
        .ZN(n13112) );
  MOAI22 U22026 ( .A1(n29173), .A2(n2332), .B1(ram[8872]), .B2(n2333), 
        .ZN(n13113) );
  MOAI22 U22027 ( .A1(n28938), .A2(n2332), .B1(ram[8873]), .B2(n2333), 
        .ZN(n13114) );
  MOAI22 U22028 ( .A1(n28703), .A2(n2332), .B1(ram[8874]), .B2(n2333), 
        .ZN(n13115) );
  MOAI22 U22029 ( .A1(n28468), .A2(n2332), .B1(ram[8875]), .B2(n2333), 
        .ZN(n13116) );
  MOAI22 U22030 ( .A1(n28233), .A2(n2332), .B1(ram[8876]), .B2(n2333), 
        .ZN(n13117) );
  MOAI22 U22031 ( .A1(n27998), .A2(n2332), .B1(ram[8877]), .B2(n2333), 
        .ZN(n13118) );
  MOAI22 U22032 ( .A1(n27763), .A2(n2332), .B1(ram[8878]), .B2(n2333), 
        .ZN(n13119) );
  MOAI22 U22033 ( .A1(n27528), .A2(n2332), .B1(ram[8879]), .B2(n2333), 
        .ZN(n13120) );
  MOAI22 U22034 ( .A1(n29173), .A2(n2334), .B1(ram[8880]), .B2(n2335), 
        .ZN(n13121) );
  MOAI22 U22035 ( .A1(n28938), .A2(n2334), .B1(ram[8881]), .B2(n2335), 
        .ZN(n13122) );
  MOAI22 U22036 ( .A1(n28703), .A2(n2334), .B1(ram[8882]), .B2(n2335), 
        .ZN(n13123) );
  MOAI22 U22037 ( .A1(n28468), .A2(n2334), .B1(ram[8883]), .B2(n2335), 
        .ZN(n13124) );
  MOAI22 U22038 ( .A1(n28233), .A2(n2334), .B1(ram[8884]), .B2(n2335), 
        .ZN(n13125) );
  MOAI22 U22039 ( .A1(n27998), .A2(n2334), .B1(ram[8885]), .B2(n2335), 
        .ZN(n13126) );
  MOAI22 U22040 ( .A1(n27763), .A2(n2334), .B1(ram[8886]), .B2(n2335), 
        .ZN(n13127) );
  MOAI22 U22041 ( .A1(n27528), .A2(n2334), .B1(ram[8887]), .B2(n2335), 
        .ZN(n13128) );
  MOAI22 U22042 ( .A1(n29173), .A2(n2336), .B1(ram[8888]), .B2(n2337), 
        .ZN(n13129) );
  MOAI22 U22043 ( .A1(n28938), .A2(n2336), .B1(ram[8889]), .B2(n2337), 
        .ZN(n13130) );
  MOAI22 U22044 ( .A1(n28703), .A2(n2336), .B1(ram[8890]), .B2(n2337), 
        .ZN(n13131) );
  MOAI22 U22045 ( .A1(n28468), .A2(n2336), .B1(ram[8891]), .B2(n2337), 
        .ZN(n13132) );
  MOAI22 U22046 ( .A1(n28233), .A2(n2336), .B1(ram[8892]), .B2(n2337), 
        .ZN(n13133) );
  MOAI22 U22047 ( .A1(n27998), .A2(n2336), .B1(ram[8893]), .B2(n2337), 
        .ZN(n13134) );
  MOAI22 U22048 ( .A1(n27763), .A2(n2336), .B1(ram[8894]), .B2(n2337), 
        .ZN(n13135) );
  MOAI22 U22049 ( .A1(n27528), .A2(n2336), .B1(ram[8895]), .B2(n2337), 
        .ZN(n13136) );
  MOAI22 U22050 ( .A1(n29173), .A2(n2338), .B1(ram[8896]), .B2(n2339), 
        .ZN(n13137) );
  MOAI22 U22051 ( .A1(n28938), .A2(n2338), .B1(ram[8897]), .B2(n2339), 
        .ZN(n13138) );
  MOAI22 U22052 ( .A1(n28703), .A2(n2338), .B1(ram[8898]), .B2(n2339), 
        .ZN(n13139) );
  MOAI22 U22053 ( .A1(n28468), .A2(n2338), .B1(ram[8899]), .B2(n2339), 
        .ZN(n13140) );
  MOAI22 U22054 ( .A1(n28233), .A2(n2338), .B1(ram[8900]), .B2(n2339), 
        .ZN(n13141) );
  MOAI22 U22055 ( .A1(n27998), .A2(n2338), .B1(ram[8901]), .B2(n2339), 
        .ZN(n13142) );
  MOAI22 U22056 ( .A1(n27763), .A2(n2338), .B1(ram[8902]), .B2(n2339), 
        .ZN(n13143) );
  MOAI22 U22057 ( .A1(n27528), .A2(n2338), .B1(ram[8903]), .B2(n2339), 
        .ZN(n13144) );
  MOAI22 U22058 ( .A1(n29173), .A2(n2340), .B1(ram[8904]), .B2(n2341), 
        .ZN(n13145) );
  MOAI22 U22059 ( .A1(n28938), .A2(n2340), .B1(ram[8905]), .B2(n2341), 
        .ZN(n13146) );
  MOAI22 U22060 ( .A1(n28703), .A2(n2340), .B1(ram[8906]), .B2(n2341), 
        .ZN(n13147) );
  MOAI22 U22061 ( .A1(n28468), .A2(n2340), .B1(ram[8907]), .B2(n2341), 
        .ZN(n13148) );
  MOAI22 U22062 ( .A1(n28233), .A2(n2340), .B1(ram[8908]), .B2(n2341), 
        .ZN(n13149) );
  MOAI22 U22063 ( .A1(n27998), .A2(n2340), .B1(ram[8909]), .B2(n2341), 
        .ZN(n13150) );
  MOAI22 U22064 ( .A1(n27763), .A2(n2340), .B1(ram[8910]), .B2(n2341), 
        .ZN(n13151) );
  MOAI22 U22065 ( .A1(n27528), .A2(n2340), .B1(ram[8911]), .B2(n2341), 
        .ZN(n13152) );
  MOAI22 U22066 ( .A1(n29173), .A2(n2342), .B1(ram[8912]), .B2(n2343), 
        .ZN(n13153) );
  MOAI22 U22067 ( .A1(n28938), .A2(n2342), .B1(ram[8913]), .B2(n2343), 
        .ZN(n13154) );
  MOAI22 U22068 ( .A1(n28703), .A2(n2342), .B1(ram[8914]), .B2(n2343), 
        .ZN(n13155) );
  MOAI22 U22069 ( .A1(n28468), .A2(n2342), .B1(ram[8915]), .B2(n2343), 
        .ZN(n13156) );
  MOAI22 U22070 ( .A1(n28233), .A2(n2342), .B1(ram[8916]), .B2(n2343), 
        .ZN(n13157) );
  MOAI22 U22071 ( .A1(n27998), .A2(n2342), .B1(ram[8917]), .B2(n2343), 
        .ZN(n13158) );
  MOAI22 U22072 ( .A1(n27763), .A2(n2342), .B1(ram[8918]), .B2(n2343), 
        .ZN(n13159) );
  MOAI22 U22073 ( .A1(n27528), .A2(n2342), .B1(ram[8919]), .B2(n2343), 
        .ZN(n13160) );
  MOAI22 U22074 ( .A1(n29173), .A2(n2344), .B1(ram[8920]), .B2(n2345), 
        .ZN(n13161) );
  MOAI22 U22075 ( .A1(n28938), .A2(n2344), .B1(ram[8921]), .B2(n2345), 
        .ZN(n13162) );
  MOAI22 U22076 ( .A1(n28703), .A2(n2344), .B1(ram[8922]), .B2(n2345), 
        .ZN(n13163) );
  MOAI22 U22077 ( .A1(n28468), .A2(n2344), .B1(ram[8923]), .B2(n2345), 
        .ZN(n13164) );
  MOAI22 U22078 ( .A1(n28233), .A2(n2344), .B1(ram[8924]), .B2(n2345), 
        .ZN(n13165) );
  MOAI22 U22079 ( .A1(n27998), .A2(n2344), .B1(ram[8925]), .B2(n2345), 
        .ZN(n13166) );
  MOAI22 U22080 ( .A1(n27763), .A2(n2344), .B1(ram[8926]), .B2(n2345), 
        .ZN(n13167) );
  MOAI22 U22081 ( .A1(n27528), .A2(n2344), .B1(ram[8927]), .B2(n2345), 
        .ZN(n13168) );
  MOAI22 U22082 ( .A1(n29173), .A2(n2346), .B1(ram[8928]), .B2(n2347), 
        .ZN(n13169) );
  MOAI22 U22083 ( .A1(n28938), .A2(n2346), .B1(ram[8929]), .B2(n2347), 
        .ZN(n13170) );
  MOAI22 U22084 ( .A1(n28703), .A2(n2346), .B1(ram[8930]), .B2(n2347), 
        .ZN(n13171) );
  MOAI22 U22085 ( .A1(n28468), .A2(n2346), .B1(ram[8931]), .B2(n2347), 
        .ZN(n13172) );
  MOAI22 U22086 ( .A1(n28233), .A2(n2346), .B1(ram[8932]), .B2(n2347), 
        .ZN(n13173) );
  MOAI22 U22087 ( .A1(n27998), .A2(n2346), .B1(ram[8933]), .B2(n2347), 
        .ZN(n13174) );
  MOAI22 U22088 ( .A1(n27763), .A2(n2346), .B1(ram[8934]), .B2(n2347), 
        .ZN(n13175) );
  MOAI22 U22089 ( .A1(n27528), .A2(n2346), .B1(ram[8935]), .B2(n2347), 
        .ZN(n13176) );
  MOAI22 U22090 ( .A1(n29173), .A2(n2348), .B1(ram[8936]), .B2(n2349), 
        .ZN(n13177) );
  MOAI22 U22091 ( .A1(n28938), .A2(n2348), .B1(ram[8937]), .B2(n2349), 
        .ZN(n13178) );
  MOAI22 U22092 ( .A1(n28703), .A2(n2348), .B1(ram[8938]), .B2(n2349), 
        .ZN(n13179) );
  MOAI22 U22093 ( .A1(n28468), .A2(n2348), .B1(ram[8939]), .B2(n2349), 
        .ZN(n13180) );
  MOAI22 U22094 ( .A1(n28233), .A2(n2348), .B1(ram[8940]), .B2(n2349), 
        .ZN(n13181) );
  MOAI22 U22095 ( .A1(n27998), .A2(n2348), .B1(ram[8941]), .B2(n2349), 
        .ZN(n13182) );
  MOAI22 U22096 ( .A1(n27763), .A2(n2348), .B1(ram[8942]), .B2(n2349), 
        .ZN(n13183) );
  MOAI22 U22097 ( .A1(n27528), .A2(n2348), .B1(ram[8943]), .B2(n2349), 
        .ZN(n13184) );
  MOAI22 U22098 ( .A1(n29174), .A2(n2350), .B1(ram[8944]), .B2(n2351), 
        .ZN(n13185) );
  MOAI22 U22099 ( .A1(n28939), .A2(n2350), .B1(ram[8945]), .B2(n2351), 
        .ZN(n13186) );
  MOAI22 U22100 ( .A1(n28704), .A2(n2350), .B1(ram[8946]), .B2(n2351), 
        .ZN(n13187) );
  MOAI22 U22101 ( .A1(n28469), .A2(n2350), .B1(ram[8947]), .B2(n2351), 
        .ZN(n13188) );
  MOAI22 U22102 ( .A1(n28234), .A2(n2350), .B1(ram[8948]), .B2(n2351), 
        .ZN(n13189) );
  MOAI22 U22103 ( .A1(n27999), .A2(n2350), .B1(ram[8949]), .B2(n2351), 
        .ZN(n13190) );
  MOAI22 U22104 ( .A1(n27764), .A2(n2350), .B1(ram[8950]), .B2(n2351), 
        .ZN(n13191) );
  MOAI22 U22105 ( .A1(n27529), .A2(n2350), .B1(ram[8951]), .B2(n2351), 
        .ZN(n13192) );
  MOAI22 U22106 ( .A1(n29174), .A2(n2352), .B1(ram[8952]), .B2(n2353), 
        .ZN(n13193) );
  MOAI22 U22107 ( .A1(n28939), .A2(n2352), .B1(ram[8953]), .B2(n2353), 
        .ZN(n13194) );
  MOAI22 U22108 ( .A1(n28704), .A2(n2352), .B1(ram[8954]), .B2(n2353), 
        .ZN(n13195) );
  MOAI22 U22109 ( .A1(n28469), .A2(n2352), .B1(ram[8955]), .B2(n2353), 
        .ZN(n13196) );
  MOAI22 U22110 ( .A1(n28234), .A2(n2352), .B1(ram[8956]), .B2(n2353), 
        .ZN(n13197) );
  MOAI22 U22111 ( .A1(n27999), .A2(n2352), .B1(ram[8957]), .B2(n2353), 
        .ZN(n13198) );
  MOAI22 U22112 ( .A1(n27764), .A2(n2352), .B1(ram[8958]), .B2(n2353), 
        .ZN(n13199) );
  MOAI22 U22113 ( .A1(n27529), .A2(n2352), .B1(ram[8959]), .B2(n2353), 
        .ZN(n13200) );
  MOAI22 U22114 ( .A1(n29174), .A2(n2354), .B1(ram[8960]), .B2(n2355), 
        .ZN(n13201) );
  MOAI22 U22115 ( .A1(n28939), .A2(n2354), .B1(ram[8961]), .B2(n2355), 
        .ZN(n13202) );
  MOAI22 U22116 ( .A1(n28704), .A2(n2354), .B1(ram[8962]), .B2(n2355), 
        .ZN(n13203) );
  MOAI22 U22117 ( .A1(n28469), .A2(n2354), .B1(ram[8963]), .B2(n2355), 
        .ZN(n13204) );
  MOAI22 U22118 ( .A1(n28234), .A2(n2354), .B1(ram[8964]), .B2(n2355), 
        .ZN(n13205) );
  MOAI22 U22119 ( .A1(n27999), .A2(n2354), .B1(ram[8965]), .B2(n2355), 
        .ZN(n13206) );
  MOAI22 U22120 ( .A1(n27764), .A2(n2354), .B1(ram[8966]), .B2(n2355), 
        .ZN(n13207) );
  MOAI22 U22121 ( .A1(n27529), .A2(n2354), .B1(ram[8967]), .B2(n2355), 
        .ZN(n13208) );
  MOAI22 U22122 ( .A1(n29174), .A2(n2356), .B1(ram[8968]), .B2(n2357), 
        .ZN(n13209) );
  MOAI22 U22123 ( .A1(n28939), .A2(n2356), .B1(ram[8969]), .B2(n2357), 
        .ZN(n13210) );
  MOAI22 U22124 ( .A1(n28704), .A2(n2356), .B1(ram[8970]), .B2(n2357), 
        .ZN(n13211) );
  MOAI22 U22125 ( .A1(n28469), .A2(n2356), .B1(ram[8971]), .B2(n2357), 
        .ZN(n13212) );
  MOAI22 U22126 ( .A1(n28234), .A2(n2356), .B1(ram[8972]), .B2(n2357), 
        .ZN(n13213) );
  MOAI22 U22127 ( .A1(n27999), .A2(n2356), .B1(ram[8973]), .B2(n2357), 
        .ZN(n13214) );
  MOAI22 U22128 ( .A1(n27764), .A2(n2356), .B1(ram[8974]), .B2(n2357), 
        .ZN(n13215) );
  MOAI22 U22129 ( .A1(n27529), .A2(n2356), .B1(ram[8975]), .B2(n2357), 
        .ZN(n13216) );
  MOAI22 U22130 ( .A1(n29174), .A2(n2358), .B1(ram[8976]), .B2(n2359), 
        .ZN(n13217) );
  MOAI22 U22131 ( .A1(n28939), .A2(n2358), .B1(ram[8977]), .B2(n2359), 
        .ZN(n13218) );
  MOAI22 U22132 ( .A1(n28704), .A2(n2358), .B1(ram[8978]), .B2(n2359), 
        .ZN(n13219) );
  MOAI22 U22133 ( .A1(n28469), .A2(n2358), .B1(ram[8979]), .B2(n2359), 
        .ZN(n13220) );
  MOAI22 U22134 ( .A1(n28234), .A2(n2358), .B1(ram[8980]), .B2(n2359), 
        .ZN(n13221) );
  MOAI22 U22135 ( .A1(n27999), .A2(n2358), .B1(ram[8981]), .B2(n2359), 
        .ZN(n13222) );
  MOAI22 U22136 ( .A1(n27764), .A2(n2358), .B1(ram[8982]), .B2(n2359), 
        .ZN(n13223) );
  MOAI22 U22137 ( .A1(n27529), .A2(n2358), .B1(ram[8983]), .B2(n2359), 
        .ZN(n13224) );
  MOAI22 U22138 ( .A1(n29174), .A2(n2360), .B1(ram[8984]), .B2(n2361), 
        .ZN(n13225) );
  MOAI22 U22139 ( .A1(n28939), .A2(n2360), .B1(ram[8985]), .B2(n2361), 
        .ZN(n13226) );
  MOAI22 U22140 ( .A1(n28704), .A2(n2360), .B1(ram[8986]), .B2(n2361), 
        .ZN(n13227) );
  MOAI22 U22141 ( .A1(n28469), .A2(n2360), .B1(ram[8987]), .B2(n2361), 
        .ZN(n13228) );
  MOAI22 U22142 ( .A1(n28234), .A2(n2360), .B1(ram[8988]), .B2(n2361), 
        .ZN(n13229) );
  MOAI22 U22143 ( .A1(n27999), .A2(n2360), .B1(ram[8989]), .B2(n2361), 
        .ZN(n13230) );
  MOAI22 U22144 ( .A1(n27764), .A2(n2360), .B1(ram[8990]), .B2(n2361), 
        .ZN(n13231) );
  MOAI22 U22145 ( .A1(n27529), .A2(n2360), .B1(ram[8991]), .B2(n2361), 
        .ZN(n13232) );
  MOAI22 U22146 ( .A1(n29174), .A2(n2362), .B1(ram[8992]), .B2(n2363), 
        .ZN(n13233) );
  MOAI22 U22147 ( .A1(n28939), .A2(n2362), .B1(ram[8993]), .B2(n2363), 
        .ZN(n13234) );
  MOAI22 U22148 ( .A1(n28704), .A2(n2362), .B1(ram[8994]), .B2(n2363), 
        .ZN(n13235) );
  MOAI22 U22149 ( .A1(n28469), .A2(n2362), .B1(ram[8995]), .B2(n2363), 
        .ZN(n13236) );
  MOAI22 U22150 ( .A1(n28234), .A2(n2362), .B1(ram[8996]), .B2(n2363), 
        .ZN(n13237) );
  MOAI22 U22151 ( .A1(n27999), .A2(n2362), .B1(ram[8997]), .B2(n2363), 
        .ZN(n13238) );
  MOAI22 U22152 ( .A1(n27764), .A2(n2362), .B1(ram[8998]), .B2(n2363), 
        .ZN(n13239) );
  MOAI22 U22153 ( .A1(n27529), .A2(n2362), .B1(ram[8999]), .B2(n2363), 
        .ZN(n13240) );
  MOAI22 U22154 ( .A1(n29174), .A2(n2364), .B1(ram[9000]), .B2(n2365), 
        .ZN(n13241) );
  MOAI22 U22155 ( .A1(n28939), .A2(n2364), .B1(ram[9001]), .B2(n2365), 
        .ZN(n13242) );
  MOAI22 U22156 ( .A1(n28704), .A2(n2364), .B1(ram[9002]), .B2(n2365), 
        .ZN(n13243) );
  MOAI22 U22157 ( .A1(n28469), .A2(n2364), .B1(ram[9003]), .B2(n2365), 
        .ZN(n13244) );
  MOAI22 U22158 ( .A1(n28234), .A2(n2364), .B1(ram[9004]), .B2(n2365), 
        .ZN(n13245) );
  MOAI22 U22159 ( .A1(n27999), .A2(n2364), .B1(ram[9005]), .B2(n2365), 
        .ZN(n13246) );
  MOAI22 U22160 ( .A1(n27764), .A2(n2364), .B1(ram[9006]), .B2(n2365), 
        .ZN(n13247) );
  MOAI22 U22161 ( .A1(n27529), .A2(n2364), .B1(ram[9007]), .B2(n2365), 
        .ZN(n13248) );
  MOAI22 U22162 ( .A1(n29174), .A2(n2366), .B1(ram[9008]), .B2(n2367), 
        .ZN(n13249) );
  MOAI22 U22163 ( .A1(n28939), .A2(n2366), .B1(ram[9009]), .B2(n2367), 
        .ZN(n13250) );
  MOAI22 U22164 ( .A1(n28704), .A2(n2366), .B1(ram[9010]), .B2(n2367), 
        .ZN(n13251) );
  MOAI22 U22165 ( .A1(n28469), .A2(n2366), .B1(ram[9011]), .B2(n2367), 
        .ZN(n13252) );
  MOAI22 U22166 ( .A1(n28234), .A2(n2366), .B1(ram[9012]), .B2(n2367), 
        .ZN(n13253) );
  MOAI22 U22167 ( .A1(n27999), .A2(n2366), .B1(ram[9013]), .B2(n2367), 
        .ZN(n13254) );
  MOAI22 U22168 ( .A1(n27764), .A2(n2366), .B1(ram[9014]), .B2(n2367), 
        .ZN(n13255) );
  MOAI22 U22169 ( .A1(n27529), .A2(n2366), .B1(ram[9015]), .B2(n2367), 
        .ZN(n13256) );
  MOAI22 U22170 ( .A1(n29174), .A2(n2368), .B1(ram[9016]), .B2(n2369), 
        .ZN(n13257) );
  MOAI22 U22171 ( .A1(n28939), .A2(n2368), .B1(ram[9017]), .B2(n2369), 
        .ZN(n13258) );
  MOAI22 U22172 ( .A1(n28704), .A2(n2368), .B1(ram[9018]), .B2(n2369), 
        .ZN(n13259) );
  MOAI22 U22173 ( .A1(n28469), .A2(n2368), .B1(ram[9019]), .B2(n2369), 
        .ZN(n13260) );
  MOAI22 U22174 ( .A1(n28234), .A2(n2368), .B1(ram[9020]), .B2(n2369), 
        .ZN(n13261) );
  MOAI22 U22175 ( .A1(n27999), .A2(n2368), .B1(ram[9021]), .B2(n2369), 
        .ZN(n13262) );
  MOAI22 U22176 ( .A1(n27764), .A2(n2368), .B1(ram[9022]), .B2(n2369), 
        .ZN(n13263) );
  MOAI22 U22177 ( .A1(n27529), .A2(n2368), .B1(ram[9023]), .B2(n2369), 
        .ZN(n13264) );
  MOAI22 U22178 ( .A1(n29174), .A2(n2370), .B1(ram[9024]), .B2(n2371), 
        .ZN(n13265) );
  MOAI22 U22179 ( .A1(n28939), .A2(n2370), .B1(ram[9025]), .B2(n2371), 
        .ZN(n13266) );
  MOAI22 U22180 ( .A1(n28704), .A2(n2370), .B1(ram[9026]), .B2(n2371), 
        .ZN(n13267) );
  MOAI22 U22181 ( .A1(n28469), .A2(n2370), .B1(ram[9027]), .B2(n2371), 
        .ZN(n13268) );
  MOAI22 U22182 ( .A1(n28234), .A2(n2370), .B1(ram[9028]), .B2(n2371), 
        .ZN(n13269) );
  MOAI22 U22183 ( .A1(n27999), .A2(n2370), .B1(ram[9029]), .B2(n2371), 
        .ZN(n13270) );
  MOAI22 U22184 ( .A1(n27764), .A2(n2370), .B1(ram[9030]), .B2(n2371), 
        .ZN(n13271) );
  MOAI22 U22185 ( .A1(n27529), .A2(n2370), .B1(ram[9031]), .B2(n2371), 
        .ZN(n13272) );
  MOAI22 U22186 ( .A1(n29174), .A2(n2372), .B1(ram[9032]), .B2(n2373), 
        .ZN(n13273) );
  MOAI22 U22187 ( .A1(n28939), .A2(n2372), .B1(ram[9033]), .B2(n2373), 
        .ZN(n13274) );
  MOAI22 U22188 ( .A1(n28704), .A2(n2372), .B1(ram[9034]), .B2(n2373), 
        .ZN(n13275) );
  MOAI22 U22189 ( .A1(n28469), .A2(n2372), .B1(ram[9035]), .B2(n2373), 
        .ZN(n13276) );
  MOAI22 U22190 ( .A1(n28234), .A2(n2372), .B1(ram[9036]), .B2(n2373), 
        .ZN(n13277) );
  MOAI22 U22191 ( .A1(n27999), .A2(n2372), .B1(ram[9037]), .B2(n2373), 
        .ZN(n13278) );
  MOAI22 U22192 ( .A1(n27764), .A2(n2372), .B1(ram[9038]), .B2(n2373), 
        .ZN(n13279) );
  MOAI22 U22193 ( .A1(n27529), .A2(n2372), .B1(ram[9039]), .B2(n2373), 
        .ZN(n13280) );
  MOAI22 U22194 ( .A1(n29174), .A2(n2374), .B1(ram[9040]), .B2(n2375), 
        .ZN(n13281) );
  MOAI22 U22195 ( .A1(n28939), .A2(n2374), .B1(ram[9041]), .B2(n2375), 
        .ZN(n13282) );
  MOAI22 U22196 ( .A1(n28704), .A2(n2374), .B1(ram[9042]), .B2(n2375), 
        .ZN(n13283) );
  MOAI22 U22197 ( .A1(n28469), .A2(n2374), .B1(ram[9043]), .B2(n2375), 
        .ZN(n13284) );
  MOAI22 U22198 ( .A1(n28234), .A2(n2374), .B1(ram[9044]), .B2(n2375), 
        .ZN(n13285) );
  MOAI22 U22199 ( .A1(n27999), .A2(n2374), .B1(ram[9045]), .B2(n2375), 
        .ZN(n13286) );
  MOAI22 U22200 ( .A1(n27764), .A2(n2374), .B1(ram[9046]), .B2(n2375), 
        .ZN(n13287) );
  MOAI22 U22201 ( .A1(n27529), .A2(n2374), .B1(ram[9047]), .B2(n2375), 
        .ZN(n13288) );
  MOAI22 U22202 ( .A1(n29175), .A2(n2376), .B1(ram[9048]), .B2(n2377), 
        .ZN(n13289) );
  MOAI22 U22203 ( .A1(n28940), .A2(n2376), .B1(ram[9049]), .B2(n2377), 
        .ZN(n13290) );
  MOAI22 U22204 ( .A1(n28705), .A2(n2376), .B1(ram[9050]), .B2(n2377), 
        .ZN(n13291) );
  MOAI22 U22205 ( .A1(n28470), .A2(n2376), .B1(ram[9051]), .B2(n2377), 
        .ZN(n13292) );
  MOAI22 U22206 ( .A1(n28235), .A2(n2376), .B1(ram[9052]), .B2(n2377), 
        .ZN(n13293) );
  MOAI22 U22207 ( .A1(n28000), .A2(n2376), .B1(ram[9053]), .B2(n2377), 
        .ZN(n13294) );
  MOAI22 U22208 ( .A1(n27765), .A2(n2376), .B1(ram[9054]), .B2(n2377), 
        .ZN(n13295) );
  MOAI22 U22209 ( .A1(n27530), .A2(n2376), .B1(ram[9055]), .B2(n2377), 
        .ZN(n13296) );
  MOAI22 U22210 ( .A1(n29175), .A2(n2378), .B1(ram[9056]), .B2(n2379), 
        .ZN(n13297) );
  MOAI22 U22211 ( .A1(n28940), .A2(n2378), .B1(ram[9057]), .B2(n2379), 
        .ZN(n13298) );
  MOAI22 U22212 ( .A1(n28705), .A2(n2378), .B1(ram[9058]), .B2(n2379), 
        .ZN(n13299) );
  MOAI22 U22213 ( .A1(n28470), .A2(n2378), .B1(ram[9059]), .B2(n2379), 
        .ZN(n13300) );
  MOAI22 U22214 ( .A1(n28235), .A2(n2378), .B1(ram[9060]), .B2(n2379), 
        .ZN(n13301) );
  MOAI22 U22215 ( .A1(n28000), .A2(n2378), .B1(ram[9061]), .B2(n2379), 
        .ZN(n13302) );
  MOAI22 U22216 ( .A1(n27765), .A2(n2378), .B1(ram[9062]), .B2(n2379), 
        .ZN(n13303) );
  MOAI22 U22217 ( .A1(n27530), .A2(n2378), .B1(ram[9063]), .B2(n2379), 
        .ZN(n13304) );
  MOAI22 U22218 ( .A1(n29175), .A2(n2380), .B1(ram[9064]), .B2(n2381), 
        .ZN(n13305) );
  MOAI22 U22219 ( .A1(n28940), .A2(n2380), .B1(ram[9065]), .B2(n2381), 
        .ZN(n13306) );
  MOAI22 U22220 ( .A1(n28705), .A2(n2380), .B1(ram[9066]), .B2(n2381), 
        .ZN(n13307) );
  MOAI22 U22221 ( .A1(n28470), .A2(n2380), .B1(ram[9067]), .B2(n2381), 
        .ZN(n13308) );
  MOAI22 U22222 ( .A1(n28235), .A2(n2380), .B1(ram[9068]), .B2(n2381), 
        .ZN(n13309) );
  MOAI22 U22223 ( .A1(n28000), .A2(n2380), .B1(ram[9069]), .B2(n2381), 
        .ZN(n13310) );
  MOAI22 U22224 ( .A1(n27765), .A2(n2380), .B1(ram[9070]), .B2(n2381), 
        .ZN(n13311) );
  MOAI22 U22225 ( .A1(n27530), .A2(n2380), .B1(ram[9071]), .B2(n2381), 
        .ZN(n13312) );
  MOAI22 U22226 ( .A1(n29175), .A2(n2382), .B1(ram[9072]), .B2(n2383), 
        .ZN(n13313) );
  MOAI22 U22227 ( .A1(n28940), .A2(n2382), .B1(ram[9073]), .B2(n2383), 
        .ZN(n13314) );
  MOAI22 U22228 ( .A1(n28705), .A2(n2382), .B1(ram[9074]), .B2(n2383), 
        .ZN(n13315) );
  MOAI22 U22229 ( .A1(n28470), .A2(n2382), .B1(ram[9075]), .B2(n2383), 
        .ZN(n13316) );
  MOAI22 U22230 ( .A1(n28235), .A2(n2382), .B1(ram[9076]), .B2(n2383), 
        .ZN(n13317) );
  MOAI22 U22231 ( .A1(n28000), .A2(n2382), .B1(ram[9077]), .B2(n2383), 
        .ZN(n13318) );
  MOAI22 U22232 ( .A1(n27765), .A2(n2382), .B1(ram[9078]), .B2(n2383), 
        .ZN(n13319) );
  MOAI22 U22233 ( .A1(n27530), .A2(n2382), .B1(ram[9079]), .B2(n2383), 
        .ZN(n13320) );
  MOAI22 U22234 ( .A1(n29175), .A2(n2384), .B1(ram[9080]), .B2(n2385), 
        .ZN(n13321) );
  MOAI22 U22235 ( .A1(n28940), .A2(n2384), .B1(ram[9081]), .B2(n2385), 
        .ZN(n13322) );
  MOAI22 U22236 ( .A1(n28705), .A2(n2384), .B1(ram[9082]), .B2(n2385), 
        .ZN(n13323) );
  MOAI22 U22237 ( .A1(n28470), .A2(n2384), .B1(ram[9083]), .B2(n2385), 
        .ZN(n13324) );
  MOAI22 U22238 ( .A1(n28235), .A2(n2384), .B1(ram[9084]), .B2(n2385), 
        .ZN(n13325) );
  MOAI22 U22239 ( .A1(n28000), .A2(n2384), .B1(ram[9085]), .B2(n2385), 
        .ZN(n13326) );
  MOAI22 U22240 ( .A1(n27765), .A2(n2384), .B1(ram[9086]), .B2(n2385), 
        .ZN(n13327) );
  MOAI22 U22241 ( .A1(n27530), .A2(n2384), .B1(ram[9087]), .B2(n2385), 
        .ZN(n13328) );
  MOAI22 U22242 ( .A1(n29175), .A2(n2386), .B1(ram[9088]), .B2(n2387), 
        .ZN(n13329) );
  MOAI22 U22243 ( .A1(n28940), .A2(n2386), .B1(ram[9089]), .B2(n2387), 
        .ZN(n13330) );
  MOAI22 U22244 ( .A1(n28705), .A2(n2386), .B1(ram[9090]), .B2(n2387), 
        .ZN(n13331) );
  MOAI22 U22245 ( .A1(n28470), .A2(n2386), .B1(ram[9091]), .B2(n2387), 
        .ZN(n13332) );
  MOAI22 U22246 ( .A1(n28235), .A2(n2386), .B1(ram[9092]), .B2(n2387), 
        .ZN(n13333) );
  MOAI22 U22247 ( .A1(n28000), .A2(n2386), .B1(ram[9093]), .B2(n2387), 
        .ZN(n13334) );
  MOAI22 U22248 ( .A1(n27765), .A2(n2386), .B1(ram[9094]), .B2(n2387), 
        .ZN(n13335) );
  MOAI22 U22249 ( .A1(n27530), .A2(n2386), .B1(ram[9095]), .B2(n2387), 
        .ZN(n13336) );
  MOAI22 U22250 ( .A1(n29175), .A2(n2388), .B1(ram[9096]), .B2(n2389), 
        .ZN(n13337) );
  MOAI22 U22251 ( .A1(n28940), .A2(n2388), .B1(ram[9097]), .B2(n2389), 
        .ZN(n13338) );
  MOAI22 U22252 ( .A1(n28705), .A2(n2388), .B1(ram[9098]), .B2(n2389), 
        .ZN(n13339) );
  MOAI22 U22253 ( .A1(n28470), .A2(n2388), .B1(ram[9099]), .B2(n2389), 
        .ZN(n13340) );
  MOAI22 U22254 ( .A1(n28235), .A2(n2388), .B1(ram[9100]), .B2(n2389), 
        .ZN(n13341) );
  MOAI22 U22255 ( .A1(n28000), .A2(n2388), .B1(ram[9101]), .B2(n2389), 
        .ZN(n13342) );
  MOAI22 U22256 ( .A1(n27765), .A2(n2388), .B1(ram[9102]), .B2(n2389), 
        .ZN(n13343) );
  MOAI22 U22257 ( .A1(n27530), .A2(n2388), .B1(ram[9103]), .B2(n2389), 
        .ZN(n13344) );
  MOAI22 U22258 ( .A1(n29175), .A2(n2390), .B1(ram[9104]), .B2(n2391), 
        .ZN(n13345) );
  MOAI22 U22259 ( .A1(n28940), .A2(n2390), .B1(ram[9105]), .B2(n2391), 
        .ZN(n13346) );
  MOAI22 U22260 ( .A1(n28705), .A2(n2390), .B1(ram[9106]), .B2(n2391), 
        .ZN(n13347) );
  MOAI22 U22261 ( .A1(n28470), .A2(n2390), .B1(ram[9107]), .B2(n2391), 
        .ZN(n13348) );
  MOAI22 U22262 ( .A1(n28235), .A2(n2390), .B1(ram[9108]), .B2(n2391), 
        .ZN(n13349) );
  MOAI22 U22263 ( .A1(n28000), .A2(n2390), .B1(ram[9109]), .B2(n2391), 
        .ZN(n13350) );
  MOAI22 U22264 ( .A1(n27765), .A2(n2390), .B1(ram[9110]), .B2(n2391), 
        .ZN(n13351) );
  MOAI22 U22265 ( .A1(n27530), .A2(n2390), .B1(ram[9111]), .B2(n2391), 
        .ZN(n13352) );
  MOAI22 U22266 ( .A1(n29175), .A2(n2392), .B1(ram[9112]), .B2(n2393), 
        .ZN(n13353) );
  MOAI22 U22267 ( .A1(n28940), .A2(n2392), .B1(ram[9113]), .B2(n2393), 
        .ZN(n13354) );
  MOAI22 U22268 ( .A1(n28705), .A2(n2392), .B1(ram[9114]), .B2(n2393), 
        .ZN(n13355) );
  MOAI22 U22269 ( .A1(n28470), .A2(n2392), .B1(ram[9115]), .B2(n2393), 
        .ZN(n13356) );
  MOAI22 U22270 ( .A1(n28235), .A2(n2392), .B1(ram[9116]), .B2(n2393), 
        .ZN(n13357) );
  MOAI22 U22271 ( .A1(n28000), .A2(n2392), .B1(ram[9117]), .B2(n2393), 
        .ZN(n13358) );
  MOAI22 U22272 ( .A1(n27765), .A2(n2392), .B1(ram[9118]), .B2(n2393), 
        .ZN(n13359) );
  MOAI22 U22273 ( .A1(n27530), .A2(n2392), .B1(ram[9119]), .B2(n2393), 
        .ZN(n13360) );
  MOAI22 U22274 ( .A1(n29175), .A2(n2394), .B1(ram[9120]), .B2(n2395), 
        .ZN(n13361) );
  MOAI22 U22275 ( .A1(n28940), .A2(n2394), .B1(ram[9121]), .B2(n2395), 
        .ZN(n13362) );
  MOAI22 U22276 ( .A1(n28705), .A2(n2394), .B1(ram[9122]), .B2(n2395), 
        .ZN(n13363) );
  MOAI22 U22277 ( .A1(n28470), .A2(n2394), .B1(ram[9123]), .B2(n2395), 
        .ZN(n13364) );
  MOAI22 U22278 ( .A1(n28235), .A2(n2394), .B1(ram[9124]), .B2(n2395), 
        .ZN(n13365) );
  MOAI22 U22279 ( .A1(n28000), .A2(n2394), .B1(ram[9125]), .B2(n2395), 
        .ZN(n13366) );
  MOAI22 U22280 ( .A1(n27765), .A2(n2394), .B1(ram[9126]), .B2(n2395), 
        .ZN(n13367) );
  MOAI22 U22281 ( .A1(n27530), .A2(n2394), .B1(ram[9127]), .B2(n2395), 
        .ZN(n13368) );
  MOAI22 U22282 ( .A1(n29175), .A2(n2396), .B1(ram[9128]), .B2(n2397), 
        .ZN(n13369) );
  MOAI22 U22283 ( .A1(n28940), .A2(n2396), .B1(ram[9129]), .B2(n2397), 
        .ZN(n13370) );
  MOAI22 U22284 ( .A1(n28705), .A2(n2396), .B1(ram[9130]), .B2(n2397), 
        .ZN(n13371) );
  MOAI22 U22285 ( .A1(n28470), .A2(n2396), .B1(ram[9131]), .B2(n2397), 
        .ZN(n13372) );
  MOAI22 U22286 ( .A1(n28235), .A2(n2396), .B1(ram[9132]), .B2(n2397), 
        .ZN(n13373) );
  MOAI22 U22287 ( .A1(n28000), .A2(n2396), .B1(ram[9133]), .B2(n2397), 
        .ZN(n13374) );
  MOAI22 U22288 ( .A1(n27765), .A2(n2396), .B1(ram[9134]), .B2(n2397), 
        .ZN(n13375) );
  MOAI22 U22289 ( .A1(n27530), .A2(n2396), .B1(ram[9135]), .B2(n2397), 
        .ZN(n13376) );
  MOAI22 U22290 ( .A1(n29175), .A2(n2398), .B1(ram[9136]), .B2(n2399), 
        .ZN(n13377) );
  MOAI22 U22291 ( .A1(n28940), .A2(n2398), .B1(ram[9137]), .B2(n2399), 
        .ZN(n13378) );
  MOAI22 U22292 ( .A1(n28705), .A2(n2398), .B1(ram[9138]), .B2(n2399), 
        .ZN(n13379) );
  MOAI22 U22293 ( .A1(n28470), .A2(n2398), .B1(ram[9139]), .B2(n2399), 
        .ZN(n13380) );
  MOAI22 U22294 ( .A1(n28235), .A2(n2398), .B1(ram[9140]), .B2(n2399), 
        .ZN(n13381) );
  MOAI22 U22295 ( .A1(n28000), .A2(n2398), .B1(ram[9141]), .B2(n2399), 
        .ZN(n13382) );
  MOAI22 U22296 ( .A1(n27765), .A2(n2398), .B1(ram[9142]), .B2(n2399), 
        .ZN(n13383) );
  MOAI22 U22297 ( .A1(n27530), .A2(n2398), .B1(ram[9143]), .B2(n2399), 
        .ZN(n13384) );
  MOAI22 U22298 ( .A1(n29175), .A2(n2400), .B1(ram[9144]), .B2(n2401), 
        .ZN(n13385) );
  MOAI22 U22299 ( .A1(n28940), .A2(n2400), .B1(ram[9145]), .B2(n2401), 
        .ZN(n13386) );
  MOAI22 U22300 ( .A1(n28705), .A2(n2400), .B1(ram[9146]), .B2(n2401), 
        .ZN(n13387) );
  MOAI22 U22301 ( .A1(n28470), .A2(n2400), .B1(ram[9147]), .B2(n2401), 
        .ZN(n13388) );
  MOAI22 U22302 ( .A1(n28235), .A2(n2400), .B1(ram[9148]), .B2(n2401), 
        .ZN(n13389) );
  MOAI22 U22303 ( .A1(n28000), .A2(n2400), .B1(ram[9149]), .B2(n2401), 
        .ZN(n13390) );
  MOAI22 U22304 ( .A1(n27765), .A2(n2400), .B1(ram[9150]), .B2(n2401), 
        .ZN(n13391) );
  MOAI22 U22305 ( .A1(n27530), .A2(n2400), .B1(ram[9151]), .B2(n2401), 
        .ZN(n13392) );
  MOAI22 U22306 ( .A1(n29176), .A2(n2402), .B1(ram[9152]), .B2(n2403), 
        .ZN(n13393) );
  MOAI22 U22307 ( .A1(n28941), .A2(n2402), .B1(ram[9153]), .B2(n2403), 
        .ZN(n13394) );
  MOAI22 U22308 ( .A1(n28706), .A2(n2402), .B1(ram[9154]), .B2(n2403), 
        .ZN(n13395) );
  MOAI22 U22309 ( .A1(n28471), .A2(n2402), .B1(ram[9155]), .B2(n2403), 
        .ZN(n13396) );
  MOAI22 U22310 ( .A1(n28236), .A2(n2402), .B1(ram[9156]), .B2(n2403), 
        .ZN(n13397) );
  MOAI22 U22311 ( .A1(n28001), .A2(n2402), .B1(ram[9157]), .B2(n2403), 
        .ZN(n13398) );
  MOAI22 U22312 ( .A1(n27766), .A2(n2402), .B1(ram[9158]), .B2(n2403), 
        .ZN(n13399) );
  MOAI22 U22313 ( .A1(n27531), .A2(n2402), .B1(ram[9159]), .B2(n2403), 
        .ZN(n13400) );
  MOAI22 U22314 ( .A1(n29176), .A2(n2404), .B1(ram[9160]), .B2(n2405), 
        .ZN(n13401) );
  MOAI22 U22315 ( .A1(n28941), .A2(n2404), .B1(ram[9161]), .B2(n2405), 
        .ZN(n13402) );
  MOAI22 U22316 ( .A1(n28706), .A2(n2404), .B1(ram[9162]), .B2(n2405), 
        .ZN(n13403) );
  MOAI22 U22317 ( .A1(n28471), .A2(n2404), .B1(ram[9163]), .B2(n2405), 
        .ZN(n13404) );
  MOAI22 U22318 ( .A1(n28236), .A2(n2404), .B1(ram[9164]), .B2(n2405), 
        .ZN(n13405) );
  MOAI22 U22319 ( .A1(n28001), .A2(n2404), .B1(ram[9165]), .B2(n2405), 
        .ZN(n13406) );
  MOAI22 U22320 ( .A1(n27766), .A2(n2404), .B1(ram[9166]), .B2(n2405), 
        .ZN(n13407) );
  MOAI22 U22321 ( .A1(n27531), .A2(n2404), .B1(ram[9167]), .B2(n2405), 
        .ZN(n13408) );
  MOAI22 U22322 ( .A1(n29176), .A2(n2406), .B1(ram[9168]), .B2(n2407), 
        .ZN(n13409) );
  MOAI22 U22323 ( .A1(n28941), .A2(n2406), .B1(ram[9169]), .B2(n2407), 
        .ZN(n13410) );
  MOAI22 U22324 ( .A1(n28706), .A2(n2406), .B1(ram[9170]), .B2(n2407), 
        .ZN(n13411) );
  MOAI22 U22325 ( .A1(n28471), .A2(n2406), .B1(ram[9171]), .B2(n2407), 
        .ZN(n13412) );
  MOAI22 U22326 ( .A1(n28236), .A2(n2406), .B1(ram[9172]), .B2(n2407), 
        .ZN(n13413) );
  MOAI22 U22327 ( .A1(n28001), .A2(n2406), .B1(ram[9173]), .B2(n2407), 
        .ZN(n13414) );
  MOAI22 U22328 ( .A1(n27766), .A2(n2406), .B1(ram[9174]), .B2(n2407), 
        .ZN(n13415) );
  MOAI22 U22329 ( .A1(n27531), .A2(n2406), .B1(ram[9175]), .B2(n2407), 
        .ZN(n13416) );
  MOAI22 U22330 ( .A1(n29176), .A2(n2408), .B1(ram[9176]), .B2(n2409), 
        .ZN(n13417) );
  MOAI22 U22331 ( .A1(n28941), .A2(n2408), .B1(ram[9177]), .B2(n2409), 
        .ZN(n13418) );
  MOAI22 U22332 ( .A1(n28706), .A2(n2408), .B1(ram[9178]), .B2(n2409), 
        .ZN(n13419) );
  MOAI22 U22333 ( .A1(n28471), .A2(n2408), .B1(ram[9179]), .B2(n2409), 
        .ZN(n13420) );
  MOAI22 U22334 ( .A1(n28236), .A2(n2408), .B1(ram[9180]), .B2(n2409), 
        .ZN(n13421) );
  MOAI22 U22335 ( .A1(n28001), .A2(n2408), .B1(ram[9181]), .B2(n2409), 
        .ZN(n13422) );
  MOAI22 U22336 ( .A1(n27766), .A2(n2408), .B1(ram[9182]), .B2(n2409), 
        .ZN(n13423) );
  MOAI22 U22337 ( .A1(n27531), .A2(n2408), .B1(ram[9183]), .B2(n2409), 
        .ZN(n13424) );
  MOAI22 U22338 ( .A1(n29176), .A2(n2410), .B1(ram[9184]), .B2(n2411), 
        .ZN(n13425) );
  MOAI22 U22339 ( .A1(n28941), .A2(n2410), .B1(ram[9185]), .B2(n2411), 
        .ZN(n13426) );
  MOAI22 U22340 ( .A1(n28706), .A2(n2410), .B1(ram[9186]), .B2(n2411), 
        .ZN(n13427) );
  MOAI22 U22341 ( .A1(n28471), .A2(n2410), .B1(ram[9187]), .B2(n2411), 
        .ZN(n13428) );
  MOAI22 U22342 ( .A1(n28236), .A2(n2410), .B1(ram[9188]), .B2(n2411), 
        .ZN(n13429) );
  MOAI22 U22343 ( .A1(n28001), .A2(n2410), .B1(ram[9189]), .B2(n2411), 
        .ZN(n13430) );
  MOAI22 U22344 ( .A1(n27766), .A2(n2410), .B1(ram[9190]), .B2(n2411), 
        .ZN(n13431) );
  MOAI22 U22345 ( .A1(n27531), .A2(n2410), .B1(ram[9191]), .B2(n2411), 
        .ZN(n13432) );
  MOAI22 U22346 ( .A1(n29176), .A2(n2412), .B1(ram[9192]), .B2(n2413), 
        .ZN(n13433) );
  MOAI22 U22347 ( .A1(n28941), .A2(n2412), .B1(ram[9193]), .B2(n2413), 
        .ZN(n13434) );
  MOAI22 U22348 ( .A1(n28706), .A2(n2412), .B1(ram[9194]), .B2(n2413), 
        .ZN(n13435) );
  MOAI22 U22349 ( .A1(n28471), .A2(n2412), .B1(ram[9195]), .B2(n2413), 
        .ZN(n13436) );
  MOAI22 U22350 ( .A1(n28236), .A2(n2412), .B1(ram[9196]), .B2(n2413), 
        .ZN(n13437) );
  MOAI22 U22351 ( .A1(n28001), .A2(n2412), .B1(ram[9197]), .B2(n2413), 
        .ZN(n13438) );
  MOAI22 U22352 ( .A1(n27766), .A2(n2412), .B1(ram[9198]), .B2(n2413), 
        .ZN(n13439) );
  MOAI22 U22353 ( .A1(n27531), .A2(n2412), .B1(ram[9199]), .B2(n2413), 
        .ZN(n13440) );
  MOAI22 U22354 ( .A1(n29176), .A2(n2414), .B1(ram[9200]), .B2(n2415), 
        .ZN(n13441) );
  MOAI22 U22355 ( .A1(n28941), .A2(n2414), .B1(ram[9201]), .B2(n2415), 
        .ZN(n13442) );
  MOAI22 U22356 ( .A1(n28706), .A2(n2414), .B1(ram[9202]), .B2(n2415), 
        .ZN(n13443) );
  MOAI22 U22357 ( .A1(n28471), .A2(n2414), .B1(ram[9203]), .B2(n2415), 
        .ZN(n13444) );
  MOAI22 U22358 ( .A1(n28236), .A2(n2414), .B1(ram[9204]), .B2(n2415), 
        .ZN(n13445) );
  MOAI22 U22359 ( .A1(n28001), .A2(n2414), .B1(ram[9205]), .B2(n2415), 
        .ZN(n13446) );
  MOAI22 U22360 ( .A1(n27766), .A2(n2414), .B1(ram[9206]), .B2(n2415), 
        .ZN(n13447) );
  MOAI22 U22361 ( .A1(n27531), .A2(n2414), .B1(ram[9207]), .B2(n2415), 
        .ZN(n13448) );
  MOAI22 U22362 ( .A1(n29176), .A2(n2416), .B1(ram[9208]), .B2(n2417), 
        .ZN(n13449) );
  MOAI22 U22363 ( .A1(n28941), .A2(n2416), .B1(ram[9209]), .B2(n2417), 
        .ZN(n13450) );
  MOAI22 U22364 ( .A1(n28706), .A2(n2416), .B1(ram[9210]), .B2(n2417), 
        .ZN(n13451) );
  MOAI22 U22365 ( .A1(n28471), .A2(n2416), .B1(ram[9211]), .B2(n2417), 
        .ZN(n13452) );
  MOAI22 U22366 ( .A1(n28236), .A2(n2416), .B1(ram[9212]), .B2(n2417), 
        .ZN(n13453) );
  MOAI22 U22367 ( .A1(n28001), .A2(n2416), .B1(ram[9213]), .B2(n2417), 
        .ZN(n13454) );
  MOAI22 U22368 ( .A1(n27766), .A2(n2416), .B1(ram[9214]), .B2(n2417), 
        .ZN(n13455) );
  MOAI22 U22369 ( .A1(n27531), .A2(n2416), .B1(ram[9215]), .B2(n2417), 
        .ZN(n13456) );
  MOAI22 U22370 ( .A1(n29176), .A2(n2418), .B1(ram[9216]), .B2(n2419), 
        .ZN(n13457) );
  MOAI22 U22371 ( .A1(n28941), .A2(n2418), .B1(ram[9217]), .B2(n2419), 
        .ZN(n13458) );
  MOAI22 U22372 ( .A1(n28706), .A2(n2418), .B1(ram[9218]), .B2(n2419), 
        .ZN(n13459) );
  MOAI22 U22373 ( .A1(n28471), .A2(n2418), .B1(ram[9219]), .B2(n2419), 
        .ZN(n13460) );
  MOAI22 U22374 ( .A1(n28236), .A2(n2418), .B1(ram[9220]), .B2(n2419), 
        .ZN(n13461) );
  MOAI22 U22375 ( .A1(n28001), .A2(n2418), .B1(ram[9221]), .B2(n2419), 
        .ZN(n13462) );
  MOAI22 U22376 ( .A1(n27766), .A2(n2418), .B1(ram[9222]), .B2(n2419), 
        .ZN(n13463) );
  MOAI22 U22377 ( .A1(n27531), .A2(n2418), .B1(ram[9223]), .B2(n2419), 
        .ZN(n13464) );
  MOAI22 U22378 ( .A1(n29176), .A2(n2421), .B1(ram[9224]), .B2(n2422), 
        .ZN(n13465) );
  MOAI22 U22379 ( .A1(n28941), .A2(n2421), .B1(ram[9225]), .B2(n2422), 
        .ZN(n13466) );
  MOAI22 U22380 ( .A1(n28706), .A2(n2421), .B1(ram[9226]), .B2(n2422), 
        .ZN(n13467) );
  MOAI22 U22381 ( .A1(n28471), .A2(n2421), .B1(ram[9227]), .B2(n2422), 
        .ZN(n13468) );
  MOAI22 U22382 ( .A1(n28236), .A2(n2421), .B1(ram[9228]), .B2(n2422), 
        .ZN(n13469) );
  MOAI22 U22383 ( .A1(n28001), .A2(n2421), .B1(ram[9229]), .B2(n2422), 
        .ZN(n13470) );
  MOAI22 U22384 ( .A1(n27766), .A2(n2421), .B1(ram[9230]), .B2(n2422), 
        .ZN(n13471) );
  MOAI22 U22385 ( .A1(n27531), .A2(n2421), .B1(ram[9231]), .B2(n2422), 
        .ZN(n13472) );
  MOAI22 U22386 ( .A1(n29176), .A2(n2423), .B1(ram[9232]), .B2(n2424), 
        .ZN(n13473) );
  MOAI22 U22387 ( .A1(n28941), .A2(n2423), .B1(ram[9233]), .B2(n2424), 
        .ZN(n13474) );
  MOAI22 U22388 ( .A1(n28706), .A2(n2423), .B1(ram[9234]), .B2(n2424), 
        .ZN(n13475) );
  MOAI22 U22389 ( .A1(n28471), .A2(n2423), .B1(ram[9235]), .B2(n2424), 
        .ZN(n13476) );
  MOAI22 U22390 ( .A1(n28236), .A2(n2423), .B1(ram[9236]), .B2(n2424), 
        .ZN(n13477) );
  MOAI22 U22391 ( .A1(n28001), .A2(n2423), .B1(ram[9237]), .B2(n2424), 
        .ZN(n13478) );
  MOAI22 U22392 ( .A1(n27766), .A2(n2423), .B1(ram[9238]), .B2(n2424), 
        .ZN(n13479) );
  MOAI22 U22393 ( .A1(n27531), .A2(n2423), .B1(ram[9239]), .B2(n2424), 
        .ZN(n13480) );
  MOAI22 U22394 ( .A1(n29176), .A2(n2425), .B1(ram[9240]), .B2(n2426), 
        .ZN(n13481) );
  MOAI22 U22395 ( .A1(n28941), .A2(n2425), .B1(ram[9241]), .B2(n2426), 
        .ZN(n13482) );
  MOAI22 U22396 ( .A1(n28706), .A2(n2425), .B1(ram[9242]), .B2(n2426), 
        .ZN(n13483) );
  MOAI22 U22397 ( .A1(n28471), .A2(n2425), .B1(ram[9243]), .B2(n2426), 
        .ZN(n13484) );
  MOAI22 U22398 ( .A1(n28236), .A2(n2425), .B1(ram[9244]), .B2(n2426), 
        .ZN(n13485) );
  MOAI22 U22399 ( .A1(n28001), .A2(n2425), .B1(ram[9245]), .B2(n2426), 
        .ZN(n13486) );
  MOAI22 U22400 ( .A1(n27766), .A2(n2425), .B1(ram[9246]), .B2(n2426), 
        .ZN(n13487) );
  MOAI22 U22401 ( .A1(n27531), .A2(n2425), .B1(ram[9247]), .B2(n2426), 
        .ZN(n13488) );
  MOAI22 U22402 ( .A1(n29176), .A2(n2427), .B1(ram[9248]), .B2(n2428), 
        .ZN(n13489) );
  MOAI22 U22403 ( .A1(n28941), .A2(n2427), .B1(ram[9249]), .B2(n2428), 
        .ZN(n13490) );
  MOAI22 U22404 ( .A1(n28706), .A2(n2427), .B1(ram[9250]), .B2(n2428), 
        .ZN(n13491) );
  MOAI22 U22405 ( .A1(n28471), .A2(n2427), .B1(ram[9251]), .B2(n2428), 
        .ZN(n13492) );
  MOAI22 U22406 ( .A1(n28236), .A2(n2427), .B1(ram[9252]), .B2(n2428), 
        .ZN(n13493) );
  MOAI22 U22407 ( .A1(n28001), .A2(n2427), .B1(ram[9253]), .B2(n2428), 
        .ZN(n13494) );
  MOAI22 U22408 ( .A1(n27766), .A2(n2427), .B1(ram[9254]), .B2(n2428), 
        .ZN(n13495) );
  MOAI22 U22409 ( .A1(n27531), .A2(n2427), .B1(ram[9255]), .B2(n2428), 
        .ZN(n13496) );
  MOAI22 U22410 ( .A1(n29177), .A2(n2429), .B1(ram[9256]), .B2(n2430), 
        .ZN(n13497) );
  MOAI22 U22411 ( .A1(n28942), .A2(n2429), .B1(ram[9257]), .B2(n2430), 
        .ZN(n13498) );
  MOAI22 U22412 ( .A1(n28707), .A2(n2429), .B1(ram[9258]), .B2(n2430), 
        .ZN(n13499) );
  MOAI22 U22413 ( .A1(n28472), .A2(n2429), .B1(ram[9259]), .B2(n2430), 
        .ZN(n13500) );
  MOAI22 U22414 ( .A1(n28237), .A2(n2429), .B1(ram[9260]), .B2(n2430), 
        .ZN(n13501) );
  MOAI22 U22415 ( .A1(n28002), .A2(n2429), .B1(ram[9261]), .B2(n2430), 
        .ZN(n13502) );
  MOAI22 U22416 ( .A1(n27767), .A2(n2429), .B1(ram[9262]), .B2(n2430), 
        .ZN(n13503) );
  MOAI22 U22417 ( .A1(n27532), .A2(n2429), .B1(ram[9263]), .B2(n2430), 
        .ZN(n13504) );
  MOAI22 U22418 ( .A1(n29177), .A2(n2431), .B1(ram[9264]), .B2(n2432), 
        .ZN(n13505) );
  MOAI22 U22419 ( .A1(n28942), .A2(n2431), .B1(ram[9265]), .B2(n2432), 
        .ZN(n13506) );
  MOAI22 U22420 ( .A1(n28707), .A2(n2431), .B1(ram[9266]), .B2(n2432), 
        .ZN(n13507) );
  MOAI22 U22421 ( .A1(n28472), .A2(n2431), .B1(ram[9267]), .B2(n2432), 
        .ZN(n13508) );
  MOAI22 U22422 ( .A1(n28237), .A2(n2431), .B1(ram[9268]), .B2(n2432), 
        .ZN(n13509) );
  MOAI22 U22423 ( .A1(n28002), .A2(n2431), .B1(ram[9269]), .B2(n2432), 
        .ZN(n13510) );
  MOAI22 U22424 ( .A1(n27767), .A2(n2431), .B1(ram[9270]), .B2(n2432), 
        .ZN(n13511) );
  MOAI22 U22425 ( .A1(n27532), .A2(n2431), .B1(ram[9271]), .B2(n2432), 
        .ZN(n13512) );
  MOAI22 U22426 ( .A1(n29177), .A2(n2433), .B1(ram[9272]), .B2(n2434), 
        .ZN(n13513) );
  MOAI22 U22427 ( .A1(n28942), .A2(n2433), .B1(ram[9273]), .B2(n2434), 
        .ZN(n13514) );
  MOAI22 U22428 ( .A1(n28707), .A2(n2433), .B1(ram[9274]), .B2(n2434), 
        .ZN(n13515) );
  MOAI22 U22429 ( .A1(n28472), .A2(n2433), .B1(ram[9275]), .B2(n2434), 
        .ZN(n13516) );
  MOAI22 U22430 ( .A1(n28237), .A2(n2433), .B1(ram[9276]), .B2(n2434), 
        .ZN(n13517) );
  MOAI22 U22431 ( .A1(n28002), .A2(n2433), .B1(ram[9277]), .B2(n2434), 
        .ZN(n13518) );
  MOAI22 U22432 ( .A1(n27767), .A2(n2433), .B1(ram[9278]), .B2(n2434), 
        .ZN(n13519) );
  MOAI22 U22433 ( .A1(n27532), .A2(n2433), .B1(ram[9279]), .B2(n2434), 
        .ZN(n13520) );
  MOAI22 U22434 ( .A1(n29177), .A2(n2435), .B1(ram[9280]), .B2(n2436), 
        .ZN(n13521) );
  MOAI22 U22435 ( .A1(n28942), .A2(n2435), .B1(ram[9281]), .B2(n2436), 
        .ZN(n13522) );
  MOAI22 U22436 ( .A1(n28707), .A2(n2435), .B1(ram[9282]), .B2(n2436), 
        .ZN(n13523) );
  MOAI22 U22437 ( .A1(n28472), .A2(n2435), .B1(ram[9283]), .B2(n2436), 
        .ZN(n13524) );
  MOAI22 U22438 ( .A1(n28237), .A2(n2435), .B1(ram[9284]), .B2(n2436), 
        .ZN(n13525) );
  MOAI22 U22439 ( .A1(n28002), .A2(n2435), .B1(ram[9285]), .B2(n2436), 
        .ZN(n13526) );
  MOAI22 U22440 ( .A1(n27767), .A2(n2435), .B1(ram[9286]), .B2(n2436), 
        .ZN(n13527) );
  MOAI22 U22441 ( .A1(n27532), .A2(n2435), .B1(ram[9287]), .B2(n2436), 
        .ZN(n13528) );
  MOAI22 U22442 ( .A1(n29177), .A2(n2437), .B1(ram[9288]), .B2(n2438), 
        .ZN(n13529) );
  MOAI22 U22443 ( .A1(n28942), .A2(n2437), .B1(ram[9289]), .B2(n2438), 
        .ZN(n13530) );
  MOAI22 U22444 ( .A1(n28707), .A2(n2437), .B1(ram[9290]), .B2(n2438), 
        .ZN(n13531) );
  MOAI22 U22445 ( .A1(n28472), .A2(n2437), .B1(ram[9291]), .B2(n2438), 
        .ZN(n13532) );
  MOAI22 U22446 ( .A1(n28237), .A2(n2437), .B1(ram[9292]), .B2(n2438), 
        .ZN(n13533) );
  MOAI22 U22447 ( .A1(n28002), .A2(n2437), .B1(ram[9293]), .B2(n2438), 
        .ZN(n13534) );
  MOAI22 U22448 ( .A1(n27767), .A2(n2437), .B1(ram[9294]), .B2(n2438), 
        .ZN(n13535) );
  MOAI22 U22449 ( .A1(n27532), .A2(n2437), .B1(ram[9295]), .B2(n2438), 
        .ZN(n13536) );
  MOAI22 U22450 ( .A1(n29177), .A2(n2439), .B1(ram[9296]), .B2(n2440), 
        .ZN(n13537) );
  MOAI22 U22451 ( .A1(n28942), .A2(n2439), .B1(ram[9297]), .B2(n2440), 
        .ZN(n13538) );
  MOAI22 U22452 ( .A1(n28707), .A2(n2439), .B1(ram[9298]), .B2(n2440), 
        .ZN(n13539) );
  MOAI22 U22453 ( .A1(n28472), .A2(n2439), .B1(ram[9299]), .B2(n2440), 
        .ZN(n13540) );
  MOAI22 U22454 ( .A1(n28237), .A2(n2439), .B1(ram[9300]), .B2(n2440), 
        .ZN(n13541) );
  MOAI22 U22455 ( .A1(n28002), .A2(n2439), .B1(ram[9301]), .B2(n2440), 
        .ZN(n13542) );
  MOAI22 U22456 ( .A1(n27767), .A2(n2439), .B1(ram[9302]), .B2(n2440), 
        .ZN(n13543) );
  MOAI22 U22457 ( .A1(n27532), .A2(n2439), .B1(ram[9303]), .B2(n2440), 
        .ZN(n13544) );
  MOAI22 U22458 ( .A1(n29177), .A2(n2441), .B1(ram[9304]), .B2(n2442), 
        .ZN(n13545) );
  MOAI22 U22459 ( .A1(n28942), .A2(n2441), .B1(ram[9305]), .B2(n2442), 
        .ZN(n13546) );
  MOAI22 U22460 ( .A1(n28707), .A2(n2441), .B1(ram[9306]), .B2(n2442), 
        .ZN(n13547) );
  MOAI22 U22461 ( .A1(n28472), .A2(n2441), .B1(ram[9307]), .B2(n2442), 
        .ZN(n13548) );
  MOAI22 U22462 ( .A1(n28237), .A2(n2441), .B1(ram[9308]), .B2(n2442), 
        .ZN(n13549) );
  MOAI22 U22463 ( .A1(n28002), .A2(n2441), .B1(ram[9309]), .B2(n2442), 
        .ZN(n13550) );
  MOAI22 U22464 ( .A1(n27767), .A2(n2441), .B1(ram[9310]), .B2(n2442), 
        .ZN(n13551) );
  MOAI22 U22465 ( .A1(n27532), .A2(n2441), .B1(ram[9311]), .B2(n2442), 
        .ZN(n13552) );
  MOAI22 U22466 ( .A1(n29177), .A2(n2443), .B1(ram[9312]), .B2(n2444), 
        .ZN(n13553) );
  MOAI22 U22467 ( .A1(n28942), .A2(n2443), .B1(ram[9313]), .B2(n2444), 
        .ZN(n13554) );
  MOAI22 U22468 ( .A1(n28707), .A2(n2443), .B1(ram[9314]), .B2(n2444), 
        .ZN(n13555) );
  MOAI22 U22469 ( .A1(n28472), .A2(n2443), .B1(ram[9315]), .B2(n2444), 
        .ZN(n13556) );
  MOAI22 U22470 ( .A1(n28237), .A2(n2443), .B1(ram[9316]), .B2(n2444), 
        .ZN(n13557) );
  MOAI22 U22471 ( .A1(n28002), .A2(n2443), .B1(ram[9317]), .B2(n2444), 
        .ZN(n13558) );
  MOAI22 U22472 ( .A1(n27767), .A2(n2443), .B1(ram[9318]), .B2(n2444), 
        .ZN(n13559) );
  MOAI22 U22473 ( .A1(n27532), .A2(n2443), .B1(ram[9319]), .B2(n2444), 
        .ZN(n13560) );
  MOAI22 U22474 ( .A1(n29177), .A2(n2445), .B1(ram[9320]), .B2(n2446), 
        .ZN(n13561) );
  MOAI22 U22475 ( .A1(n28942), .A2(n2445), .B1(ram[9321]), .B2(n2446), 
        .ZN(n13562) );
  MOAI22 U22476 ( .A1(n28707), .A2(n2445), .B1(ram[9322]), .B2(n2446), 
        .ZN(n13563) );
  MOAI22 U22477 ( .A1(n28472), .A2(n2445), .B1(ram[9323]), .B2(n2446), 
        .ZN(n13564) );
  MOAI22 U22478 ( .A1(n28237), .A2(n2445), .B1(ram[9324]), .B2(n2446), 
        .ZN(n13565) );
  MOAI22 U22479 ( .A1(n28002), .A2(n2445), .B1(ram[9325]), .B2(n2446), 
        .ZN(n13566) );
  MOAI22 U22480 ( .A1(n27767), .A2(n2445), .B1(ram[9326]), .B2(n2446), 
        .ZN(n13567) );
  MOAI22 U22481 ( .A1(n27532), .A2(n2445), .B1(ram[9327]), .B2(n2446), 
        .ZN(n13568) );
  MOAI22 U22482 ( .A1(n29177), .A2(n2447), .B1(ram[9328]), .B2(n2448), 
        .ZN(n13569) );
  MOAI22 U22483 ( .A1(n28942), .A2(n2447), .B1(ram[9329]), .B2(n2448), 
        .ZN(n13570) );
  MOAI22 U22484 ( .A1(n28707), .A2(n2447), .B1(ram[9330]), .B2(n2448), 
        .ZN(n13571) );
  MOAI22 U22485 ( .A1(n28472), .A2(n2447), .B1(ram[9331]), .B2(n2448), 
        .ZN(n13572) );
  MOAI22 U22486 ( .A1(n28237), .A2(n2447), .B1(ram[9332]), .B2(n2448), 
        .ZN(n13573) );
  MOAI22 U22487 ( .A1(n28002), .A2(n2447), .B1(ram[9333]), .B2(n2448), 
        .ZN(n13574) );
  MOAI22 U22488 ( .A1(n27767), .A2(n2447), .B1(ram[9334]), .B2(n2448), 
        .ZN(n13575) );
  MOAI22 U22489 ( .A1(n27532), .A2(n2447), .B1(ram[9335]), .B2(n2448), 
        .ZN(n13576) );
  MOAI22 U22490 ( .A1(n29177), .A2(n2449), .B1(ram[9336]), .B2(n2450), 
        .ZN(n13577) );
  MOAI22 U22491 ( .A1(n28942), .A2(n2449), .B1(ram[9337]), .B2(n2450), 
        .ZN(n13578) );
  MOAI22 U22492 ( .A1(n28707), .A2(n2449), .B1(ram[9338]), .B2(n2450), 
        .ZN(n13579) );
  MOAI22 U22493 ( .A1(n28472), .A2(n2449), .B1(ram[9339]), .B2(n2450), 
        .ZN(n13580) );
  MOAI22 U22494 ( .A1(n28237), .A2(n2449), .B1(ram[9340]), .B2(n2450), 
        .ZN(n13581) );
  MOAI22 U22495 ( .A1(n28002), .A2(n2449), .B1(ram[9341]), .B2(n2450), 
        .ZN(n13582) );
  MOAI22 U22496 ( .A1(n27767), .A2(n2449), .B1(ram[9342]), .B2(n2450), 
        .ZN(n13583) );
  MOAI22 U22497 ( .A1(n27532), .A2(n2449), .B1(ram[9343]), .B2(n2450), 
        .ZN(n13584) );
  MOAI22 U22498 ( .A1(n29177), .A2(n2451), .B1(ram[9344]), .B2(n2452), 
        .ZN(n13585) );
  MOAI22 U22499 ( .A1(n28942), .A2(n2451), .B1(ram[9345]), .B2(n2452), 
        .ZN(n13586) );
  MOAI22 U22500 ( .A1(n28707), .A2(n2451), .B1(ram[9346]), .B2(n2452), 
        .ZN(n13587) );
  MOAI22 U22501 ( .A1(n28472), .A2(n2451), .B1(ram[9347]), .B2(n2452), 
        .ZN(n13588) );
  MOAI22 U22502 ( .A1(n28237), .A2(n2451), .B1(ram[9348]), .B2(n2452), 
        .ZN(n13589) );
  MOAI22 U22503 ( .A1(n28002), .A2(n2451), .B1(ram[9349]), .B2(n2452), 
        .ZN(n13590) );
  MOAI22 U22504 ( .A1(n27767), .A2(n2451), .B1(ram[9350]), .B2(n2452), 
        .ZN(n13591) );
  MOAI22 U22505 ( .A1(n27532), .A2(n2451), .B1(ram[9351]), .B2(n2452), 
        .ZN(n13592) );
  MOAI22 U22506 ( .A1(n29177), .A2(n2453), .B1(ram[9352]), .B2(n2454), 
        .ZN(n13593) );
  MOAI22 U22507 ( .A1(n28942), .A2(n2453), .B1(ram[9353]), .B2(n2454), 
        .ZN(n13594) );
  MOAI22 U22508 ( .A1(n28707), .A2(n2453), .B1(ram[9354]), .B2(n2454), 
        .ZN(n13595) );
  MOAI22 U22509 ( .A1(n28472), .A2(n2453), .B1(ram[9355]), .B2(n2454), 
        .ZN(n13596) );
  MOAI22 U22510 ( .A1(n28237), .A2(n2453), .B1(ram[9356]), .B2(n2454), 
        .ZN(n13597) );
  MOAI22 U22511 ( .A1(n28002), .A2(n2453), .B1(ram[9357]), .B2(n2454), 
        .ZN(n13598) );
  MOAI22 U22512 ( .A1(n27767), .A2(n2453), .B1(ram[9358]), .B2(n2454), 
        .ZN(n13599) );
  MOAI22 U22513 ( .A1(n27532), .A2(n2453), .B1(ram[9359]), .B2(n2454), 
        .ZN(n13600) );
  MOAI22 U22514 ( .A1(n29178), .A2(n2455), .B1(ram[9360]), .B2(n2456), 
        .ZN(n13601) );
  MOAI22 U22515 ( .A1(n28943), .A2(n2455), .B1(ram[9361]), .B2(n2456), 
        .ZN(n13602) );
  MOAI22 U22516 ( .A1(n28708), .A2(n2455), .B1(ram[9362]), .B2(n2456), 
        .ZN(n13603) );
  MOAI22 U22517 ( .A1(n28473), .A2(n2455), .B1(ram[9363]), .B2(n2456), 
        .ZN(n13604) );
  MOAI22 U22518 ( .A1(n28238), .A2(n2455), .B1(ram[9364]), .B2(n2456), 
        .ZN(n13605) );
  MOAI22 U22519 ( .A1(n28003), .A2(n2455), .B1(ram[9365]), .B2(n2456), 
        .ZN(n13606) );
  MOAI22 U22520 ( .A1(n27768), .A2(n2455), .B1(ram[9366]), .B2(n2456), 
        .ZN(n13607) );
  MOAI22 U22521 ( .A1(n27533), .A2(n2455), .B1(ram[9367]), .B2(n2456), 
        .ZN(n13608) );
  MOAI22 U22522 ( .A1(n29178), .A2(n2457), .B1(ram[9368]), .B2(n2458), 
        .ZN(n13609) );
  MOAI22 U22523 ( .A1(n28943), .A2(n2457), .B1(ram[9369]), .B2(n2458), 
        .ZN(n13610) );
  MOAI22 U22524 ( .A1(n28708), .A2(n2457), .B1(ram[9370]), .B2(n2458), 
        .ZN(n13611) );
  MOAI22 U22525 ( .A1(n28473), .A2(n2457), .B1(ram[9371]), .B2(n2458), 
        .ZN(n13612) );
  MOAI22 U22526 ( .A1(n28238), .A2(n2457), .B1(ram[9372]), .B2(n2458), 
        .ZN(n13613) );
  MOAI22 U22527 ( .A1(n28003), .A2(n2457), .B1(ram[9373]), .B2(n2458), 
        .ZN(n13614) );
  MOAI22 U22528 ( .A1(n27768), .A2(n2457), .B1(ram[9374]), .B2(n2458), 
        .ZN(n13615) );
  MOAI22 U22529 ( .A1(n27533), .A2(n2457), .B1(ram[9375]), .B2(n2458), 
        .ZN(n13616) );
  MOAI22 U22530 ( .A1(n29178), .A2(n2459), .B1(ram[9376]), .B2(n2460), 
        .ZN(n13617) );
  MOAI22 U22531 ( .A1(n28943), .A2(n2459), .B1(ram[9377]), .B2(n2460), 
        .ZN(n13618) );
  MOAI22 U22532 ( .A1(n28708), .A2(n2459), .B1(ram[9378]), .B2(n2460), 
        .ZN(n13619) );
  MOAI22 U22533 ( .A1(n28473), .A2(n2459), .B1(ram[9379]), .B2(n2460), 
        .ZN(n13620) );
  MOAI22 U22534 ( .A1(n28238), .A2(n2459), .B1(ram[9380]), .B2(n2460), 
        .ZN(n13621) );
  MOAI22 U22535 ( .A1(n28003), .A2(n2459), .B1(ram[9381]), .B2(n2460), 
        .ZN(n13622) );
  MOAI22 U22536 ( .A1(n27768), .A2(n2459), .B1(ram[9382]), .B2(n2460), 
        .ZN(n13623) );
  MOAI22 U22537 ( .A1(n27533), .A2(n2459), .B1(ram[9383]), .B2(n2460), 
        .ZN(n13624) );
  MOAI22 U22538 ( .A1(n29178), .A2(n2461), .B1(ram[9384]), .B2(n2462), 
        .ZN(n13625) );
  MOAI22 U22539 ( .A1(n28943), .A2(n2461), .B1(ram[9385]), .B2(n2462), 
        .ZN(n13626) );
  MOAI22 U22540 ( .A1(n28708), .A2(n2461), .B1(ram[9386]), .B2(n2462), 
        .ZN(n13627) );
  MOAI22 U22541 ( .A1(n28473), .A2(n2461), .B1(ram[9387]), .B2(n2462), 
        .ZN(n13628) );
  MOAI22 U22542 ( .A1(n28238), .A2(n2461), .B1(ram[9388]), .B2(n2462), 
        .ZN(n13629) );
  MOAI22 U22543 ( .A1(n28003), .A2(n2461), .B1(ram[9389]), .B2(n2462), 
        .ZN(n13630) );
  MOAI22 U22544 ( .A1(n27768), .A2(n2461), .B1(ram[9390]), .B2(n2462), 
        .ZN(n13631) );
  MOAI22 U22545 ( .A1(n27533), .A2(n2461), .B1(ram[9391]), .B2(n2462), 
        .ZN(n13632) );
  MOAI22 U22546 ( .A1(n29178), .A2(n2463), .B1(ram[9392]), .B2(n2464), 
        .ZN(n13633) );
  MOAI22 U22547 ( .A1(n28943), .A2(n2463), .B1(ram[9393]), .B2(n2464), 
        .ZN(n13634) );
  MOAI22 U22548 ( .A1(n28708), .A2(n2463), .B1(ram[9394]), .B2(n2464), 
        .ZN(n13635) );
  MOAI22 U22549 ( .A1(n28473), .A2(n2463), .B1(ram[9395]), .B2(n2464), 
        .ZN(n13636) );
  MOAI22 U22550 ( .A1(n28238), .A2(n2463), .B1(ram[9396]), .B2(n2464), 
        .ZN(n13637) );
  MOAI22 U22551 ( .A1(n28003), .A2(n2463), .B1(ram[9397]), .B2(n2464), 
        .ZN(n13638) );
  MOAI22 U22552 ( .A1(n27768), .A2(n2463), .B1(ram[9398]), .B2(n2464), 
        .ZN(n13639) );
  MOAI22 U22553 ( .A1(n27533), .A2(n2463), .B1(ram[9399]), .B2(n2464), 
        .ZN(n13640) );
  MOAI22 U22554 ( .A1(n29178), .A2(n2465), .B1(ram[9400]), .B2(n2466), 
        .ZN(n13641) );
  MOAI22 U22555 ( .A1(n28943), .A2(n2465), .B1(ram[9401]), .B2(n2466), 
        .ZN(n13642) );
  MOAI22 U22556 ( .A1(n28708), .A2(n2465), .B1(ram[9402]), .B2(n2466), 
        .ZN(n13643) );
  MOAI22 U22557 ( .A1(n28473), .A2(n2465), .B1(ram[9403]), .B2(n2466), 
        .ZN(n13644) );
  MOAI22 U22558 ( .A1(n28238), .A2(n2465), .B1(ram[9404]), .B2(n2466), 
        .ZN(n13645) );
  MOAI22 U22559 ( .A1(n28003), .A2(n2465), .B1(ram[9405]), .B2(n2466), 
        .ZN(n13646) );
  MOAI22 U22560 ( .A1(n27768), .A2(n2465), .B1(ram[9406]), .B2(n2466), 
        .ZN(n13647) );
  MOAI22 U22561 ( .A1(n27533), .A2(n2465), .B1(ram[9407]), .B2(n2466), 
        .ZN(n13648) );
  MOAI22 U22562 ( .A1(n29178), .A2(n2467), .B1(ram[9408]), .B2(n2468), 
        .ZN(n13649) );
  MOAI22 U22563 ( .A1(n28943), .A2(n2467), .B1(ram[9409]), .B2(n2468), 
        .ZN(n13650) );
  MOAI22 U22564 ( .A1(n28708), .A2(n2467), .B1(ram[9410]), .B2(n2468), 
        .ZN(n13651) );
  MOAI22 U22565 ( .A1(n28473), .A2(n2467), .B1(ram[9411]), .B2(n2468), 
        .ZN(n13652) );
  MOAI22 U22566 ( .A1(n28238), .A2(n2467), .B1(ram[9412]), .B2(n2468), 
        .ZN(n13653) );
  MOAI22 U22567 ( .A1(n28003), .A2(n2467), .B1(ram[9413]), .B2(n2468), 
        .ZN(n13654) );
  MOAI22 U22568 ( .A1(n27768), .A2(n2467), .B1(ram[9414]), .B2(n2468), 
        .ZN(n13655) );
  MOAI22 U22569 ( .A1(n27533), .A2(n2467), .B1(ram[9415]), .B2(n2468), 
        .ZN(n13656) );
  MOAI22 U22570 ( .A1(n29178), .A2(n2469), .B1(ram[9416]), .B2(n2470), 
        .ZN(n13657) );
  MOAI22 U22571 ( .A1(n28943), .A2(n2469), .B1(ram[9417]), .B2(n2470), 
        .ZN(n13658) );
  MOAI22 U22572 ( .A1(n28708), .A2(n2469), .B1(ram[9418]), .B2(n2470), 
        .ZN(n13659) );
  MOAI22 U22573 ( .A1(n28473), .A2(n2469), .B1(ram[9419]), .B2(n2470), 
        .ZN(n13660) );
  MOAI22 U22574 ( .A1(n28238), .A2(n2469), .B1(ram[9420]), .B2(n2470), 
        .ZN(n13661) );
  MOAI22 U22575 ( .A1(n28003), .A2(n2469), .B1(ram[9421]), .B2(n2470), 
        .ZN(n13662) );
  MOAI22 U22576 ( .A1(n27768), .A2(n2469), .B1(ram[9422]), .B2(n2470), 
        .ZN(n13663) );
  MOAI22 U22577 ( .A1(n27533), .A2(n2469), .B1(ram[9423]), .B2(n2470), 
        .ZN(n13664) );
  MOAI22 U22578 ( .A1(n29178), .A2(n2471), .B1(ram[9424]), .B2(n2472), 
        .ZN(n13665) );
  MOAI22 U22579 ( .A1(n28943), .A2(n2471), .B1(ram[9425]), .B2(n2472), 
        .ZN(n13666) );
  MOAI22 U22580 ( .A1(n28708), .A2(n2471), .B1(ram[9426]), .B2(n2472), 
        .ZN(n13667) );
  MOAI22 U22581 ( .A1(n28473), .A2(n2471), .B1(ram[9427]), .B2(n2472), 
        .ZN(n13668) );
  MOAI22 U22582 ( .A1(n28238), .A2(n2471), .B1(ram[9428]), .B2(n2472), 
        .ZN(n13669) );
  MOAI22 U22583 ( .A1(n28003), .A2(n2471), .B1(ram[9429]), .B2(n2472), 
        .ZN(n13670) );
  MOAI22 U22584 ( .A1(n27768), .A2(n2471), .B1(ram[9430]), .B2(n2472), 
        .ZN(n13671) );
  MOAI22 U22585 ( .A1(n27533), .A2(n2471), .B1(ram[9431]), .B2(n2472), 
        .ZN(n13672) );
  MOAI22 U22586 ( .A1(n29178), .A2(n2473), .B1(ram[9432]), .B2(n2474), 
        .ZN(n13673) );
  MOAI22 U22587 ( .A1(n28943), .A2(n2473), .B1(ram[9433]), .B2(n2474), 
        .ZN(n13674) );
  MOAI22 U22588 ( .A1(n28708), .A2(n2473), .B1(ram[9434]), .B2(n2474), 
        .ZN(n13675) );
  MOAI22 U22589 ( .A1(n28473), .A2(n2473), .B1(ram[9435]), .B2(n2474), 
        .ZN(n13676) );
  MOAI22 U22590 ( .A1(n28238), .A2(n2473), .B1(ram[9436]), .B2(n2474), 
        .ZN(n13677) );
  MOAI22 U22591 ( .A1(n28003), .A2(n2473), .B1(ram[9437]), .B2(n2474), 
        .ZN(n13678) );
  MOAI22 U22592 ( .A1(n27768), .A2(n2473), .B1(ram[9438]), .B2(n2474), 
        .ZN(n13679) );
  MOAI22 U22593 ( .A1(n27533), .A2(n2473), .B1(ram[9439]), .B2(n2474), 
        .ZN(n13680) );
  MOAI22 U22594 ( .A1(n29178), .A2(n2475), .B1(ram[9440]), .B2(n2476), 
        .ZN(n13681) );
  MOAI22 U22595 ( .A1(n28943), .A2(n2475), .B1(ram[9441]), .B2(n2476), 
        .ZN(n13682) );
  MOAI22 U22596 ( .A1(n28708), .A2(n2475), .B1(ram[9442]), .B2(n2476), 
        .ZN(n13683) );
  MOAI22 U22597 ( .A1(n28473), .A2(n2475), .B1(ram[9443]), .B2(n2476), 
        .ZN(n13684) );
  MOAI22 U22598 ( .A1(n28238), .A2(n2475), .B1(ram[9444]), .B2(n2476), 
        .ZN(n13685) );
  MOAI22 U22599 ( .A1(n28003), .A2(n2475), .B1(ram[9445]), .B2(n2476), 
        .ZN(n13686) );
  MOAI22 U22600 ( .A1(n27768), .A2(n2475), .B1(ram[9446]), .B2(n2476), 
        .ZN(n13687) );
  MOAI22 U22601 ( .A1(n27533), .A2(n2475), .B1(ram[9447]), .B2(n2476), 
        .ZN(n13688) );
  MOAI22 U22602 ( .A1(n29178), .A2(n2477), .B1(ram[9448]), .B2(n2478), 
        .ZN(n13689) );
  MOAI22 U22603 ( .A1(n28943), .A2(n2477), .B1(ram[9449]), .B2(n2478), 
        .ZN(n13690) );
  MOAI22 U22604 ( .A1(n28708), .A2(n2477), .B1(ram[9450]), .B2(n2478), 
        .ZN(n13691) );
  MOAI22 U22605 ( .A1(n28473), .A2(n2477), .B1(ram[9451]), .B2(n2478), 
        .ZN(n13692) );
  MOAI22 U22606 ( .A1(n28238), .A2(n2477), .B1(ram[9452]), .B2(n2478), 
        .ZN(n13693) );
  MOAI22 U22607 ( .A1(n28003), .A2(n2477), .B1(ram[9453]), .B2(n2478), 
        .ZN(n13694) );
  MOAI22 U22608 ( .A1(n27768), .A2(n2477), .B1(ram[9454]), .B2(n2478), 
        .ZN(n13695) );
  MOAI22 U22609 ( .A1(n27533), .A2(n2477), .B1(ram[9455]), .B2(n2478), 
        .ZN(n13696) );
  MOAI22 U22610 ( .A1(n29178), .A2(n2479), .B1(ram[9456]), .B2(n2480), 
        .ZN(n13697) );
  MOAI22 U22611 ( .A1(n28943), .A2(n2479), .B1(ram[9457]), .B2(n2480), 
        .ZN(n13698) );
  MOAI22 U22612 ( .A1(n28708), .A2(n2479), .B1(ram[9458]), .B2(n2480), 
        .ZN(n13699) );
  MOAI22 U22613 ( .A1(n28473), .A2(n2479), .B1(ram[9459]), .B2(n2480), 
        .ZN(n13700) );
  MOAI22 U22614 ( .A1(n28238), .A2(n2479), .B1(ram[9460]), .B2(n2480), 
        .ZN(n13701) );
  MOAI22 U22615 ( .A1(n28003), .A2(n2479), .B1(ram[9461]), .B2(n2480), 
        .ZN(n13702) );
  MOAI22 U22616 ( .A1(n27768), .A2(n2479), .B1(ram[9462]), .B2(n2480), 
        .ZN(n13703) );
  MOAI22 U22617 ( .A1(n27533), .A2(n2479), .B1(ram[9463]), .B2(n2480), 
        .ZN(n13704) );
  MOAI22 U22618 ( .A1(n29179), .A2(n2481), .B1(ram[9464]), .B2(n2482), 
        .ZN(n13705) );
  MOAI22 U22619 ( .A1(n28944), .A2(n2481), .B1(ram[9465]), .B2(n2482), 
        .ZN(n13706) );
  MOAI22 U22620 ( .A1(n28709), .A2(n2481), .B1(ram[9466]), .B2(n2482), 
        .ZN(n13707) );
  MOAI22 U22621 ( .A1(n28474), .A2(n2481), .B1(ram[9467]), .B2(n2482), 
        .ZN(n13708) );
  MOAI22 U22622 ( .A1(n28239), .A2(n2481), .B1(ram[9468]), .B2(n2482), 
        .ZN(n13709) );
  MOAI22 U22623 ( .A1(n28004), .A2(n2481), .B1(ram[9469]), .B2(n2482), 
        .ZN(n13710) );
  MOAI22 U22624 ( .A1(n27769), .A2(n2481), .B1(ram[9470]), .B2(n2482), 
        .ZN(n13711) );
  MOAI22 U22625 ( .A1(n27534), .A2(n2481), .B1(ram[9471]), .B2(n2482), 
        .ZN(n13712) );
  MOAI22 U22626 ( .A1(n29179), .A2(n2483), .B1(ram[9472]), .B2(n2484), 
        .ZN(n13713) );
  MOAI22 U22627 ( .A1(n28944), .A2(n2483), .B1(ram[9473]), .B2(n2484), 
        .ZN(n13714) );
  MOAI22 U22628 ( .A1(n28709), .A2(n2483), .B1(ram[9474]), .B2(n2484), 
        .ZN(n13715) );
  MOAI22 U22629 ( .A1(n28474), .A2(n2483), .B1(ram[9475]), .B2(n2484), 
        .ZN(n13716) );
  MOAI22 U22630 ( .A1(n28239), .A2(n2483), .B1(ram[9476]), .B2(n2484), 
        .ZN(n13717) );
  MOAI22 U22631 ( .A1(n28004), .A2(n2483), .B1(ram[9477]), .B2(n2484), 
        .ZN(n13718) );
  MOAI22 U22632 ( .A1(n27769), .A2(n2483), .B1(ram[9478]), .B2(n2484), 
        .ZN(n13719) );
  MOAI22 U22633 ( .A1(n27534), .A2(n2483), .B1(ram[9479]), .B2(n2484), 
        .ZN(n13720) );
  MOAI22 U22634 ( .A1(n29179), .A2(n2485), .B1(ram[9480]), .B2(n2486), 
        .ZN(n13721) );
  MOAI22 U22635 ( .A1(n28944), .A2(n2485), .B1(ram[9481]), .B2(n2486), 
        .ZN(n13722) );
  MOAI22 U22636 ( .A1(n28709), .A2(n2485), .B1(ram[9482]), .B2(n2486), 
        .ZN(n13723) );
  MOAI22 U22637 ( .A1(n28474), .A2(n2485), .B1(ram[9483]), .B2(n2486), 
        .ZN(n13724) );
  MOAI22 U22638 ( .A1(n28239), .A2(n2485), .B1(ram[9484]), .B2(n2486), 
        .ZN(n13725) );
  MOAI22 U22639 ( .A1(n28004), .A2(n2485), .B1(ram[9485]), .B2(n2486), 
        .ZN(n13726) );
  MOAI22 U22640 ( .A1(n27769), .A2(n2485), .B1(ram[9486]), .B2(n2486), 
        .ZN(n13727) );
  MOAI22 U22641 ( .A1(n27534), .A2(n2485), .B1(ram[9487]), .B2(n2486), 
        .ZN(n13728) );
  MOAI22 U22642 ( .A1(n29179), .A2(n2487), .B1(ram[9488]), .B2(n2488), 
        .ZN(n13729) );
  MOAI22 U22643 ( .A1(n28944), .A2(n2487), .B1(ram[9489]), .B2(n2488), 
        .ZN(n13730) );
  MOAI22 U22644 ( .A1(n28709), .A2(n2487), .B1(ram[9490]), .B2(n2488), 
        .ZN(n13731) );
  MOAI22 U22645 ( .A1(n28474), .A2(n2487), .B1(ram[9491]), .B2(n2488), 
        .ZN(n13732) );
  MOAI22 U22646 ( .A1(n28239), .A2(n2487), .B1(ram[9492]), .B2(n2488), 
        .ZN(n13733) );
  MOAI22 U22647 ( .A1(n28004), .A2(n2487), .B1(ram[9493]), .B2(n2488), 
        .ZN(n13734) );
  MOAI22 U22648 ( .A1(n27769), .A2(n2487), .B1(ram[9494]), .B2(n2488), 
        .ZN(n13735) );
  MOAI22 U22649 ( .A1(n27534), .A2(n2487), .B1(ram[9495]), .B2(n2488), 
        .ZN(n13736) );
  MOAI22 U22650 ( .A1(n29179), .A2(n2489), .B1(ram[9496]), .B2(n2490), 
        .ZN(n13737) );
  MOAI22 U22651 ( .A1(n28944), .A2(n2489), .B1(ram[9497]), .B2(n2490), 
        .ZN(n13738) );
  MOAI22 U22652 ( .A1(n28709), .A2(n2489), .B1(ram[9498]), .B2(n2490), 
        .ZN(n13739) );
  MOAI22 U22653 ( .A1(n28474), .A2(n2489), .B1(ram[9499]), .B2(n2490), 
        .ZN(n13740) );
  MOAI22 U22654 ( .A1(n28239), .A2(n2489), .B1(ram[9500]), .B2(n2490), 
        .ZN(n13741) );
  MOAI22 U22655 ( .A1(n28004), .A2(n2489), .B1(ram[9501]), .B2(n2490), 
        .ZN(n13742) );
  MOAI22 U22656 ( .A1(n27769), .A2(n2489), .B1(ram[9502]), .B2(n2490), 
        .ZN(n13743) );
  MOAI22 U22657 ( .A1(n27534), .A2(n2489), .B1(ram[9503]), .B2(n2490), 
        .ZN(n13744) );
  MOAI22 U22658 ( .A1(n29179), .A2(n2491), .B1(ram[9504]), .B2(n2492), 
        .ZN(n13745) );
  MOAI22 U22659 ( .A1(n28944), .A2(n2491), .B1(ram[9505]), .B2(n2492), 
        .ZN(n13746) );
  MOAI22 U22660 ( .A1(n28709), .A2(n2491), .B1(ram[9506]), .B2(n2492), 
        .ZN(n13747) );
  MOAI22 U22661 ( .A1(n28474), .A2(n2491), .B1(ram[9507]), .B2(n2492), 
        .ZN(n13748) );
  MOAI22 U22662 ( .A1(n28239), .A2(n2491), .B1(ram[9508]), .B2(n2492), 
        .ZN(n13749) );
  MOAI22 U22663 ( .A1(n28004), .A2(n2491), .B1(ram[9509]), .B2(n2492), 
        .ZN(n13750) );
  MOAI22 U22664 ( .A1(n27769), .A2(n2491), .B1(ram[9510]), .B2(n2492), 
        .ZN(n13751) );
  MOAI22 U22665 ( .A1(n27534), .A2(n2491), .B1(ram[9511]), .B2(n2492), 
        .ZN(n13752) );
  MOAI22 U22666 ( .A1(n29179), .A2(n2493), .B1(ram[9512]), .B2(n2494), 
        .ZN(n13753) );
  MOAI22 U22667 ( .A1(n28944), .A2(n2493), .B1(ram[9513]), .B2(n2494), 
        .ZN(n13754) );
  MOAI22 U22668 ( .A1(n28709), .A2(n2493), .B1(ram[9514]), .B2(n2494), 
        .ZN(n13755) );
  MOAI22 U22669 ( .A1(n28474), .A2(n2493), .B1(ram[9515]), .B2(n2494), 
        .ZN(n13756) );
  MOAI22 U22670 ( .A1(n28239), .A2(n2493), .B1(ram[9516]), .B2(n2494), 
        .ZN(n13757) );
  MOAI22 U22671 ( .A1(n28004), .A2(n2493), .B1(ram[9517]), .B2(n2494), 
        .ZN(n13758) );
  MOAI22 U22672 ( .A1(n27769), .A2(n2493), .B1(ram[9518]), .B2(n2494), 
        .ZN(n13759) );
  MOAI22 U22673 ( .A1(n27534), .A2(n2493), .B1(ram[9519]), .B2(n2494), 
        .ZN(n13760) );
  MOAI22 U22674 ( .A1(n29179), .A2(n2495), .B1(ram[9520]), .B2(n2496), 
        .ZN(n13761) );
  MOAI22 U22675 ( .A1(n28944), .A2(n2495), .B1(ram[9521]), .B2(n2496), 
        .ZN(n13762) );
  MOAI22 U22676 ( .A1(n28709), .A2(n2495), .B1(ram[9522]), .B2(n2496), 
        .ZN(n13763) );
  MOAI22 U22677 ( .A1(n28474), .A2(n2495), .B1(ram[9523]), .B2(n2496), 
        .ZN(n13764) );
  MOAI22 U22678 ( .A1(n28239), .A2(n2495), .B1(ram[9524]), .B2(n2496), 
        .ZN(n13765) );
  MOAI22 U22679 ( .A1(n28004), .A2(n2495), .B1(ram[9525]), .B2(n2496), 
        .ZN(n13766) );
  MOAI22 U22680 ( .A1(n27769), .A2(n2495), .B1(ram[9526]), .B2(n2496), 
        .ZN(n13767) );
  MOAI22 U22681 ( .A1(n27534), .A2(n2495), .B1(ram[9527]), .B2(n2496), 
        .ZN(n13768) );
  MOAI22 U22682 ( .A1(n29179), .A2(n2497), .B1(ram[9528]), .B2(n2498), 
        .ZN(n13769) );
  MOAI22 U22683 ( .A1(n28944), .A2(n2497), .B1(ram[9529]), .B2(n2498), 
        .ZN(n13770) );
  MOAI22 U22684 ( .A1(n28709), .A2(n2497), .B1(ram[9530]), .B2(n2498), 
        .ZN(n13771) );
  MOAI22 U22685 ( .A1(n28474), .A2(n2497), .B1(ram[9531]), .B2(n2498), 
        .ZN(n13772) );
  MOAI22 U22686 ( .A1(n28239), .A2(n2497), .B1(ram[9532]), .B2(n2498), 
        .ZN(n13773) );
  MOAI22 U22687 ( .A1(n28004), .A2(n2497), .B1(ram[9533]), .B2(n2498), 
        .ZN(n13774) );
  MOAI22 U22688 ( .A1(n27769), .A2(n2497), .B1(ram[9534]), .B2(n2498), 
        .ZN(n13775) );
  MOAI22 U22689 ( .A1(n27534), .A2(n2497), .B1(ram[9535]), .B2(n2498), 
        .ZN(n13776) );
  MOAI22 U22690 ( .A1(n29179), .A2(n2499), .B1(ram[9536]), .B2(n2500), 
        .ZN(n13777) );
  MOAI22 U22691 ( .A1(n28944), .A2(n2499), .B1(ram[9537]), .B2(n2500), 
        .ZN(n13778) );
  MOAI22 U22692 ( .A1(n28709), .A2(n2499), .B1(ram[9538]), .B2(n2500), 
        .ZN(n13779) );
  MOAI22 U22693 ( .A1(n28474), .A2(n2499), .B1(ram[9539]), .B2(n2500), 
        .ZN(n13780) );
  MOAI22 U22694 ( .A1(n28239), .A2(n2499), .B1(ram[9540]), .B2(n2500), 
        .ZN(n13781) );
  MOAI22 U22695 ( .A1(n28004), .A2(n2499), .B1(ram[9541]), .B2(n2500), 
        .ZN(n13782) );
  MOAI22 U22696 ( .A1(n27769), .A2(n2499), .B1(ram[9542]), .B2(n2500), 
        .ZN(n13783) );
  MOAI22 U22697 ( .A1(n27534), .A2(n2499), .B1(ram[9543]), .B2(n2500), 
        .ZN(n13784) );
  MOAI22 U22698 ( .A1(n29179), .A2(n2501), .B1(ram[9544]), .B2(n2502), 
        .ZN(n13785) );
  MOAI22 U22699 ( .A1(n28944), .A2(n2501), .B1(ram[9545]), .B2(n2502), 
        .ZN(n13786) );
  MOAI22 U22700 ( .A1(n28709), .A2(n2501), .B1(ram[9546]), .B2(n2502), 
        .ZN(n13787) );
  MOAI22 U22701 ( .A1(n28474), .A2(n2501), .B1(ram[9547]), .B2(n2502), 
        .ZN(n13788) );
  MOAI22 U22702 ( .A1(n28239), .A2(n2501), .B1(ram[9548]), .B2(n2502), 
        .ZN(n13789) );
  MOAI22 U22703 ( .A1(n28004), .A2(n2501), .B1(ram[9549]), .B2(n2502), 
        .ZN(n13790) );
  MOAI22 U22704 ( .A1(n27769), .A2(n2501), .B1(ram[9550]), .B2(n2502), 
        .ZN(n13791) );
  MOAI22 U22705 ( .A1(n27534), .A2(n2501), .B1(ram[9551]), .B2(n2502), 
        .ZN(n13792) );
  MOAI22 U22706 ( .A1(n29179), .A2(n2503), .B1(ram[9552]), .B2(n2504), 
        .ZN(n13793) );
  MOAI22 U22707 ( .A1(n28944), .A2(n2503), .B1(ram[9553]), .B2(n2504), 
        .ZN(n13794) );
  MOAI22 U22708 ( .A1(n28709), .A2(n2503), .B1(ram[9554]), .B2(n2504), 
        .ZN(n13795) );
  MOAI22 U22709 ( .A1(n28474), .A2(n2503), .B1(ram[9555]), .B2(n2504), 
        .ZN(n13796) );
  MOAI22 U22710 ( .A1(n28239), .A2(n2503), .B1(ram[9556]), .B2(n2504), 
        .ZN(n13797) );
  MOAI22 U22711 ( .A1(n28004), .A2(n2503), .B1(ram[9557]), .B2(n2504), 
        .ZN(n13798) );
  MOAI22 U22712 ( .A1(n27769), .A2(n2503), .B1(ram[9558]), .B2(n2504), 
        .ZN(n13799) );
  MOAI22 U22713 ( .A1(n27534), .A2(n2503), .B1(ram[9559]), .B2(n2504), 
        .ZN(n13800) );
  MOAI22 U22714 ( .A1(n29179), .A2(n2505), .B1(ram[9560]), .B2(n2506), 
        .ZN(n13801) );
  MOAI22 U22715 ( .A1(n28944), .A2(n2505), .B1(ram[9561]), .B2(n2506), 
        .ZN(n13802) );
  MOAI22 U22716 ( .A1(n28709), .A2(n2505), .B1(ram[9562]), .B2(n2506), 
        .ZN(n13803) );
  MOAI22 U22717 ( .A1(n28474), .A2(n2505), .B1(ram[9563]), .B2(n2506), 
        .ZN(n13804) );
  MOAI22 U22718 ( .A1(n28239), .A2(n2505), .B1(ram[9564]), .B2(n2506), 
        .ZN(n13805) );
  MOAI22 U22719 ( .A1(n28004), .A2(n2505), .B1(ram[9565]), .B2(n2506), 
        .ZN(n13806) );
  MOAI22 U22720 ( .A1(n27769), .A2(n2505), .B1(ram[9566]), .B2(n2506), 
        .ZN(n13807) );
  MOAI22 U22721 ( .A1(n27534), .A2(n2505), .B1(ram[9567]), .B2(n2506), 
        .ZN(n13808) );
  MOAI22 U22722 ( .A1(n29180), .A2(n2507), .B1(ram[9568]), .B2(n2508), 
        .ZN(n13809) );
  MOAI22 U22723 ( .A1(n28945), .A2(n2507), .B1(ram[9569]), .B2(n2508), 
        .ZN(n13810) );
  MOAI22 U22724 ( .A1(n28710), .A2(n2507), .B1(ram[9570]), .B2(n2508), 
        .ZN(n13811) );
  MOAI22 U22725 ( .A1(n28475), .A2(n2507), .B1(ram[9571]), .B2(n2508), 
        .ZN(n13812) );
  MOAI22 U22726 ( .A1(n28240), .A2(n2507), .B1(ram[9572]), .B2(n2508), 
        .ZN(n13813) );
  MOAI22 U22727 ( .A1(n28005), .A2(n2507), .B1(ram[9573]), .B2(n2508), 
        .ZN(n13814) );
  MOAI22 U22728 ( .A1(n27770), .A2(n2507), .B1(ram[9574]), .B2(n2508), 
        .ZN(n13815) );
  MOAI22 U22729 ( .A1(n27535), .A2(n2507), .B1(ram[9575]), .B2(n2508), 
        .ZN(n13816) );
  MOAI22 U22730 ( .A1(n29180), .A2(n2509), .B1(ram[9576]), .B2(n2510), 
        .ZN(n13817) );
  MOAI22 U22731 ( .A1(n28945), .A2(n2509), .B1(ram[9577]), .B2(n2510), 
        .ZN(n13818) );
  MOAI22 U22732 ( .A1(n28710), .A2(n2509), .B1(ram[9578]), .B2(n2510), 
        .ZN(n13819) );
  MOAI22 U22733 ( .A1(n28475), .A2(n2509), .B1(ram[9579]), .B2(n2510), 
        .ZN(n13820) );
  MOAI22 U22734 ( .A1(n28240), .A2(n2509), .B1(ram[9580]), .B2(n2510), 
        .ZN(n13821) );
  MOAI22 U22735 ( .A1(n28005), .A2(n2509), .B1(ram[9581]), .B2(n2510), 
        .ZN(n13822) );
  MOAI22 U22736 ( .A1(n27770), .A2(n2509), .B1(ram[9582]), .B2(n2510), 
        .ZN(n13823) );
  MOAI22 U22737 ( .A1(n27535), .A2(n2509), .B1(ram[9583]), .B2(n2510), 
        .ZN(n13824) );
  MOAI22 U22738 ( .A1(n29180), .A2(n2511), .B1(ram[9584]), .B2(n2512), 
        .ZN(n13825) );
  MOAI22 U22739 ( .A1(n28945), .A2(n2511), .B1(ram[9585]), .B2(n2512), 
        .ZN(n13826) );
  MOAI22 U22740 ( .A1(n28710), .A2(n2511), .B1(ram[9586]), .B2(n2512), 
        .ZN(n13827) );
  MOAI22 U22741 ( .A1(n28475), .A2(n2511), .B1(ram[9587]), .B2(n2512), 
        .ZN(n13828) );
  MOAI22 U22742 ( .A1(n28240), .A2(n2511), .B1(ram[9588]), .B2(n2512), 
        .ZN(n13829) );
  MOAI22 U22743 ( .A1(n28005), .A2(n2511), .B1(ram[9589]), .B2(n2512), 
        .ZN(n13830) );
  MOAI22 U22744 ( .A1(n27770), .A2(n2511), .B1(ram[9590]), .B2(n2512), 
        .ZN(n13831) );
  MOAI22 U22745 ( .A1(n27535), .A2(n2511), .B1(ram[9591]), .B2(n2512), 
        .ZN(n13832) );
  MOAI22 U22746 ( .A1(n29180), .A2(n2513), .B1(ram[9592]), .B2(n2514), 
        .ZN(n13833) );
  MOAI22 U22747 ( .A1(n28945), .A2(n2513), .B1(ram[9593]), .B2(n2514), 
        .ZN(n13834) );
  MOAI22 U22748 ( .A1(n28710), .A2(n2513), .B1(ram[9594]), .B2(n2514), 
        .ZN(n13835) );
  MOAI22 U22749 ( .A1(n28475), .A2(n2513), .B1(ram[9595]), .B2(n2514), 
        .ZN(n13836) );
  MOAI22 U22750 ( .A1(n28240), .A2(n2513), .B1(ram[9596]), .B2(n2514), 
        .ZN(n13837) );
  MOAI22 U22751 ( .A1(n28005), .A2(n2513), .B1(ram[9597]), .B2(n2514), 
        .ZN(n13838) );
  MOAI22 U22752 ( .A1(n27770), .A2(n2513), .B1(ram[9598]), .B2(n2514), 
        .ZN(n13839) );
  MOAI22 U22753 ( .A1(n27535), .A2(n2513), .B1(ram[9599]), .B2(n2514), 
        .ZN(n13840) );
  MOAI22 U22754 ( .A1(n29180), .A2(n2515), .B1(ram[9600]), .B2(n2516), 
        .ZN(n13841) );
  MOAI22 U22755 ( .A1(n28945), .A2(n2515), .B1(ram[9601]), .B2(n2516), 
        .ZN(n13842) );
  MOAI22 U22756 ( .A1(n28710), .A2(n2515), .B1(ram[9602]), .B2(n2516), 
        .ZN(n13843) );
  MOAI22 U22757 ( .A1(n28475), .A2(n2515), .B1(ram[9603]), .B2(n2516), 
        .ZN(n13844) );
  MOAI22 U22758 ( .A1(n28240), .A2(n2515), .B1(ram[9604]), .B2(n2516), 
        .ZN(n13845) );
  MOAI22 U22759 ( .A1(n28005), .A2(n2515), .B1(ram[9605]), .B2(n2516), 
        .ZN(n13846) );
  MOAI22 U22760 ( .A1(n27770), .A2(n2515), .B1(ram[9606]), .B2(n2516), 
        .ZN(n13847) );
  MOAI22 U22761 ( .A1(n27535), .A2(n2515), .B1(ram[9607]), .B2(n2516), 
        .ZN(n13848) );
  MOAI22 U22762 ( .A1(n29180), .A2(n2517), .B1(ram[9608]), .B2(n2518), 
        .ZN(n13849) );
  MOAI22 U22763 ( .A1(n28945), .A2(n2517), .B1(ram[9609]), .B2(n2518), 
        .ZN(n13850) );
  MOAI22 U22764 ( .A1(n28710), .A2(n2517), .B1(ram[9610]), .B2(n2518), 
        .ZN(n13851) );
  MOAI22 U22765 ( .A1(n28475), .A2(n2517), .B1(ram[9611]), .B2(n2518), 
        .ZN(n13852) );
  MOAI22 U22766 ( .A1(n28240), .A2(n2517), .B1(ram[9612]), .B2(n2518), 
        .ZN(n13853) );
  MOAI22 U22767 ( .A1(n28005), .A2(n2517), .B1(ram[9613]), .B2(n2518), 
        .ZN(n13854) );
  MOAI22 U22768 ( .A1(n27770), .A2(n2517), .B1(ram[9614]), .B2(n2518), 
        .ZN(n13855) );
  MOAI22 U22769 ( .A1(n27535), .A2(n2517), .B1(ram[9615]), .B2(n2518), 
        .ZN(n13856) );
  MOAI22 U22770 ( .A1(n29180), .A2(n2519), .B1(ram[9616]), .B2(n2520), 
        .ZN(n13857) );
  MOAI22 U22771 ( .A1(n28945), .A2(n2519), .B1(ram[9617]), .B2(n2520), 
        .ZN(n13858) );
  MOAI22 U22772 ( .A1(n28710), .A2(n2519), .B1(ram[9618]), .B2(n2520), 
        .ZN(n13859) );
  MOAI22 U22773 ( .A1(n28475), .A2(n2519), .B1(ram[9619]), .B2(n2520), 
        .ZN(n13860) );
  MOAI22 U22774 ( .A1(n28240), .A2(n2519), .B1(ram[9620]), .B2(n2520), 
        .ZN(n13861) );
  MOAI22 U22775 ( .A1(n28005), .A2(n2519), .B1(ram[9621]), .B2(n2520), 
        .ZN(n13862) );
  MOAI22 U22776 ( .A1(n27770), .A2(n2519), .B1(ram[9622]), .B2(n2520), 
        .ZN(n13863) );
  MOAI22 U22777 ( .A1(n27535), .A2(n2519), .B1(ram[9623]), .B2(n2520), 
        .ZN(n13864) );
  MOAI22 U22778 ( .A1(n29180), .A2(n2521), .B1(ram[9624]), .B2(n2522), 
        .ZN(n13865) );
  MOAI22 U22779 ( .A1(n28945), .A2(n2521), .B1(ram[9625]), .B2(n2522), 
        .ZN(n13866) );
  MOAI22 U22780 ( .A1(n28710), .A2(n2521), .B1(ram[9626]), .B2(n2522), 
        .ZN(n13867) );
  MOAI22 U22781 ( .A1(n28475), .A2(n2521), .B1(ram[9627]), .B2(n2522), 
        .ZN(n13868) );
  MOAI22 U22782 ( .A1(n28240), .A2(n2521), .B1(ram[9628]), .B2(n2522), 
        .ZN(n13869) );
  MOAI22 U22783 ( .A1(n28005), .A2(n2521), .B1(ram[9629]), .B2(n2522), 
        .ZN(n13870) );
  MOAI22 U22784 ( .A1(n27770), .A2(n2521), .B1(ram[9630]), .B2(n2522), 
        .ZN(n13871) );
  MOAI22 U22785 ( .A1(n27535), .A2(n2521), .B1(ram[9631]), .B2(n2522), 
        .ZN(n13872) );
  MOAI22 U22786 ( .A1(n29180), .A2(n2523), .B1(ram[9632]), .B2(n2524), 
        .ZN(n13873) );
  MOAI22 U22787 ( .A1(n28945), .A2(n2523), .B1(ram[9633]), .B2(n2524), 
        .ZN(n13874) );
  MOAI22 U22788 ( .A1(n28710), .A2(n2523), .B1(ram[9634]), .B2(n2524), 
        .ZN(n13875) );
  MOAI22 U22789 ( .A1(n28475), .A2(n2523), .B1(ram[9635]), .B2(n2524), 
        .ZN(n13876) );
  MOAI22 U22790 ( .A1(n28240), .A2(n2523), .B1(ram[9636]), .B2(n2524), 
        .ZN(n13877) );
  MOAI22 U22791 ( .A1(n28005), .A2(n2523), .B1(ram[9637]), .B2(n2524), 
        .ZN(n13878) );
  MOAI22 U22792 ( .A1(n27770), .A2(n2523), .B1(ram[9638]), .B2(n2524), 
        .ZN(n13879) );
  MOAI22 U22793 ( .A1(n27535), .A2(n2523), .B1(ram[9639]), .B2(n2524), 
        .ZN(n13880) );
  MOAI22 U22794 ( .A1(n29180), .A2(n2525), .B1(ram[9640]), .B2(n2526), 
        .ZN(n13881) );
  MOAI22 U22795 ( .A1(n28945), .A2(n2525), .B1(ram[9641]), .B2(n2526), 
        .ZN(n13882) );
  MOAI22 U22796 ( .A1(n28710), .A2(n2525), .B1(ram[9642]), .B2(n2526), 
        .ZN(n13883) );
  MOAI22 U22797 ( .A1(n28475), .A2(n2525), .B1(ram[9643]), .B2(n2526), 
        .ZN(n13884) );
  MOAI22 U22798 ( .A1(n28240), .A2(n2525), .B1(ram[9644]), .B2(n2526), 
        .ZN(n13885) );
  MOAI22 U22799 ( .A1(n28005), .A2(n2525), .B1(ram[9645]), .B2(n2526), 
        .ZN(n13886) );
  MOAI22 U22800 ( .A1(n27770), .A2(n2525), .B1(ram[9646]), .B2(n2526), 
        .ZN(n13887) );
  MOAI22 U22801 ( .A1(n27535), .A2(n2525), .B1(ram[9647]), .B2(n2526), 
        .ZN(n13888) );
  MOAI22 U22802 ( .A1(n29180), .A2(n2527), .B1(ram[9648]), .B2(n2528), 
        .ZN(n13889) );
  MOAI22 U22803 ( .A1(n28945), .A2(n2527), .B1(ram[9649]), .B2(n2528), 
        .ZN(n13890) );
  MOAI22 U22804 ( .A1(n28710), .A2(n2527), .B1(ram[9650]), .B2(n2528), 
        .ZN(n13891) );
  MOAI22 U22805 ( .A1(n28475), .A2(n2527), .B1(ram[9651]), .B2(n2528), 
        .ZN(n13892) );
  MOAI22 U22806 ( .A1(n28240), .A2(n2527), .B1(ram[9652]), .B2(n2528), 
        .ZN(n13893) );
  MOAI22 U22807 ( .A1(n28005), .A2(n2527), .B1(ram[9653]), .B2(n2528), 
        .ZN(n13894) );
  MOAI22 U22808 ( .A1(n27770), .A2(n2527), .B1(ram[9654]), .B2(n2528), 
        .ZN(n13895) );
  MOAI22 U22809 ( .A1(n27535), .A2(n2527), .B1(ram[9655]), .B2(n2528), 
        .ZN(n13896) );
  MOAI22 U22810 ( .A1(n29180), .A2(n2529), .B1(ram[9656]), .B2(n2530), 
        .ZN(n13897) );
  MOAI22 U22811 ( .A1(n28945), .A2(n2529), .B1(ram[9657]), .B2(n2530), 
        .ZN(n13898) );
  MOAI22 U22812 ( .A1(n28710), .A2(n2529), .B1(ram[9658]), .B2(n2530), 
        .ZN(n13899) );
  MOAI22 U22813 ( .A1(n28475), .A2(n2529), .B1(ram[9659]), .B2(n2530), 
        .ZN(n13900) );
  MOAI22 U22814 ( .A1(n28240), .A2(n2529), .B1(ram[9660]), .B2(n2530), 
        .ZN(n13901) );
  MOAI22 U22815 ( .A1(n28005), .A2(n2529), .B1(ram[9661]), .B2(n2530), 
        .ZN(n13902) );
  MOAI22 U22816 ( .A1(n27770), .A2(n2529), .B1(ram[9662]), .B2(n2530), 
        .ZN(n13903) );
  MOAI22 U22817 ( .A1(n27535), .A2(n2529), .B1(ram[9663]), .B2(n2530), 
        .ZN(n13904) );
  MOAI22 U22818 ( .A1(n29180), .A2(n2531), .B1(ram[9664]), .B2(n2532), 
        .ZN(n13905) );
  MOAI22 U22819 ( .A1(n28945), .A2(n2531), .B1(ram[9665]), .B2(n2532), 
        .ZN(n13906) );
  MOAI22 U22820 ( .A1(n28710), .A2(n2531), .B1(ram[9666]), .B2(n2532), 
        .ZN(n13907) );
  MOAI22 U22821 ( .A1(n28475), .A2(n2531), .B1(ram[9667]), .B2(n2532), 
        .ZN(n13908) );
  MOAI22 U22822 ( .A1(n28240), .A2(n2531), .B1(ram[9668]), .B2(n2532), 
        .ZN(n13909) );
  MOAI22 U22823 ( .A1(n28005), .A2(n2531), .B1(ram[9669]), .B2(n2532), 
        .ZN(n13910) );
  MOAI22 U22824 ( .A1(n27770), .A2(n2531), .B1(ram[9670]), .B2(n2532), 
        .ZN(n13911) );
  MOAI22 U22825 ( .A1(n27535), .A2(n2531), .B1(ram[9671]), .B2(n2532), 
        .ZN(n13912) );
  MOAI22 U22826 ( .A1(n29181), .A2(n2533), .B1(ram[9672]), .B2(n2534), 
        .ZN(n13913) );
  MOAI22 U22827 ( .A1(n28946), .A2(n2533), .B1(ram[9673]), .B2(n2534), 
        .ZN(n13914) );
  MOAI22 U22828 ( .A1(n28711), .A2(n2533), .B1(ram[9674]), .B2(n2534), 
        .ZN(n13915) );
  MOAI22 U22829 ( .A1(n28476), .A2(n2533), .B1(ram[9675]), .B2(n2534), 
        .ZN(n13916) );
  MOAI22 U22830 ( .A1(n28241), .A2(n2533), .B1(ram[9676]), .B2(n2534), 
        .ZN(n13917) );
  MOAI22 U22831 ( .A1(n28006), .A2(n2533), .B1(ram[9677]), .B2(n2534), 
        .ZN(n13918) );
  MOAI22 U22832 ( .A1(n27771), .A2(n2533), .B1(ram[9678]), .B2(n2534), 
        .ZN(n13919) );
  MOAI22 U22833 ( .A1(n27536), .A2(n2533), .B1(ram[9679]), .B2(n2534), 
        .ZN(n13920) );
  MOAI22 U22834 ( .A1(n29181), .A2(n2535), .B1(ram[9680]), .B2(n2536), 
        .ZN(n13921) );
  MOAI22 U22835 ( .A1(n28946), .A2(n2535), .B1(ram[9681]), .B2(n2536), 
        .ZN(n13922) );
  MOAI22 U22836 ( .A1(n28711), .A2(n2535), .B1(ram[9682]), .B2(n2536), 
        .ZN(n13923) );
  MOAI22 U22837 ( .A1(n28476), .A2(n2535), .B1(ram[9683]), .B2(n2536), 
        .ZN(n13924) );
  MOAI22 U22838 ( .A1(n28241), .A2(n2535), .B1(ram[9684]), .B2(n2536), 
        .ZN(n13925) );
  MOAI22 U22839 ( .A1(n28006), .A2(n2535), .B1(ram[9685]), .B2(n2536), 
        .ZN(n13926) );
  MOAI22 U22840 ( .A1(n27771), .A2(n2535), .B1(ram[9686]), .B2(n2536), 
        .ZN(n13927) );
  MOAI22 U22841 ( .A1(n27536), .A2(n2535), .B1(ram[9687]), .B2(n2536), 
        .ZN(n13928) );
  MOAI22 U22842 ( .A1(n29181), .A2(n2537), .B1(ram[9688]), .B2(n2538), 
        .ZN(n13929) );
  MOAI22 U22843 ( .A1(n28946), .A2(n2537), .B1(ram[9689]), .B2(n2538), 
        .ZN(n13930) );
  MOAI22 U22844 ( .A1(n28711), .A2(n2537), .B1(ram[9690]), .B2(n2538), 
        .ZN(n13931) );
  MOAI22 U22845 ( .A1(n28476), .A2(n2537), .B1(ram[9691]), .B2(n2538), 
        .ZN(n13932) );
  MOAI22 U22846 ( .A1(n28241), .A2(n2537), .B1(ram[9692]), .B2(n2538), 
        .ZN(n13933) );
  MOAI22 U22847 ( .A1(n28006), .A2(n2537), .B1(ram[9693]), .B2(n2538), 
        .ZN(n13934) );
  MOAI22 U22848 ( .A1(n27771), .A2(n2537), .B1(ram[9694]), .B2(n2538), 
        .ZN(n13935) );
  MOAI22 U22849 ( .A1(n27536), .A2(n2537), .B1(ram[9695]), .B2(n2538), 
        .ZN(n13936) );
  MOAI22 U22850 ( .A1(n29181), .A2(n2539), .B1(ram[9696]), .B2(n2540), 
        .ZN(n13937) );
  MOAI22 U22851 ( .A1(n28946), .A2(n2539), .B1(ram[9697]), .B2(n2540), 
        .ZN(n13938) );
  MOAI22 U22852 ( .A1(n28711), .A2(n2539), .B1(ram[9698]), .B2(n2540), 
        .ZN(n13939) );
  MOAI22 U22853 ( .A1(n28476), .A2(n2539), .B1(ram[9699]), .B2(n2540), 
        .ZN(n13940) );
  MOAI22 U22854 ( .A1(n28241), .A2(n2539), .B1(ram[9700]), .B2(n2540), 
        .ZN(n13941) );
  MOAI22 U22855 ( .A1(n28006), .A2(n2539), .B1(ram[9701]), .B2(n2540), 
        .ZN(n13942) );
  MOAI22 U22856 ( .A1(n27771), .A2(n2539), .B1(ram[9702]), .B2(n2540), 
        .ZN(n13943) );
  MOAI22 U22857 ( .A1(n27536), .A2(n2539), .B1(ram[9703]), .B2(n2540), 
        .ZN(n13944) );
  MOAI22 U22858 ( .A1(n29181), .A2(n2541), .B1(ram[9704]), .B2(n2542), 
        .ZN(n13945) );
  MOAI22 U22859 ( .A1(n28946), .A2(n2541), .B1(ram[9705]), .B2(n2542), 
        .ZN(n13946) );
  MOAI22 U22860 ( .A1(n28711), .A2(n2541), .B1(ram[9706]), .B2(n2542), 
        .ZN(n13947) );
  MOAI22 U22861 ( .A1(n28476), .A2(n2541), .B1(ram[9707]), .B2(n2542), 
        .ZN(n13948) );
  MOAI22 U22862 ( .A1(n28241), .A2(n2541), .B1(ram[9708]), .B2(n2542), 
        .ZN(n13949) );
  MOAI22 U22863 ( .A1(n28006), .A2(n2541), .B1(ram[9709]), .B2(n2542), 
        .ZN(n13950) );
  MOAI22 U22864 ( .A1(n27771), .A2(n2541), .B1(ram[9710]), .B2(n2542), 
        .ZN(n13951) );
  MOAI22 U22865 ( .A1(n27536), .A2(n2541), .B1(ram[9711]), .B2(n2542), 
        .ZN(n13952) );
  MOAI22 U22866 ( .A1(n29181), .A2(n2543), .B1(ram[9712]), .B2(n2544), 
        .ZN(n13953) );
  MOAI22 U22867 ( .A1(n28946), .A2(n2543), .B1(ram[9713]), .B2(n2544), 
        .ZN(n13954) );
  MOAI22 U22868 ( .A1(n28711), .A2(n2543), .B1(ram[9714]), .B2(n2544), 
        .ZN(n13955) );
  MOAI22 U22869 ( .A1(n28476), .A2(n2543), .B1(ram[9715]), .B2(n2544), 
        .ZN(n13956) );
  MOAI22 U22870 ( .A1(n28241), .A2(n2543), .B1(ram[9716]), .B2(n2544), 
        .ZN(n13957) );
  MOAI22 U22871 ( .A1(n28006), .A2(n2543), .B1(ram[9717]), .B2(n2544), 
        .ZN(n13958) );
  MOAI22 U22872 ( .A1(n27771), .A2(n2543), .B1(ram[9718]), .B2(n2544), 
        .ZN(n13959) );
  MOAI22 U22873 ( .A1(n27536), .A2(n2543), .B1(ram[9719]), .B2(n2544), 
        .ZN(n13960) );
  MOAI22 U22874 ( .A1(n29181), .A2(n2545), .B1(ram[9720]), .B2(n2546), 
        .ZN(n13961) );
  MOAI22 U22875 ( .A1(n28946), .A2(n2545), .B1(ram[9721]), .B2(n2546), 
        .ZN(n13962) );
  MOAI22 U22876 ( .A1(n28711), .A2(n2545), .B1(ram[9722]), .B2(n2546), 
        .ZN(n13963) );
  MOAI22 U22877 ( .A1(n28476), .A2(n2545), .B1(ram[9723]), .B2(n2546), 
        .ZN(n13964) );
  MOAI22 U22878 ( .A1(n28241), .A2(n2545), .B1(ram[9724]), .B2(n2546), 
        .ZN(n13965) );
  MOAI22 U22879 ( .A1(n28006), .A2(n2545), .B1(ram[9725]), .B2(n2546), 
        .ZN(n13966) );
  MOAI22 U22880 ( .A1(n27771), .A2(n2545), .B1(ram[9726]), .B2(n2546), 
        .ZN(n13967) );
  MOAI22 U22881 ( .A1(n27536), .A2(n2545), .B1(ram[9727]), .B2(n2546), 
        .ZN(n13968) );
  MOAI22 U22882 ( .A1(n29181), .A2(n2547), .B1(ram[9728]), .B2(n2548), 
        .ZN(n13969) );
  MOAI22 U22883 ( .A1(n28946), .A2(n2547), .B1(ram[9729]), .B2(n2548), 
        .ZN(n13970) );
  MOAI22 U22884 ( .A1(n28711), .A2(n2547), .B1(ram[9730]), .B2(n2548), 
        .ZN(n13971) );
  MOAI22 U22885 ( .A1(n28476), .A2(n2547), .B1(ram[9731]), .B2(n2548), 
        .ZN(n13972) );
  MOAI22 U22886 ( .A1(n28241), .A2(n2547), .B1(ram[9732]), .B2(n2548), 
        .ZN(n13973) );
  MOAI22 U22887 ( .A1(n28006), .A2(n2547), .B1(ram[9733]), .B2(n2548), 
        .ZN(n13974) );
  MOAI22 U22888 ( .A1(n27771), .A2(n2547), .B1(ram[9734]), .B2(n2548), 
        .ZN(n13975) );
  MOAI22 U22889 ( .A1(n27536), .A2(n2547), .B1(ram[9735]), .B2(n2548), 
        .ZN(n13976) );
  MOAI22 U22890 ( .A1(n29181), .A2(n2550), .B1(ram[9736]), .B2(n2551), 
        .ZN(n13977) );
  MOAI22 U22891 ( .A1(n28946), .A2(n2550), .B1(ram[9737]), .B2(n2551), 
        .ZN(n13978) );
  MOAI22 U22892 ( .A1(n28711), .A2(n2550), .B1(ram[9738]), .B2(n2551), 
        .ZN(n13979) );
  MOAI22 U22893 ( .A1(n28476), .A2(n2550), .B1(ram[9739]), .B2(n2551), 
        .ZN(n13980) );
  MOAI22 U22894 ( .A1(n28241), .A2(n2550), .B1(ram[9740]), .B2(n2551), 
        .ZN(n13981) );
  MOAI22 U22895 ( .A1(n28006), .A2(n2550), .B1(ram[9741]), .B2(n2551), 
        .ZN(n13982) );
  MOAI22 U22896 ( .A1(n27771), .A2(n2550), .B1(ram[9742]), .B2(n2551), 
        .ZN(n13983) );
  MOAI22 U22897 ( .A1(n27536), .A2(n2550), .B1(ram[9743]), .B2(n2551), 
        .ZN(n13984) );
  MOAI22 U22898 ( .A1(n29181), .A2(n2552), .B1(ram[9744]), .B2(n2553), 
        .ZN(n13985) );
  MOAI22 U22899 ( .A1(n28946), .A2(n2552), .B1(ram[9745]), .B2(n2553), 
        .ZN(n13986) );
  MOAI22 U22900 ( .A1(n28711), .A2(n2552), .B1(ram[9746]), .B2(n2553), 
        .ZN(n13987) );
  MOAI22 U22901 ( .A1(n28476), .A2(n2552), .B1(ram[9747]), .B2(n2553), 
        .ZN(n13988) );
  MOAI22 U22902 ( .A1(n28241), .A2(n2552), .B1(ram[9748]), .B2(n2553), 
        .ZN(n13989) );
  MOAI22 U22903 ( .A1(n28006), .A2(n2552), .B1(ram[9749]), .B2(n2553), 
        .ZN(n13990) );
  MOAI22 U22904 ( .A1(n27771), .A2(n2552), .B1(ram[9750]), .B2(n2553), 
        .ZN(n13991) );
  MOAI22 U22905 ( .A1(n27536), .A2(n2552), .B1(ram[9751]), .B2(n2553), 
        .ZN(n13992) );
  MOAI22 U22906 ( .A1(n29181), .A2(n2554), .B1(ram[9752]), .B2(n2555), 
        .ZN(n13993) );
  MOAI22 U22907 ( .A1(n28946), .A2(n2554), .B1(ram[9753]), .B2(n2555), 
        .ZN(n13994) );
  MOAI22 U22908 ( .A1(n28711), .A2(n2554), .B1(ram[9754]), .B2(n2555), 
        .ZN(n13995) );
  MOAI22 U22909 ( .A1(n28476), .A2(n2554), .B1(ram[9755]), .B2(n2555), 
        .ZN(n13996) );
  MOAI22 U22910 ( .A1(n28241), .A2(n2554), .B1(ram[9756]), .B2(n2555), 
        .ZN(n13997) );
  MOAI22 U22911 ( .A1(n28006), .A2(n2554), .B1(ram[9757]), .B2(n2555), 
        .ZN(n13998) );
  MOAI22 U22912 ( .A1(n27771), .A2(n2554), .B1(ram[9758]), .B2(n2555), 
        .ZN(n13999) );
  MOAI22 U22913 ( .A1(n27536), .A2(n2554), .B1(ram[9759]), .B2(n2555), 
        .ZN(n14000) );
  MOAI22 U22914 ( .A1(n29181), .A2(n2556), .B1(ram[9760]), .B2(n2557), 
        .ZN(n14001) );
  MOAI22 U22915 ( .A1(n28946), .A2(n2556), .B1(ram[9761]), .B2(n2557), 
        .ZN(n14002) );
  MOAI22 U22916 ( .A1(n28711), .A2(n2556), .B1(ram[9762]), .B2(n2557), 
        .ZN(n14003) );
  MOAI22 U22917 ( .A1(n28476), .A2(n2556), .B1(ram[9763]), .B2(n2557), 
        .ZN(n14004) );
  MOAI22 U22918 ( .A1(n28241), .A2(n2556), .B1(ram[9764]), .B2(n2557), 
        .ZN(n14005) );
  MOAI22 U22919 ( .A1(n28006), .A2(n2556), .B1(ram[9765]), .B2(n2557), 
        .ZN(n14006) );
  MOAI22 U22920 ( .A1(n27771), .A2(n2556), .B1(ram[9766]), .B2(n2557), 
        .ZN(n14007) );
  MOAI22 U22921 ( .A1(n27536), .A2(n2556), .B1(ram[9767]), .B2(n2557), 
        .ZN(n14008) );
  MOAI22 U22922 ( .A1(n29181), .A2(n2558), .B1(ram[9768]), .B2(n2559), 
        .ZN(n14009) );
  MOAI22 U22923 ( .A1(n28946), .A2(n2558), .B1(ram[9769]), .B2(n2559), 
        .ZN(n14010) );
  MOAI22 U22924 ( .A1(n28711), .A2(n2558), .B1(ram[9770]), .B2(n2559), 
        .ZN(n14011) );
  MOAI22 U22925 ( .A1(n28476), .A2(n2558), .B1(ram[9771]), .B2(n2559), 
        .ZN(n14012) );
  MOAI22 U22926 ( .A1(n28241), .A2(n2558), .B1(ram[9772]), .B2(n2559), 
        .ZN(n14013) );
  MOAI22 U22927 ( .A1(n28006), .A2(n2558), .B1(ram[9773]), .B2(n2559), 
        .ZN(n14014) );
  MOAI22 U22928 ( .A1(n27771), .A2(n2558), .B1(ram[9774]), .B2(n2559), 
        .ZN(n14015) );
  MOAI22 U22929 ( .A1(n27536), .A2(n2558), .B1(ram[9775]), .B2(n2559), 
        .ZN(n14016) );
  MOAI22 U22930 ( .A1(n29182), .A2(n2560), .B1(ram[9776]), .B2(n2561), 
        .ZN(n14017) );
  MOAI22 U22931 ( .A1(n28947), .A2(n2560), .B1(ram[9777]), .B2(n2561), 
        .ZN(n14018) );
  MOAI22 U22932 ( .A1(n28712), .A2(n2560), .B1(ram[9778]), .B2(n2561), 
        .ZN(n14019) );
  MOAI22 U22933 ( .A1(n28477), .A2(n2560), .B1(ram[9779]), .B2(n2561), 
        .ZN(n14020) );
  MOAI22 U22934 ( .A1(n28242), .A2(n2560), .B1(ram[9780]), .B2(n2561), 
        .ZN(n14021) );
  MOAI22 U22935 ( .A1(n28007), .A2(n2560), .B1(ram[9781]), .B2(n2561), 
        .ZN(n14022) );
  MOAI22 U22936 ( .A1(n27772), .A2(n2560), .B1(ram[9782]), .B2(n2561), 
        .ZN(n14023) );
  MOAI22 U22937 ( .A1(n27537), .A2(n2560), .B1(ram[9783]), .B2(n2561), 
        .ZN(n14024) );
  MOAI22 U22938 ( .A1(n29182), .A2(n2562), .B1(ram[9784]), .B2(n2563), 
        .ZN(n14025) );
  MOAI22 U22939 ( .A1(n28947), .A2(n2562), .B1(ram[9785]), .B2(n2563), 
        .ZN(n14026) );
  MOAI22 U22940 ( .A1(n28712), .A2(n2562), .B1(ram[9786]), .B2(n2563), 
        .ZN(n14027) );
  MOAI22 U22941 ( .A1(n28477), .A2(n2562), .B1(ram[9787]), .B2(n2563), 
        .ZN(n14028) );
  MOAI22 U22942 ( .A1(n28242), .A2(n2562), .B1(ram[9788]), .B2(n2563), 
        .ZN(n14029) );
  MOAI22 U22943 ( .A1(n28007), .A2(n2562), .B1(ram[9789]), .B2(n2563), 
        .ZN(n14030) );
  MOAI22 U22944 ( .A1(n27772), .A2(n2562), .B1(ram[9790]), .B2(n2563), 
        .ZN(n14031) );
  MOAI22 U22945 ( .A1(n27537), .A2(n2562), .B1(ram[9791]), .B2(n2563), 
        .ZN(n14032) );
  MOAI22 U22946 ( .A1(n29182), .A2(n2564), .B1(ram[9792]), .B2(n2565), 
        .ZN(n14033) );
  MOAI22 U22947 ( .A1(n28947), .A2(n2564), .B1(ram[9793]), .B2(n2565), 
        .ZN(n14034) );
  MOAI22 U22948 ( .A1(n28712), .A2(n2564), .B1(ram[9794]), .B2(n2565), 
        .ZN(n14035) );
  MOAI22 U22949 ( .A1(n28477), .A2(n2564), .B1(ram[9795]), .B2(n2565), 
        .ZN(n14036) );
  MOAI22 U22950 ( .A1(n28242), .A2(n2564), .B1(ram[9796]), .B2(n2565), 
        .ZN(n14037) );
  MOAI22 U22951 ( .A1(n28007), .A2(n2564), .B1(ram[9797]), .B2(n2565), 
        .ZN(n14038) );
  MOAI22 U22952 ( .A1(n27772), .A2(n2564), .B1(ram[9798]), .B2(n2565), 
        .ZN(n14039) );
  MOAI22 U22953 ( .A1(n27537), .A2(n2564), .B1(ram[9799]), .B2(n2565), 
        .ZN(n14040) );
  MOAI22 U22954 ( .A1(n29182), .A2(n2566), .B1(ram[9800]), .B2(n2567), 
        .ZN(n14041) );
  MOAI22 U22955 ( .A1(n28947), .A2(n2566), .B1(ram[9801]), .B2(n2567), 
        .ZN(n14042) );
  MOAI22 U22956 ( .A1(n28712), .A2(n2566), .B1(ram[9802]), .B2(n2567), 
        .ZN(n14043) );
  MOAI22 U22957 ( .A1(n28477), .A2(n2566), .B1(ram[9803]), .B2(n2567), 
        .ZN(n14044) );
  MOAI22 U22958 ( .A1(n28242), .A2(n2566), .B1(ram[9804]), .B2(n2567), 
        .ZN(n14045) );
  MOAI22 U22959 ( .A1(n28007), .A2(n2566), .B1(ram[9805]), .B2(n2567), 
        .ZN(n14046) );
  MOAI22 U22960 ( .A1(n27772), .A2(n2566), .B1(ram[9806]), .B2(n2567), 
        .ZN(n14047) );
  MOAI22 U22961 ( .A1(n27537), .A2(n2566), .B1(ram[9807]), .B2(n2567), 
        .ZN(n14048) );
  MOAI22 U22962 ( .A1(n29182), .A2(n2568), .B1(ram[9808]), .B2(n2569), 
        .ZN(n14049) );
  MOAI22 U22963 ( .A1(n28947), .A2(n2568), .B1(ram[9809]), .B2(n2569), 
        .ZN(n14050) );
  MOAI22 U22964 ( .A1(n28712), .A2(n2568), .B1(ram[9810]), .B2(n2569), 
        .ZN(n14051) );
  MOAI22 U22965 ( .A1(n28477), .A2(n2568), .B1(ram[9811]), .B2(n2569), 
        .ZN(n14052) );
  MOAI22 U22966 ( .A1(n28242), .A2(n2568), .B1(ram[9812]), .B2(n2569), 
        .ZN(n14053) );
  MOAI22 U22967 ( .A1(n28007), .A2(n2568), .B1(ram[9813]), .B2(n2569), 
        .ZN(n14054) );
  MOAI22 U22968 ( .A1(n27772), .A2(n2568), .B1(ram[9814]), .B2(n2569), 
        .ZN(n14055) );
  MOAI22 U22969 ( .A1(n27537), .A2(n2568), .B1(ram[9815]), .B2(n2569), 
        .ZN(n14056) );
  MOAI22 U22970 ( .A1(n29182), .A2(n2570), .B1(ram[9816]), .B2(n2571), 
        .ZN(n14057) );
  MOAI22 U22971 ( .A1(n28947), .A2(n2570), .B1(ram[9817]), .B2(n2571), 
        .ZN(n14058) );
  MOAI22 U22972 ( .A1(n28712), .A2(n2570), .B1(ram[9818]), .B2(n2571), 
        .ZN(n14059) );
  MOAI22 U22973 ( .A1(n28477), .A2(n2570), .B1(ram[9819]), .B2(n2571), 
        .ZN(n14060) );
  MOAI22 U22974 ( .A1(n28242), .A2(n2570), .B1(ram[9820]), .B2(n2571), 
        .ZN(n14061) );
  MOAI22 U22975 ( .A1(n28007), .A2(n2570), .B1(ram[9821]), .B2(n2571), 
        .ZN(n14062) );
  MOAI22 U22976 ( .A1(n27772), .A2(n2570), .B1(ram[9822]), .B2(n2571), 
        .ZN(n14063) );
  MOAI22 U22977 ( .A1(n27537), .A2(n2570), .B1(ram[9823]), .B2(n2571), 
        .ZN(n14064) );
  MOAI22 U22978 ( .A1(n29182), .A2(n2572), .B1(ram[9824]), .B2(n2573), 
        .ZN(n14065) );
  MOAI22 U22979 ( .A1(n28947), .A2(n2572), .B1(ram[9825]), .B2(n2573), 
        .ZN(n14066) );
  MOAI22 U22980 ( .A1(n28712), .A2(n2572), .B1(ram[9826]), .B2(n2573), 
        .ZN(n14067) );
  MOAI22 U22981 ( .A1(n28477), .A2(n2572), .B1(ram[9827]), .B2(n2573), 
        .ZN(n14068) );
  MOAI22 U22982 ( .A1(n28242), .A2(n2572), .B1(ram[9828]), .B2(n2573), 
        .ZN(n14069) );
  MOAI22 U22983 ( .A1(n28007), .A2(n2572), .B1(ram[9829]), .B2(n2573), 
        .ZN(n14070) );
  MOAI22 U22984 ( .A1(n27772), .A2(n2572), .B1(ram[9830]), .B2(n2573), 
        .ZN(n14071) );
  MOAI22 U22985 ( .A1(n27537), .A2(n2572), .B1(ram[9831]), .B2(n2573), 
        .ZN(n14072) );
  MOAI22 U22986 ( .A1(n29182), .A2(n2574), .B1(ram[9832]), .B2(n2575), 
        .ZN(n14073) );
  MOAI22 U22987 ( .A1(n28947), .A2(n2574), .B1(ram[9833]), .B2(n2575), 
        .ZN(n14074) );
  MOAI22 U22988 ( .A1(n28712), .A2(n2574), .B1(ram[9834]), .B2(n2575), 
        .ZN(n14075) );
  MOAI22 U22989 ( .A1(n28477), .A2(n2574), .B1(ram[9835]), .B2(n2575), 
        .ZN(n14076) );
  MOAI22 U22990 ( .A1(n28242), .A2(n2574), .B1(ram[9836]), .B2(n2575), 
        .ZN(n14077) );
  MOAI22 U22991 ( .A1(n28007), .A2(n2574), .B1(ram[9837]), .B2(n2575), 
        .ZN(n14078) );
  MOAI22 U22992 ( .A1(n27772), .A2(n2574), .B1(ram[9838]), .B2(n2575), 
        .ZN(n14079) );
  MOAI22 U22993 ( .A1(n27537), .A2(n2574), .B1(ram[9839]), .B2(n2575), 
        .ZN(n14080) );
  MOAI22 U22994 ( .A1(n29182), .A2(n2576), .B1(ram[9840]), .B2(n2577), 
        .ZN(n14081) );
  MOAI22 U22995 ( .A1(n28947), .A2(n2576), .B1(ram[9841]), .B2(n2577), 
        .ZN(n14082) );
  MOAI22 U22996 ( .A1(n28712), .A2(n2576), .B1(ram[9842]), .B2(n2577), 
        .ZN(n14083) );
  MOAI22 U22997 ( .A1(n28477), .A2(n2576), .B1(ram[9843]), .B2(n2577), 
        .ZN(n14084) );
  MOAI22 U22998 ( .A1(n28242), .A2(n2576), .B1(ram[9844]), .B2(n2577), 
        .ZN(n14085) );
  MOAI22 U22999 ( .A1(n28007), .A2(n2576), .B1(ram[9845]), .B2(n2577), 
        .ZN(n14086) );
  MOAI22 U23000 ( .A1(n27772), .A2(n2576), .B1(ram[9846]), .B2(n2577), 
        .ZN(n14087) );
  MOAI22 U23001 ( .A1(n27537), .A2(n2576), .B1(ram[9847]), .B2(n2577), 
        .ZN(n14088) );
  MOAI22 U23002 ( .A1(n29182), .A2(n2578), .B1(ram[9848]), .B2(n2579), 
        .ZN(n14089) );
  MOAI22 U23003 ( .A1(n28947), .A2(n2578), .B1(ram[9849]), .B2(n2579), 
        .ZN(n14090) );
  MOAI22 U23004 ( .A1(n28712), .A2(n2578), .B1(ram[9850]), .B2(n2579), 
        .ZN(n14091) );
  MOAI22 U23005 ( .A1(n28477), .A2(n2578), .B1(ram[9851]), .B2(n2579), 
        .ZN(n14092) );
  MOAI22 U23006 ( .A1(n28242), .A2(n2578), .B1(ram[9852]), .B2(n2579), 
        .ZN(n14093) );
  MOAI22 U23007 ( .A1(n28007), .A2(n2578), .B1(ram[9853]), .B2(n2579), 
        .ZN(n14094) );
  MOAI22 U23008 ( .A1(n27772), .A2(n2578), .B1(ram[9854]), .B2(n2579), 
        .ZN(n14095) );
  MOAI22 U23009 ( .A1(n27537), .A2(n2578), .B1(ram[9855]), .B2(n2579), 
        .ZN(n14096) );
  MOAI22 U23010 ( .A1(n29182), .A2(n2580), .B1(ram[9856]), .B2(n2581), 
        .ZN(n14097) );
  MOAI22 U23011 ( .A1(n28947), .A2(n2580), .B1(ram[9857]), .B2(n2581), 
        .ZN(n14098) );
  MOAI22 U23012 ( .A1(n28712), .A2(n2580), .B1(ram[9858]), .B2(n2581), 
        .ZN(n14099) );
  MOAI22 U23013 ( .A1(n28477), .A2(n2580), .B1(ram[9859]), .B2(n2581), 
        .ZN(n14100) );
  MOAI22 U23014 ( .A1(n28242), .A2(n2580), .B1(ram[9860]), .B2(n2581), 
        .ZN(n14101) );
  MOAI22 U23015 ( .A1(n28007), .A2(n2580), .B1(ram[9861]), .B2(n2581), 
        .ZN(n14102) );
  MOAI22 U23016 ( .A1(n27772), .A2(n2580), .B1(ram[9862]), .B2(n2581), 
        .ZN(n14103) );
  MOAI22 U23017 ( .A1(n27537), .A2(n2580), .B1(ram[9863]), .B2(n2581), 
        .ZN(n14104) );
  MOAI22 U23018 ( .A1(n29182), .A2(n2582), .B1(ram[9864]), .B2(n2583), 
        .ZN(n14105) );
  MOAI22 U23019 ( .A1(n28947), .A2(n2582), .B1(ram[9865]), .B2(n2583), 
        .ZN(n14106) );
  MOAI22 U23020 ( .A1(n28712), .A2(n2582), .B1(ram[9866]), .B2(n2583), 
        .ZN(n14107) );
  MOAI22 U23021 ( .A1(n28477), .A2(n2582), .B1(ram[9867]), .B2(n2583), 
        .ZN(n14108) );
  MOAI22 U23022 ( .A1(n28242), .A2(n2582), .B1(ram[9868]), .B2(n2583), 
        .ZN(n14109) );
  MOAI22 U23023 ( .A1(n28007), .A2(n2582), .B1(ram[9869]), .B2(n2583), 
        .ZN(n14110) );
  MOAI22 U23024 ( .A1(n27772), .A2(n2582), .B1(ram[9870]), .B2(n2583), 
        .ZN(n14111) );
  MOAI22 U23025 ( .A1(n27537), .A2(n2582), .B1(ram[9871]), .B2(n2583), 
        .ZN(n14112) );
  MOAI22 U23026 ( .A1(n29182), .A2(n2584), .B1(ram[9872]), .B2(n2585), 
        .ZN(n14113) );
  MOAI22 U23027 ( .A1(n28947), .A2(n2584), .B1(ram[9873]), .B2(n2585), 
        .ZN(n14114) );
  MOAI22 U23028 ( .A1(n28712), .A2(n2584), .B1(ram[9874]), .B2(n2585), 
        .ZN(n14115) );
  MOAI22 U23029 ( .A1(n28477), .A2(n2584), .B1(ram[9875]), .B2(n2585), 
        .ZN(n14116) );
  MOAI22 U23030 ( .A1(n28242), .A2(n2584), .B1(ram[9876]), .B2(n2585), 
        .ZN(n14117) );
  MOAI22 U23031 ( .A1(n28007), .A2(n2584), .B1(ram[9877]), .B2(n2585), 
        .ZN(n14118) );
  MOAI22 U23032 ( .A1(n27772), .A2(n2584), .B1(ram[9878]), .B2(n2585), 
        .ZN(n14119) );
  MOAI22 U23033 ( .A1(n27537), .A2(n2584), .B1(ram[9879]), .B2(n2585), 
        .ZN(n14120) );
  MOAI22 U23034 ( .A1(n29183), .A2(n2586), .B1(ram[9880]), .B2(n2587), 
        .ZN(n14121) );
  MOAI22 U23035 ( .A1(n28948), .A2(n2586), .B1(ram[9881]), .B2(n2587), 
        .ZN(n14122) );
  MOAI22 U23036 ( .A1(n28713), .A2(n2586), .B1(ram[9882]), .B2(n2587), 
        .ZN(n14123) );
  MOAI22 U23037 ( .A1(n28478), .A2(n2586), .B1(ram[9883]), .B2(n2587), 
        .ZN(n14124) );
  MOAI22 U23038 ( .A1(n28243), .A2(n2586), .B1(ram[9884]), .B2(n2587), 
        .ZN(n14125) );
  MOAI22 U23039 ( .A1(n28008), .A2(n2586), .B1(ram[9885]), .B2(n2587), 
        .ZN(n14126) );
  MOAI22 U23040 ( .A1(n27773), .A2(n2586), .B1(ram[9886]), .B2(n2587), 
        .ZN(n14127) );
  MOAI22 U23041 ( .A1(n27538), .A2(n2586), .B1(ram[9887]), .B2(n2587), 
        .ZN(n14128) );
  MOAI22 U23042 ( .A1(n29183), .A2(n2588), .B1(ram[9888]), .B2(n2589), 
        .ZN(n14129) );
  MOAI22 U23043 ( .A1(n28948), .A2(n2588), .B1(ram[9889]), .B2(n2589), 
        .ZN(n14130) );
  MOAI22 U23044 ( .A1(n28713), .A2(n2588), .B1(ram[9890]), .B2(n2589), 
        .ZN(n14131) );
  MOAI22 U23045 ( .A1(n28478), .A2(n2588), .B1(ram[9891]), .B2(n2589), 
        .ZN(n14132) );
  MOAI22 U23046 ( .A1(n28243), .A2(n2588), .B1(ram[9892]), .B2(n2589), 
        .ZN(n14133) );
  MOAI22 U23047 ( .A1(n28008), .A2(n2588), .B1(ram[9893]), .B2(n2589), 
        .ZN(n14134) );
  MOAI22 U23048 ( .A1(n27773), .A2(n2588), .B1(ram[9894]), .B2(n2589), 
        .ZN(n14135) );
  MOAI22 U23049 ( .A1(n27538), .A2(n2588), .B1(ram[9895]), .B2(n2589), 
        .ZN(n14136) );
  MOAI22 U23050 ( .A1(n29183), .A2(n2590), .B1(ram[9896]), .B2(n2591), 
        .ZN(n14137) );
  MOAI22 U23051 ( .A1(n28948), .A2(n2590), .B1(ram[9897]), .B2(n2591), 
        .ZN(n14138) );
  MOAI22 U23052 ( .A1(n28713), .A2(n2590), .B1(ram[9898]), .B2(n2591), 
        .ZN(n14139) );
  MOAI22 U23053 ( .A1(n28478), .A2(n2590), .B1(ram[9899]), .B2(n2591), 
        .ZN(n14140) );
  MOAI22 U23054 ( .A1(n28243), .A2(n2590), .B1(ram[9900]), .B2(n2591), 
        .ZN(n14141) );
  MOAI22 U23055 ( .A1(n28008), .A2(n2590), .B1(ram[9901]), .B2(n2591), 
        .ZN(n14142) );
  MOAI22 U23056 ( .A1(n27773), .A2(n2590), .B1(ram[9902]), .B2(n2591), 
        .ZN(n14143) );
  MOAI22 U23057 ( .A1(n27538), .A2(n2590), .B1(ram[9903]), .B2(n2591), 
        .ZN(n14144) );
  MOAI22 U23058 ( .A1(n29183), .A2(n2592), .B1(ram[9904]), .B2(n2593), 
        .ZN(n14145) );
  MOAI22 U23059 ( .A1(n28948), .A2(n2592), .B1(ram[9905]), .B2(n2593), 
        .ZN(n14146) );
  MOAI22 U23060 ( .A1(n28713), .A2(n2592), .B1(ram[9906]), .B2(n2593), 
        .ZN(n14147) );
  MOAI22 U23061 ( .A1(n28478), .A2(n2592), .B1(ram[9907]), .B2(n2593), 
        .ZN(n14148) );
  MOAI22 U23062 ( .A1(n28243), .A2(n2592), .B1(ram[9908]), .B2(n2593), 
        .ZN(n14149) );
  MOAI22 U23063 ( .A1(n28008), .A2(n2592), .B1(ram[9909]), .B2(n2593), 
        .ZN(n14150) );
  MOAI22 U23064 ( .A1(n27773), .A2(n2592), .B1(ram[9910]), .B2(n2593), 
        .ZN(n14151) );
  MOAI22 U23065 ( .A1(n27538), .A2(n2592), .B1(ram[9911]), .B2(n2593), 
        .ZN(n14152) );
  MOAI22 U23066 ( .A1(n29183), .A2(n2594), .B1(ram[9912]), .B2(n2595), 
        .ZN(n14153) );
  MOAI22 U23067 ( .A1(n28948), .A2(n2594), .B1(ram[9913]), .B2(n2595), 
        .ZN(n14154) );
  MOAI22 U23068 ( .A1(n28713), .A2(n2594), .B1(ram[9914]), .B2(n2595), 
        .ZN(n14155) );
  MOAI22 U23069 ( .A1(n28478), .A2(n2594), .B1(ram[9915]), .B2(n2595), 
        .ZN(n14156) );
  MOAI22 U23070 ( .A1(n28243), .A2(n2594), .B1(ram[9916]), .B2(n2595), 
        .ZN(n14157) );
  MOAI22 U23071 ( .A1(n28008), .A2(n2594), .B1(ram[9917]), .B2(n2595), 
        .ZN(n14158) );
  MOAI22 U23072 ( .A1(n27773), .A2(n2594), .B1(ram[9918]), .B2(n2595), 
        .ZN(n14159) );
  MOAI22 U23073 ( .A1(n27538), .A2(n2594), .B1(ram[9919]), .B2(n2595), 
        .ZN(n14160) );
  MOAI22 U23074 ( .A1(n29183), .A2(n2596), .B1(ram[9920]), .B2(n2597), 
        .ZN(n14161) );
  MOAI22 U23075 ( .A1(n28948), .A2(n2596), .B1(ram[9921]), .B2(n2597), 
        .ZN(n14162) );
  MOAI22 U23076 ( .A1(n28713), .A2(n2596), .B1(ram[9922]), .B2(n2597), 
        .ZN(n14163) );
  MOAI22 U23077 ( .A1(n28478), .A2(n2596), .B1(ram[9923]), .B2(n2597), 
        .ZN(n14164) );
  MOAI22 U23078 ( .A1(n28243), .A2(n2596), .B1(ram[9924]), .B2(n2597), 
        .ZN(n14165) );
  MOAI22 U23079 ( .A1(n28008), .A2(n2596), .B1(ram[9925]), .B2(n2597), 
        .ZN(n14166) );
  MOAI22 U23080 ( .A1(n27773), .A2(n2596), .B1(ram[9926]), .B2(n2597), 
        .ZN(n14167) );
  MOAI22 U23081 ( .A1(n27538), .A2(n2596), .B1(ram[9927]), .B2(n2597), 
        .ZN(n14168) );
  MOAI22 U23082 ( .A1(n29183), .A2(n2598), .B1(ram[9928]), .B2(n2599), 
        .ZN(n14169) );
  MOAI22 U23083 ( .A1(n28948), .A2(n2598), .B1(ram[9929]), .B2(n2599), 
        .ZN(n14170) );
  MOAI22 U23084 ( .A1(n28713), .A2(n2598), .B1(ram[9930]), .B2(n2599), 
        .ZN(n14171) );
  MOAI22 U23085 ( .A1(n28478), .A2(n2598), .B1(ram[9931]), .B2(n2599), 
        .ZN(n14172) );
  MOAI22 U23086 ( .A1(n28243), .A2(n2598), .B1(ram[9932]), .B2(n2599), 
        .ZN(n14173) );
  MOAI22 U23087 ( .A1(n28008), .A2(n2598), .B1(ram[9933]), .B2(n2599), 
        .ZN(n14174) );
  MOAI22 U23088 ( .A1(n27773), .A2(n2598), .B1(ram[9934]), .B2(n2599), 
        .ZN(n14175) );
  MOAI22 U23089 ( .A1(n27538), .A2(n2598), .B1(ram[9935]), .B2(n2599), 
        .ZN(n14176) );
  MOAI22 U23090 ( .A1(n29183), .A2(n2600), .B1(ram[9936]), .B2(n2601), 
        .ZN(n14177) );
  MOAI22 U23091 ( .A1(n28948), .A2(n2600), .B1(ram[9937]), .B2(n2601), 
        .ZN(n14178) );
  MOAI22 U23092 ( .A1(n28713), .A2(n2600), .B1(ram[9938]), .B2(n2601), 
        .ZN(n14179) );
  MOAI22 U23093 ( .A1(n28478), .A2(n2600), .B1(ram[9939]), .B2(n2601), 
        .ZN(n14180) );
  MOAI22 U23094 ( .A1(n28243), .A2(n2600), .B1(ram[9940]), .B2(n2601), 
        .ZN(n14181) );
  MOAI22 U23095 ( .A1(n28008), .A2(n2600), .B1(ram[9941]), .B2(n2601), 
        .ZN(n14182) );
  MOAI22 U23096 ( .A1(n27773), .A2(n2600), .B1(ram[9942]), .B2(n2601), 
        .ZN(n14183) );
  MOAI22 U23097 ( .A1(n27538), .A2(n2600), .B1(ram[9943]), .B2(n2601), 
        .ZN(n14184) );
  MOAI22 U23098 ( .A1(n29183), .A2(n2602), .B1(ram[9944]), .B2(n2603), 
        .ZN(n14185) );
  MOAI22 U23099 ( .A1(n28948), .A2(n2602), .B1(ram[9945]), .B2(n2603), 
        .ZN(n14186) );
  MOAI22 U23100 ( .A1(n28713), .A2(n2602), .B1(ram[9946]), .B2(n2603), 
        .ZN(n14187) );
  MOAI22 U23101 ( .A1(n28478), .A2(n2602), .B1(ram[9947]), .B2(n2603), 
        .ZN(n14188) );
  MOAI22 U23102 ( .A1(n28243), .A2(n2602), .B1(ram[9948]), .B2(n2603), 
        .ZN(n14189) );
  MOAI22 U23103 ( .A1(n28008), .A2(n2602), .B1(ram[9949]), .B2(n2603), 
        .ZN(n14190) );
  MOAI22 U23104 ( .A1(n27773), .A2(n2602), .B1(ram[9950]), .B2(n2603), 
        .ZN(n14191) );
  MOAI22 U23105 ( .A1(n27538), .A2(n2602), .B1(ram[9951]), .B2(n2603), 
        .ZN(n14192) );
  MOAI22 U23106 ( .A1(n29183), .A2(n2604), .B1(ram[9952]), .B2(n2605), 
        .ZN(n14193) );
  MOAI22 U23107 ( .A1(n28948), .A2(n2604), .B1(ram[9953]), .B2(n2605), 
        .ZN(n14194) );
  MOAI22 U23108 ( .A1(n28713), .A2(n2604), .B1(ram[9954]), .B2(n2605), 
        .ZN(n14195) );
  MOAI22 U23109 ( .A1(n28478), .A2(n2604), .B1(ram[9955]), .B2(n2605), 
        .ZN(n14196) );
  MOAI22 U23110 ( .A1(n28243), .A2(n2604), .B1(ram[9956]), .B2(n2605), 
        .ZN(n14197) );
  MOAI22 U23111 ( .A1(n28008), .A2(n2604), .B1(ram[9957]), .B2(n2605), 
        .ZN(n14198) );
  MOAI22 U23112 ( .A1(n27773), .A2(n2604), .B1(ram[9958]), .B2(n2605), 
        .ZN(n14199) );
  MOAI22 U23113 ( .A1(n27538), .A2(n2604), .B1(ram[9959]), .B2(n2605), 
        .ZN(n14200) );
  MOAI22 U23114 ( .A1(n29183), .A2(n2606), .B1(ram[9960]), .B2(n2607), 
        .ZN(n14201) );
  MOAI22 U23115 ( .A1(n28948), .A2(n2606), .B1(ram[9961]), .B2(n2607), 
        .ZN(n14202) );
  MOAI22 U23116 ( .A1(n28713), .A2(n2606), .B1(ram[9962]), .B2(n2607), 
        .ZN(n14203) );
  MOAI22 U23117 ( .A1(n28478), .A2(n2606), .B1(ram[9963]), .B2(n2607), 
        .ZN(n14204) );
  MOAI22 U23118 ( .A1(n28243), .A2(n2606), .B1(ram[9964]), .B2(n2607), 
        .ZN(n14205) );
  MOAI22 U23119 ( .A1(n28008), .A2(n2606), .B1(ram[9965]), .B2(n2607), 
        .ZN(n14206) );
  MOAI22 U23120 ( .A1(n27773), .A2(n2606), .B1(ram[9966]), .B2(n2607), 
        .ZN(n14207) );
  MOAI22 U23121 ( .A1(n27538), .A2(n2606), .B1(ram[9967]), .B2(n2607), 
        .ZN(n14208) );
  MOAI22 U23122 ( .A1(n29183), .A2(n2608), .B1(ram[9968]), .B2(n2609), 
        .ZN(n14209) );
  MOAI22 U23123 ( .A1(n28948), .A2(n2608), .B1(ram[9969]), .B2(n2609), 
        .ZN(n14210) );
  MOAI22 U23124 ( .A1(n28713), .A2(n2608), .B1(ram[9970]), .B2(n2609), 
        .ZN(n14211) );
  MOAI22 U23125 ( .A1(n28478), .A2(n2608), .B1(ram[9971]), .B2(n2609), 
        .ZN(n14212) );
  MOAI22 U23126 ( .A1(n28243), .A2(n2608), .B1(ram[9972]), .B2(n2609), 
        .ZN(n14213) );
  MOAI22 U23127 ( .A1(n28008), .A2(n2608), .B1(ram[9973]), .B2(n2609), 
        .ZN(n14214) );
  MOAI22 U23128 ( .A1(n27773), .A2(n2608), .B1(ram[9974]), .B2(n2609), 
        .ZN(n14215) );
  MOAI22 U23129 ( .A1(n27538), .A2(n2608), .B1(ram[9975]), .B2(n2609), 
        .ZN(n14216) );
  MOAI22 U23130 ( .A1(n29183), .A2(n2610), .B1(ram[9976]), .B2(n2611), 
        .ZN(n14217) );
  MOAI22 U23131 ( .A1(n28948), .A2(n2610), .B1(ram[9977]), .B2(n2611), 
        .ZN(n14218) );
  MOAI22 U23132 ( .A1(n28713), .A2(n2610), .B1(ram[9978]), .B2(n2611), 
        .ZN(n14219) );
  MOAI22 U23133 ( .A1(n28478), .A2(n2610), .B1(ram[9979]), .B2(n2611), 
        .ZN(n14220) );
  MOAI22 U23134 ( .A1(n28243), .A2(n2610), .B1(ram[9980]), .B2(n2611), 
        .ZN(n14221) );
  MOAI22 U23135 ( .A1(n28008), .A2(n2610), .B1(ram[9981]), .B2(n2611), 
        .ZN(n14222) );
  MOAI22 U23136 ( .A1(n27773), .A2(n2610), .B1(ram[9982]), .B2(n2611), 
        .ZN(n14223) );
  MOAI22 U23137 ( .A1(n27538), .A2(n2610), .B1(ram[9983]), .B2(n2611), 
        .ZN(n14224) );
  MOAI22 U23138 ( .A1(n29184), .A2(n2612), .B1(ram[9984]), .B2(n2613), 
        .ZN(n14225) );
  MOAI22 U23139 ( .A1(n28949), .A2(n2612), .B1(ram[9985]), .B2(n2613), 
        .ZN(n14226) );
  MOAI22 U23140 ( .A1(n28714), .A2(n2612), .B1(ram[9986]), .B2(n2613), 
        .ZN(n14227) );
  MOAI22 U23141 ( .A1(n28479), .A2(n2612), .B1(ram[9987]), .B2(n2613), 
        .ZN(n14228) );
  MOAI22 U23142 ( .A1(n28244), .A2(n2612), .B1(ram[9988]), .B2(n2613), 
        .ZN(n14229) );
  MOAI22 U23143 ( .A1(n28009), .A2(n2612), .B1(ram[9989]), .B2(n2613), 
        .ZN(n14230) );
  MOAI22 U23144 ( .A1(n27774), .A2(n2612), .B1(ram[9990]), .B2(n2613), 
        .ZN(n14231) );
  MOAI22 U23145 ( .A1(n27539), .A2(n2612), .B1(ram[9991]), .B2(n2613), 
        .ZN(n14232) );
  MOAI22 U23146 ( .A1(n29184), .A2(n2614), .B1(ram[9992]), .B2(n2615), 
        .ZN(n14233) );
  MOAI22 U23147 ( .A1(n28949), .A2(n2614), .B1(ram[9993]), .B2(n2615), 
        .ZN(n14234) );
  MOAI22 U23148 ( .A1(n28714), .A2(n2614), .B1(ram[9994]), .B2(n2615), 
        .ZN(n14235) );
  MOAI22 U23149 ( .A1(n28479), .A2(n2614), .B1(ram[9995]), .B2(n2615), 
        .ZN(n14236) );
  MOAI22 U23150 ( .A1(n28244), .A2(n2614), .B1(ram[9996]), .B2(n2615), 
        .ZN(n14237) );
  MOAI22 U23151 ( .A1(n28009), .A2(n2614), .B1(ram[9997]), .B2(n2615), 
        .ZN(n14238) );
  MOAI22 U23152 ( .A1(n27774), .A2(n2614), .B1(ram[9998]), .B2(n2615), 
        .ZN(n14239) );
  MOAI22 U23153 ( .A1(n27539), .A2(n2614), .B1(ram[9999]), .B2(n2615), 
        .ZN(n14240) );
  MOAI22 U23154 ( .A1(n29184), .A2(n2616), .B1(ram[10000]), .B2(n2617), 
        .ZN(n14241) );
  MOAI22 U23155 ( .A1(n28949), .A2(n2616), .B1(ram[10001]), .B2(n2617), 
        .ZN(n14242) );
  MOAI22 U23156 ( .A1(n28714), .A2(n2616), .B1(ram[10002]), .B2(n2617), 
        .ZN(n14243) );
  MOAI22 U23157 ( .A1(n28479), .A2(n2616), .B1(ram[10003]), .B2(n2617), 
        .ZN(n14244) );
  MOAI22 U23158 ( .A1(n28244), .A2(n2616), .B1(ram[10004]), .B2(n2617), 
        .ZN(n14245) );
  MOAI22 U23159 ( .A1(n28009), .A2(n2616), .B1(ram[10005]), .B2(n2617), 
        .ZN(n14246) );
  MOAI22 U23160 ( .A1(n27774), .A2(n2616), .B1(ram[10006]), .B2(n2617), 
        .ZN(n14247) );
  MOAI22 U23161 ( .A1(n27539), .A2(n2616), .B1(ram[10007]), .B2(n2617), 
        .ZN(n14248) );
  MOAI22 U23162 ( .A1(n29184), .A2(n2618), .B1(ram[10008]), .B2(n2619), 
        .ZN(n14249) );
  MOAI22 U23163 ( .A1(n28949), .A2(n2618), .B1(ram[10009]), .B2(n2619), 
        .ZN(n14250) );
  MOAI22 U23164 ( .A1(n28714), .A2(n2618), .B1(ram[10010]), .B2(n2619), 
        .ZN(n14251) );
  MOAI22 U23165 ( .A1(n28479), .A2(n2618), .B1(ram[10011]), .B2(n2619), 
        .ZN(n14252) );
  MOAI22 U23166 ( .A1(n28244), .A2(n2618), .B1(ram[10012]), .B2(n2619), 
        .ZN(n14253) );
  MOAI22 U23167 ( .A1(n28009), .A2(n2618), .B1(ram[10013]), .B2(n2619), 
        .ZN(n14254) );
  MOAI22 U23168 ( .A1(n27774), .A2(n2618), .B1(ram[10014]), .B2(n2619), 
        .ZN(n14255) );
  MOAI22 U23169 ( .A1(n27539), .A2(n2618), .B1(ram[10015]), .B2(n2619), 
        .ZN(n14256) );
  MOAI22 U23170 ( .A1(n29184), .A2(n2620), .B1(ram[10016]), .B2(n2621), 
        .ZN(n14257) );
  MOAI22 U23171 ( .A1(n28949), .A2(n2620), .B1(ram[10017]), .B2(n2621), 
        .ZN(n14258) );
  MOAI22 U23172 ( .A1(n28714), .A2(n2620), .B1(ram[10018]), .B2(n2621), 
        .ZN(n14259) );
  MOAI22 U23173 ( .A1(n28479), .A2(n2620), .B1(ram[10019]), .B2(n2621), 
        .ZN(n14260) );
  MOAI22 U23174 ( .A1(n28244), .A2(n2620), .B1(ram[10020]), .B2(n2621), 
        .ZN(n14261) );
  MOAI22 U23175 ( .A1(n28009), .A2(n2620), .B1(ram[10021]), .B2(n2621), 
        .ZN(n14262) );
  MOAI22 U23176 ( .A1(n27774), .A2(n2620), .B1(ram[10022]), .B2(n2621), 
        .ZN(n14263) );
  MOAI22 U23177 ( .A1(n27539), .A2(n2620), .B1(ram[10023]), .B2(n2621), 
        .ZN(n14264) );
  MOAI22 U23178 ( .A1(n29184), .A2(n2622), .B1(ram[10024]), .B2(n2623), 
        .ZN(n14265) );
  MOAI22 U23179 ( .A1(n28949), .A2(n2622), .B1(ram[10025]), .B2(n2623), 
        .ZN(n14266) );
  MOAI22 U23180 ( .A1(n28714), .A2(n2622), .B1(ram[10026]), .B2(n2623), 
        .ZN(n14267) );
  MOAI22 U23181 ( .A1(n28479), .A2(n2622), .B1(ram[10027]), .B2(n2623), 
        .ZN(n14268) );
  MOAI22 U23182 ( .A1(n28244), .A2(n2622), .B1(ram[10028]), .B2(n2623), 
        .ZN(n14269) );
  MOAI22 U23183 ( .A1(n28009), .A2(n2622), .B1(ram[10029]), .B2(n2623), 
        .ZN(n14270) );
  MOAI22 U23184 ( .A1(n27774), .A2(n2622), .B1(ram[10030]), .B2(n2623), 
        .ZN(n14271) );
  MOAI22 U23185 ( .A1(n27539), .A2(n2622), .B1(ram[10031]), .B2(n2623), 
        .ZN(n14272) );
  MOAI22 U23186 ( .A1(n29184), .A2(n2624), .B1(ram[10032]), .B2(n2625), 
        .ZN(n14273) );
  MOAI22 U23187 ( .A1(n28949), .A2(n2624), .B1(ram[10033]), .B2(n2625), 
        .ZN(n14274) );
  MOAI22 U23188 ( .A1(n28714), .A2(n2624), .B1(ram[10034]), .B2(n2625), 
        .ZN(n14275) );
  MOAI22 U23189 ( .A1(n28479), .A2(n2624), .B1(ram[10035]), .B2(n2625), 
        .ZN(n14276) );
  MOAI22 U23190 ( .A1(n28244), .A2(n2624), .B1(ram[10036]), .B2(n2625), 
        .ZN(n14277) );
  MOAI22 U23191 ( .A1(n28009), .A2(n2624), .B1(ram[10037]), .B2(n2625), 
        .ZN(n14278) );
  MOAI22 U23192 ( .A1(n27774), .A2(n2624), .B1(ram[10038]), .B2(n2625), 
        .ZN(n14279) );
  MOAI22 U23193 ( .A1(n27539), .A2(n2624), .B1(ram[10039]), .B2(n2625), 
        .ZN(n14280) );
  MOAI22 U23194 ( .A1(n29184), .A2(n2626), .B1(ram[10040]), .B2(n2627), 
        .ZN(n14281) );
  MOAI22 U23195 ( .A1(n28949), .A2(n2626), .B1(ram[10041]), .B2(n2627), 
        .ZN(n14282) );
  MOAI22 U23196 ( .A1(n28714), .A2(n2626), .B1(ram[10042]), .B2(n2627), 
        .ZN(n14283) );
  MOAI22 U23197 ( .A1(n28479), .A2(n2626), .B1(ram[10043]), .B2(n2627), 
        .ZN(n14284) );
  MOAI22 U23198 ( .A1(n28244), .A2(n2626), .B1(ram[10044]), .B2(n2627), 
        .ZN(n14285) );
  MOAI22 U23199 ( .A1(n28009), .A2(n2626), .B1(ram[10045]), .B2(n2627), 
        .ZN(n14286) );
  MOAI22 U23200 ( .A1(n27774), .A2(n2626), .B1(ram[10046]), .B2(n2627), 
        .ZN(n14287) );
  MOAI22 U23201 ( .A1(n27539), .A2(n2626), .B1(ram[10047]), .B2(n2627), 
        .ZN(n14288) );
  MOAI22 U23202 ( .A1(n29184), .A2(n2628), .B1(ram[10048]), .B2(n2629), 
        .ZN(n14289) );
  MOAI22 U23203 ( .A1(n28949), .A2(n2628), .B1(ram[10049]), .B2(n2629), 
        .ZN(n14290) );
  MOAI22 U23204 ( .A1(n28714), .A2(n2628), .B1(ram[10050]), .B2(n2629), 
        .ZN(n14291) );
  MOAI22 U23205 ( .A1(n28479), .A2(n2628), .B1(ram[10051]), .B2(n2629), 
        .ZN(n14292) );
  MOAI22 U23206 ( .A1(n28244), .A2(n2628), .B1(ram[10052]), .B2(n2629), 
        .ZN(n14293) );
  MOAI22 U23207 ( .A1(n28009), .A2(n2628), .B1(ram[10053]), .B2(n2629), 
        .ZN(n14294) );
  MOAI22 U23208 ( .A1(n27774), .A2(n2628), .B1(ram[10054]), .B2(n2629), 
        .ZN(n14295) );
  MOAI22 U23209 ( .A1(n27539), .A2(n2628), .B1(ram[10055]), .B2(n2629), 
        .ZN(n14296) );
  MOAI22 U23210 ( .A1(n29184), .A2(n2630), .B1(ram[10056]), .B2(n2631), 
        .ZN(n14297) );
  MOAI22 U23211 ( .A1(n28949), .A2(n2630), .B1(ram[10057]), .B2(n2631), 
        .ZN(n14298) );
  MOAI22 U23212 ( .A1(n28714), .A2(n2630), .B1(ram[10058]), .B2(n2631), 
        .ZN(n14299) );
  MOAI22 U23213 ( .A1(n28479), .A2(n2630), .B1(ram[10059]), .B2(n2631), 
        .ZN(n14300) );
  MOAI22 U23214 ( .A1(n28244), .A2(n2630), .B1(ram[10060]), .B2(n2631), 
        .ZN(n14301) );
  MOAI22 U23215 ( .A1(n28009), .A2(n2630), .B1(ram[10061]), .B2(n2631), 
        .ZN(n14302) );
  MOAI22 U23216 ( .A1(n27774), .A2(n2630), .B1(ram[10062]), .B2(n2631), 
        .ZN(n14303) );
  MOAI22 U23217 ( .A1(n27539), .A2(n2630), .B1(ram[10063]), .B2(n2631), 
        .ZN(n14304) );
  MOAI22 U23218 ( .A1(n29184), .A2(n2632), .B1(ram[10064]), .B2(n2633), 
        .ZN(n14305) );
  MOAI22 U23219 ( .A1(n28949), .A2(n2632), .B1(ram[10065]), .B2(n2633), 
        .ZN(n14306) );
  MOAI22 U23220 ( .A1(n28714), .A2(n2632), .B1(ram[10066]), .B2(n2633), 
        .ZN(n14307) );
  MOAI22 U23221 ( .A1(n28479), .A2(n2632), .B1(ram[10067]), .B2(n2633), 
        .ZN(n14308) );
  MOAI22 U23222 ( .A1(n28244), .A2(n2632), .B1(ram[10068]), .B2(n2633), 
        .ZN(n14309) );
  MOAI22 U23223 ( .A1(n28009), .A2(n2632), .B1(ram[10069]), .B2(n2633), 
        .ZN(n14310) );
  MOAI22 U23224 ( .A1(n27774), .A2(n2632), .B1(ram[10070]), .B2(n2633), 
        .ZN(n14311) );
  MOAI22 U23225 ( .A1(n27539), .A2(n2632), .B1(ram[10071]), .B2(n2633), 
        .ZN(n14312) );
  MOAI22 U23226 ( .A1(n29184), .A2(n2634), .B1(ram[10072]), .B2(n2635), 
        .ZN(n14313) );
  MOAI22 U23227 ( .A1(n28949), .A2(n2634), .B1(ram[10073]), .B2(n2635), 
        .ZN(n14314) );
  MOAI22 U23228 ( .A1(n28714), .A2(n2634), .B1(ram[10074]), .B2(n2635), 
        .ZN(n14315) );
  MOAI22 U23229 ( .A1(n28479), .A2(n2634), .B1(ram[10075]), .B2(n2635), 
        .ZN(n14316) );
  MOAI22 U23230 ( .A1(n28244), .A2(n2634), .B1(ram[10076]), .B2(n2635), 
        .ZN(n14317) );
  MOAI22 U23231 ( .A1(n28009), .A2(n2634), .B1(ram[10077]), .B2(n2635), 
        .ZN(n14318) );
  MOAI22 U23232 ( .A1(n27774), .A2(n2634), .B1(ram[10078]), .B2(n2635), 
        .ZN(n14319) );
  MOAI22 U23233 ( .A1(n27539), .A2(n2634), .B1(ram[10079]), .B2(n2635), 
        .ZN(n14320) );
  MOAI22 U23234 ( .A1(n29184), .A2(n2636), .B1(ram[10080]), .B2(n2637), 
        .ZN(n14321) );
  MOAI22 U23235 ( .A1(n28949), .A2(n2636), .B1(ram[10081]), .B2(n2637), 
        .ZN(n14322) );
  MOAI22 U23236 ( .A1(n28714), .A2(n2636), .B1(ram[10082]), .B2(n2637), 
        .ZN(n14323) );
  MOAI22 U23237 ( .A1(n28479), .A2(n2636), .B1(ram[10083]), .B2(n2637), 
        .ZN(n14324) );
  MOAI22 U23238 ( .A1(n28244), .A2(n2636), .B1(ram[10084]), .B2(n2637), 
        .ZN(n14325) );
  MOAI22 U23239 ( .A1(n28009), .A2(n2636), .B1(ram[10085]), .B2(n2637), 
        .ZN(n14326) );
  MOAI22 U23240 ( .A1(n27774), .A2(n2636), .B1(ram[10086]), .B2(n2637), 
        .ZN(n14327) );
  MOAI22 U23241 ( .A1(n27539), .A2(n2636), .B1(ram[10087]), .B2(n2637), 
        .ZN(n14328) );
  MOAI22 U23242 ( .A1(n29185), .A2(n2638), .B1(ram[10088]), .B2(n2639), 
        .ZN(n14329) );
  MOAI22 U23243 ( .A1(n28950), .A2(n2638), .B1(ram[10089]), .B2(n2639), 
        .ZN(n14330) );
  MOAI22 U23244 ( .A1(n28715), .A2(n2638), .B1(ram[10090]), .B2(n2639), 
        .ZN(n14331) );
  MOAI22 U23245 ( .A1(n28480), .A2(n2638), .B1(ram[10091]), .B2(n2639), 
        .ZN(n14332) );
  MOAI22 U23246 ( .A1(n28245), .A2(n2638), .B1(ram[10092]), .B2(n2639), 
        .ZN(n14333) );
  MOAI22 U23247 ( .A1(n28010), .A2(n2638), .B1(ram[10093]), .B2(n2639), 
        .ZN(n14334) );
  MOAI22 U23248 ( .A1(n27775), .A2(n2638), .B1(ram[10094]), .B2(n2639), 
        .ZN(n14335) );
  MOAI22 U23249 ( .A1(n27540), .A2(n2638), .B1(ram[10095]), .B2(n2639), 
        .ZN(n14336) );
  MOAI22 U23250 ( .A1(n29185), .A2(n2640), .B1(ram[10096]), .B2(n2641), 
        .ZN(n14337) );
  MOAI22 U23251 ( .A1(n28950), .A2(n2640), .B1(ram[10097]), .B2(n2641), 
        .ZN(n14338) );
  MOAI22 U23252 ( .A1(n28715), .A2(n2640), .B1(ram[10098]), .B2(n2641), 
        .ZN(n14339) );
  MOAI22 U23253 ( .A1(n28480), .A2(n2640), .B1(ram[10099]), .B2(n2641), 
        .ZN(n14340) );
  MOAI22 U23254 ( .A1(n28245), .A2(n2640), .B1(ram[10100]), .B2(n2641), 
        .ZN(n14341) );
  MOAI22 U23255 ( .A1(n28010), .A2(n2640), .B1(ram[10101]), .B2(n2641), 
        .ZN(n14342) );
  MOAI22 U23256 ( .A1(n27775), .A2(n2640), .B1(ram[10102]), .B2(n2641), 
        .ZN(n14343) );
  MOAI22 U23257 ( .A1(n27540), .A2(n2640), .B1(ram[10103]), .B2(n2641), 
        .ZN(n14344) );
  MOAI22 U23258 ( .A1(n29185), .A2(n2642), .B1(ram[10104]), .B2(n2643), 
        .ZN(n14345) );
  MOAI22 U23259 ( .A1(n28950), .A2(n2642), .B1(ram[10105]), .B2(n2643), 
        .ZN(n14346) );
  MOAI22 U23260 ( .A1(n28715), .A2(n2642), .B1(ram[10106]), .B2(n2643), 
        .ZN(n14347) );
  MOAI22 U23261 ( .A1(n28480), .A2(n2642), .B1(ram[10107]), .B2(n2643), 
        .ZN(n14348) );
  MOAI22 U23262 ( .A1(n28245), .A2(n2642), .B1(ram[10108]), .B2(n2643), 
        .ZN(n14349) );
  MOAI22 U23263 ( .A1(n28010), .A2(n2642), .B1(ram[10109]), .B2(n2643), 
        .ZN(n14350) );
  MOAI22 U23264 ( .A1(n27775), .A2(n2642), .B1(ram[10110]), .B2(n2643), 
        .ZN(n14351) );
  MOAI22 U23265 ( .A1(n27540), .A2(n2642), .B1(ram[10111]), .B2(n2643), 
        .ZN(n14352) );
  MOAI22 U23266 ( .A1(n29185), .A2(n2644), .B1(ram[10112]), .B2(n2645), 
        .ZN(n14353) );
  MOAI22 U23267 ( .A1(n28950), .A2(n2644), .B1(ram[10113]), .B2(n2645), 
        .ZN(n14354) );
  MOAI22 U23268 ( .A1(n28715), .A2(n2644), .B1(ram[10114]), .B2(n2645), 
        .ZN(n14355) );
  MOAI22 U23269 ( .A1(n28480), .A2(n2644), .B1(ram[10115]), .B2(n2645), 
        .ZN(n14356) );
  MOAI22 U23270 ( .A1(n28245), .A2(n2644), .B1(ram[10116]), .B2(n2645), 
        .ZN(n14357) );
  MOAI22 U23271 ( .A1(n28010), .A2(n2644), .B1(ram[10117]), .B2(n2645), 
        .ZN(n14358) );
  MOAI22 U23272 ( .A1(n27775), .A2(n2644), .B1(ram[10118]), .B2(n2645), 
        .ZN(n14359) );
  MOAI22 U23273 ( .A1(n27540), .A2(n2644), .B1(ram[10119]), .B2(n2645), 
        .ZN(n14360) );
  MOAI22 U23274 ( .A1(n29185), .A2(n2646), .B1(ram[10120]), .B2(n2647), 
        .ZN(n14361) );
  MOAI22 U23275 ( .A1(n28950), .A2(n2646), .B1(ram[10121]), .B2(n2647), 
        .ZN(n14362) );
  MOAI22 U23276 ( .A1(n28715), .A2(n2646), .B1(ram[10122]), .B2(n2647), 
        .ZN(n14363) );
  MOAI22 U23277 ( .A1(n28480), .A2(n2646), .B1(ram[10123]), .B2(n2647), 
        .ZN(n14364) );
  MOAI22 U23278 ( .A1(n28245), .A2(n2646), .B1(ram[10124]), .B2(n2647), 
        .ZN(n14365) );
  MOAI22 U23279 ( .A1(n28010), .A2(n2646), .B1(ram[10125]), .B2(n2647), 
        .ZN(n14366) );
  MOAI22 U23280 ( .A1(n27775), .A2(n2646), .B1(ram[10126]), .B2(n2647), 
        .ZN(n14367) );
  MOAI22 U23281 ( .A1(n27540), .A2(n2646), .B1(ram[10127]), .B2(n2647), 
        .ZN(n14368) );
  MOAI22 U23282 ( .A1(n29185), .A2(n2648), .B1(ram[10128]), .B2(n2649), 
        .ZN(n14369) );
  MOAI22 U23283 ( .A1(n28950), .A2(n2648), .B1(ram[10129]), .B2(n2649), 
        .ZN(n14370) );
  MOAI22 U23284 ( .A1(n28715), .A2(n2648), .B1(ram[10130]), .B2(n2649), 
        .ZN(n14371) );
  MOAI22 U23285 ( .A1(n28480), .A2(n2648), .B1(ram[10131]), .B2(n2649), 
        .ZN(n14372) );
  MOAI22 U23286 ( .A1(n28245), .A2(n2648), .B1(ram[10132]), .B2(n2649), 
        .ZN(n14373) );
  MOAI22 U23287 ( .A1(n28010), .A2(n2648), .B1(ram[10133]), .B2(n2649), 
        .ZN(n14374) );
  MOAI22 U23288 ( .A1(n27775), .A2(n2648), .B1(ram[10134]), .B2(n2649), 
        .ZN(n14375) );
  MOAI22 U23289 ( .A1(n27540), .A2(n2648), .B1(ram[10135]), .B2(n2649), 
        .ZN(n14376) );
  MOAI22 U23290 ( .A1(n29185), .A2(n2650), .B1(ram[10136]), .B2(n2651), 
        .ZN(n14377) );
  MOAI22 U23291 ( .A1(n28950), .A2(n2650), .B1(ram[10137]), .B2(n2651), 
        .ZN(n14378) );
  MOAI22 U23292 ( .A1(n28715), .A2(n2650), .B1(ram[10138]), .B2(n2651), 
        .ZN(n14379) );
  MOAI22 U23293 ( .A1(n28480), .A2(n2650), .B1(ram[10139]), .B2(n2651), 
        .ZN(n14380) );
  MOAI22 U23294 ( .A1(n28245), .A2(n2650), .B1(ram[10140]), .B2(n2651), 
        .ZN(n14381) );
  MOAI22 U23295 ( .A1(n28010), .A2(n2650), .B1(ram[10141]), .B2(n2651), 
        .ZN(n14382) );
  MOAI22 U23296 ( .A1(n27775), .A2(n2650), .B1(ram[10142]), .B2(n2651), 
        .ZN(n14383) );
  MOAI22 U23297 ( .A1(n27540), .A2(n2650), .B1(ram[10143]), .B2(n2651), 
        .ZN(n14384) );
  MOAI22 U23298 ( .A1(n29185), .A2(n2652), .B1(ram[10144]), .B2(n2653), 
        .ZN(n14385) );
  MOAI22 U23299 ( .A1(n28950), .A2(n2652), .B1(ram[10145]), .B2(n2653), 
        .ZN(n14386) );
  MOAI22 U23300 ( .A1(n28715), .A2(n2652), .B1(ram[10146]), .B2(n2653), 
        .ZN(n14387) );
  MOAI22 U23301 ( .A1(n28480), .A2(n2652), .B1(ram[10147]), .B2(n2653), 
        .ZN(n14388) );
  MOAI22 U23302 ( .A1(n28245), .A2(n2652), .B1(ram[10148]), .B2(n2653), 
        .ZN(n14389) );
  MOAI22 U23303 ( .A1(n28010), .A2(n2652), .B1(ram[10149]), .B2(n2653), 
        .ZN(n14390) );
  MOAI22 U23304 ( .A1(n27775), .A2(n2652), .B1(ram[10150]), .B2(n2653), 
        .ZN(n14391) );
  MOAI22 U23305 ( .A1(n27540), .A2(n2652), .B1(ram[10151]), .B2(n2653), 
        .ZN(n14392) );
  MOAI22 U23306 ( .A1(n29185), .A2(n2654), .B1(ram[10152]), .B2(n2655), 
        .ZN(n14393) );
  MOAI22 U23307 ( .A1(n28950), .A2(n2654), .B1(ram[10153]), .B2(n2655), 
        .ZN(n14394) );
  MOAI22 U23308 ( .A1(n28715), .A2(n2654), .B1(ram[10154]), .B2(n2655), 
        .ZN(n14395) );
  MOAI22 U23309 ( .A1(n28480), .A2(n2654), .B1(ram[10155]), .B2(n2655), 
        .ZN(n14396) );
  MOAI22 U23310 ( .A1(n28245), .A2(n2654), .B1(ram[10156]), .B2(n2655), 
        .ZN(n14397) );
  MOAI22 U23311 ( .A1(n28010), .A2(n2654), .B1(ram[10157]), .B2(n2655), 
        .ZN(n14398) );
  MOAI22 U23312 ( .A1(n27775), .A2(n2654), .B1(ram[10158]), .B2(n2655), 
        .ZN(n14399) );
  MOAI22 U23313 ( .A1(n27540), .A2(n2654), .B1(ram[10159]), .B2(n2655), 
        .ZN(n14400) );
  MOAI22 U23314 ( .A1(n29185), .A2(n2656), .B1(ram[10160]), .B2(n2657), 
        .ZN(n14401) );
  MOAI22 U23315 ( .A1(n28950), .A2(n2656), .B1(ram[10161]), .B2(n2657), 
        .ZN(n14402) );
  MOAI22 U23316 ( .A1(n28715), .A2(n2656), .B1(ram[10162]), .B2(n2657), 
        .ZN(n14403) );
  MOAI22 U23317 ( .A1(n28480), .A2(n2656), .B1(ram[10163]), .B2(n2657), 
        .ZN(n14404) );
  MOAI22 U23318 ( .A1(n28245), .A2(n2656), .B1(ram[10164]), .B2(n2657), 
        .ZN(n14405) );
  MOAI22 U23319 ( .A1(n28010), .A2(n2656), .B1(ram[10165]), .B2(n2657), 
        .ZN(n14406) );
  MOAI22 U23320 ( .A1(n27775), .A2(n2656), .B1(ram[10166]), .B2(n2657), 
        .ZN(n14407) );
  MOAI22 U23321 ( .A1(n27540), .A2(n2656), .B1(ram[10167]), .B2(n2657), 
        .ZN(n14408) );
  MOAI22 U23322 ( .A1(n29185), .A2(n2658), .B1(ram[10168]), .B2(n2659), 
        .ZN(n14409) );
  MOAI22 U23323 ( .A1(n28950), .A2(n2658), .B1(ram[10169]), .B2(n2659), 
        .ZN(n14410) );
  MOAI22 U23324 ( .A1(n28715), .A2(n2658), .B1(ram[10170]), .B2(n2659), 
        .ZN(n14411) );
  MOAI22 U23325 ( .A1(n28480), .A2(n2658), .B1(ram[10171]), .B2(n2659), 
        .ZN(n14412) );
  MOAI22 U23326 ( .A1(n28245), .A2(n2658), .B1(ram[10172]), .B2(n2659), 
        .ZN(n14413) );
  MOAI22 U23327 ( .A1(n28010), .A2(n2658), .B1(ram[10173]), .B2(n2659), 
        .ZN(n14414) );
  MOAI22 U23328 ( .A1(n27775), .A2(n2658), .B1(ram[10174]), .B2(n2659), 
        .ZN(n14415) );
  MOAI22 U23329 ( .A1(n27540), .A2(n2658), .B1(ram[10175]), .B2(n2659), 
        .ZN(n14416) );
  MOAI22 U23330 ( .A1(n29185), .A2(n2660), .B1(ram[10176]), .B2(n2661), 
        .ZN(n14417) );
  MOAI22 U23331 ( .A1(n28950), .A2(n2660), .B1(ram[10177]), .B2(n2661), 
        .ZN(n14418) );
  MOAI22 U23332 ( .A1(n28715), .A2(n2660), .B1(ram[10178]), .B2(n2661), 
        .ZN(n14419) );
  MOAI22 U23333 ( .A1(n28480), .A2(n2660), .B1(ram[10179]), .B2(n2661), 
        .ZN(n14420) );
  MOAI22 U23334 ( .A1(n28245), .A2(n2660), .B1(ram[10180]), .B2(n2661), 
        .ZN(n14421) );
  MOAI22 U23335 ( .A1(n28010), .A2(n2660), .B1(ram[10181]), .B2(n2661), 
        .ZN(n14422) );
  MOAI22 U23336 ( .A1(n27775), .A2(n2660), .B1(ram[10182]), .B2(n2661), 
        .ZN(n14423) );
  MOAI22 U23337 ( .A1(n27540), .A2(n2660), .B1(ram[10183]), .B2(n2661), 
        .ZN(n14424) );
  MOAI22 U23338 ( .A1(n29185), .A2(n2662), .B1(ram[10184]), .B2(n2663), 
        .ZN(n14425) );
  MOAI22 U23339 ( .A1(n28950), .A2(n2662), .B1(ram[10185]), .B2(n2663), 
        .ZN(n14426) );
  MOAI22 U23340 ( .A1(n28715), .A2(n2662), .B1(ram[10186]), .B2(n2663), 
        .ZN(n14427) );
  MOAI22 U23341 ( .A1(n28480), .A2(n2662), .B1(ram[10187]), .B2(n2663), 
        .ZN(n14428) );
  MOAI22 U23342 ( .A1(n28245), .A2(n2662), .B1(ram[10188]), .B2(n2663), 
        .ZN(n14429) );
  MOAI22 U23343 ( .A1(n28010), .A2(n2662), .B1(ram[10189]), .B2(n2663), 
        .ZN(n14430) );
  MOAI22 U23344 ( .A1(n27775), .A2(n2662), .B1(ram[10190]), .B2(n2663), 
        .ZN(n14431) );
  MOAI22 U23345 ( .A1(n27540), .A2(n2662), .B1(ram[10191]), .B2(n2663), 
        .ZN(n14432) );
  MOAI22 U23346 ( .A1(n29186), .A2(n2664), .B1(ram[10192]), .B2(n2665), 
        .ZN(n14433) );
  MOAI22 U23347 ( .A1(n28951), .A2(n2664), .B1(ram[10193]), .B2(n2665), 
        .ZN(n14434) );
  MOAI22 U23348 ( .A1(n28716), .A2(n2664), .B1(ram[10194]), .B2(n2665), 
        .ZN(n14435) );
  MOAI22 U23349 ( .A1(n28481), .A2(n2664), .B1(ram[10195]), .B2(n2665), 
        .ZN(n14436) );
  MOAI22 U23350 ( .A1(n28246), .A2(n2664), .B1(ram[10196]), .B2(n2665), 
        .ZN(n14437) );
  MOAI22 U23351 ( .A1(n28011), .A2(n2664), .B1(ram[10197]), .B2(n2665), 
        .ZN(n14438) );
  MOAI22 U23352 ( .A1(n27776), .A2(n2664), .B1(ram[10198]), .B2(n2665), 
        .ZN(n14439) );
  MOAI22 U23353 ( .A1(n27541), .A2(n2664), .B1(ram[10199]), .B2(n2665), 
        .ZN(n14440) );
  MOAI22 U23354 ( .A1(n29186), .A2(n2666), .B1(ram[10200]), .B2(n2667), 
        .ZN(n14441) );
  MOAI22 U23355 ( .A1(n28951), .A2(n2666), .B1(ram[10201]), .B2(n2667), 
        .ZN(n14442) );
  MOAI22 U23356 ( .A1(n28716), .A2(n2666), .B1(ram[10202]), .B2(n2667), 
        .ZN(n14443) );
  MOAI22 U23357 ( .A1(n28481), .A2(n2666), .B1(ram[10203]), .B2(n2667), 
        .ZN(n14444) );
  MOAI22 U23358 ( .A1(n28246), .A2(n2666), .B1(ram[10204]), .B2(n2667), 
        .ZN(n14445) );
  MOAI22 U23359 ( .A1(n28011), .A2(n2666), .B1(ram[10205]), .B2(n2667), 
        .ZN(n14446) );
  MOAI22 U23360 ( .A1(n27776), .A2(n2666), .B1(ram[10206]), .B2(n2667), 
        .ZN(n14447) );
  MOAI22 U23361 ( .A1(n27541), .A2(n2666), .B1(ram[10207]), .B2(n2667), 
        .ZN(n14448) );
  MOAI22 U23362 ( .A1(n29186), .A2(n2668), .B1(ram[10208]), .B2(n2669), 
        .ZN(n14449) );
  MOAI22 U23363 ( .A1(n28951), .A2(n2668), .B1(ram[10209]), .B2(n2669), 
        .ZN(n14450) );
  MOAI22 U23364 ( .A1(n28716), .A2(n2668), .B1(ram[10210]), .B2(n2669), 
        .ZN(n14451) );
  MOAI22 U23365 ( .A1(n28481), .A2(n2668), .B1(ram[10211]), .B2(n2669), 
        .ZN(n14452) );
  MOAI22 U23366 ( .A1(n28246), .A2(n2668), .B1(ram[10212]), .B2(n2669), 
        .ZN(n14453) );
  MOAI22 U23367 ( .A1(n28011), .A2(n2668), .B1(ram[10213]), .B2(n2669), 
        .ZN(n14454) );
  MOAI22 U23368 ( .A1(n27776), .A2(n2668), .B1(ram[10214]), .B2(n2669), 
        .ZN(n14455) );
  MOAI22 U23369 ( .A1(n27541), .A2(n2668), .B1(ram[10215]), .B2(n2669), 
        .ZN(n14456) );
  MOAI22 U23370 ( .A1(n29186), .A2(n2670), .B1(ram[10216]), .B2(n2671), 
        .ZN(n14457) );
  MOAI22 U23371 ( .A1(n28951), .A2(n2670), .B1(ram[10217]), .B2(n2671), 
        .ZN(n14458) );
  MOAI22 U23372 ( .A1(n28716), .A2(n2670), .B1(ram[10218]), .B2(n2671), 
        .ZN(n14459) );
  MOAI22 U23373 ( .A1(n28481), .A2(n2670), .B1(ram[10219]), .B2(n2671), 
        .ZN(n14460) );
  MOAI22 U23374 ( .A1(n28246), .A2(n2670), .B1(ram[10220]), .B2(n2671), 
        .ZN(n14461) );
  MOAI22 U23375 ( .A1(n28011), .A2(n2670), .B1(ram[10221]), .B2(n2671), 
        .ZN(n14462) );
  MOAI22 U23376 ( .A1(n27776), .A2(n2670), .B1(ram[10222]), .B2(n2671), 
        .ZN(n14463) );
  MOAI22 U23377 ( .A1(n27541), .A2(n2670), .B1(ram[10223]), .B2(n2671), 
        .ZN(n14464) );
  MOAI22 U23378 ( .A1(n29186), .A2(n2672), .B1(ram[10224]), .B2(n2673), 
        .ZN(n14465) );
  MOAI22 U23379 ( .A1(n28951), .A2(n2672), .B1(ram[10225]), .B2(n2673), 
        .ZN(n14466) );
  MOAI22 U23380 ( .A1(n28716), .A2(n2672), .B1(ram[10226]), .B2(n2673), 
        .ZN(n14467) );
  MOAI22 U23381 ( .A1(n28481), .A2(n2672), .B1(ram[10227]), .B2(n2673), 
        .ZN(n14468) );
  MOAI22 U23382 ( .A1(n28246), .A2(n2672), .B1(ram[10228]), .B2(n2673), 
        .ZN(n14469) );
  MOAI22 U23383 ( .A1(n28011), .A2(n2672), .B1(ram[10229]), .B2(n2673), 
        .ZN(n14470) );
  MOAI22 U23384 ( .A1(n27776), .A2(n2672), .B1(ram[10230]), .B2(n2673), 
        .ZN(n14471) );
  MOAI22 U23385 ( .A1(n27541), .A2(n2672), .B1(ram[10231]), .B2(n2673), 
        .ZN(n14472) );
  MOAI22 U23386 ( .A1(n29186), .A2(n2674), .B1(ram[10232]), .B2(n2675), 
        .ZN(n14473) );
  MOAI22 U23387 ( .A1(n28951), .A2(n2674), .B1(ram[10233]), .B2(n2675), 
        .ZN(n14474) );
  MOAI22 U23388 ( .A1(n28716), .A2(n2674), .B1(ram[10234]), .B2(n2675), 
        .ZN(n14475) );
  MOAI22 U23389 ( .A1(n28481), .A2(n2674), .B1(ram[10235]), .B2(n2675), 
        .ZN(n14476) );
  MOAI22 U23390 ( .A1(n28246), .A2(n2674), .B1(ram[10236]), .B2(n2675), 
        .ZN(n14477) );
  MOAI22 U23391 ( .A1(n28011), .A2(n2674), .B1(ram[10237]), .B2(n2675), 
        .ZN(n14478) );
  MOAI22 U23392 ( .A1(n27776), .A2(n2674), .B1(ram[10238]), .B2(n2675), 
        .ZN(n14479) );
  MOAI22 U23393 ( .A1(n27541), .A2(n2674), .B1(ram[10239]), .B2(n2675), 
        .ZN(n14480) );
  MOAI22 U23394 ( .A1(n29186), .A2(n2676), .B1(ram[10240]), .B2(n2677), 
        .ZN(n14481) );
  MOAI22 U23395 ( .A1(n28951), .A2(n2676), .B1(ram[10241]), .B2(n2677), 
        .ZN(n14482) );
  MOAI22 U23396 ( .A1(n28716), .A2(n2676), .B1(ram[10242]), .B2(n2677), 
        .ZN(n14483) );
  MOAI22 U23397 ( .A1(n28481), .A2(n2676), .B1(ram[10243]), .B2(n2677), 
        .ZN(n14484) );
  MOAI22 U23398 ( .A1(n28246), .A2(n2676), .B1(ram[10244]), .B2(n2677), 
        .ZN(n14485) );
  MOAI22 U23399 ( .A1(n28011), .A2(n2676), .B1(ram[10245]), .B2(n2677), 
        .ZN(n14486) );
  MOAI22 U23400 ( .A1(n27776), .A2(n2676), .B1(ram[10246]), .B2(n2677), 
        .ZN(n14487) );
  MOAI22 U23401 ( .A1(n27541), .A2(n2676), .B1(ram[10247]), .B2(n2677), 
        .ZN(n14488) );
  MOAI22 U23402 ( .A1(n29186), .A2(n2679), .B1(ram[10248]), .B2(n2680), 
        .ZN(n14489) );
  MOAI22 U23403 ( .A1(n28951), .A2(n2679), .B1(ram[10249]), .B2(n2680), 
        .ZN(n14490) );
  MOAI22 U23404 ( .A1(n28716), .A2(n2679), .B1(ram[10250]), .B2(n2680), 
        .ZN(n14491) );
  MOAI22 U23405 ( .A1(n28481), .A2(n2679), .B1(ram[10251]), .B2(n2680), 
        .ZN(n14492) );
  MOAI22 U23406 ( .A1(n28246), .A2(n2679), .B1(ram[10252]), .B2(n2680), 
        .ZN(n14493) );
  MOAI22 U23407 ( .A1(n28011), .A2(n2679), .B1(ram[10253]), .B2(n2680), 
        .ZN(n14494) );
  MOAI22 U23408 ( .A1(n27776), .A2(n2679), .B1(ram[10254]), .B2(n2680), 
        .ZN(n14495) );
  MOAI22 U23409 ( .A1(n27541), .A2(n2679), .B1(ram[10255]), .B2(n2680), 
        .ZN(n14496) );
  MOAI22 U23410 ( .A1(n29186), .A2(n2681), .B1(ram[10256]), .B2(n2682), 
        .ZN(n14497) );
  MOAI22 U23411 ( .A1(n28951), .A2(n2681), .B1(ram[10257]), .B2(n2682), 
        .ZN(n14498) );
  MOAI22 U23412 ( .A1(n28716), .A2(n2681), .B1(ram[10258]), .B2(n2682), 
        .ZN(n14499) );
  MOAI22 U23413 ( .A1(n28481), .A2(n2681), .B1(ram[10259]), .B2(n2682), 
        .ZN(n14500) );
  MOAI22 U23414 ( .A1(n28246), .A2(n2681), .B1(ram[10260]), .B2(n2682), 
        .ZN(n14501) );
  MOAI22 U23415 ( .A1(n28011), .A2(n2681), .B1(ram[10261]), .B2(n2682), 
        .ZN(n14502) );
  MOAI22 U23416 ( .A1(n27776), .A2(n2681), .B1(ram[10262]), .B2(n2682), 
        .ZN(n14503) );
  MOAI22 U23417 ( .A1(n27541), .A2(n2681), .B1(ram[10263]), .B2(n2682), 
        .ZN(n14504) );
  MOAI22 U23418 ( .A1(n29186), .A2(n2683), .B1(ram[10264]), .B2(n2684), 
        .ZN(n14505) );
  MOAI22 U23419 ( .A1(n28951), .A2(n2683), .B1(ram[10265]), .B2(n2684), 
        .ZN(n14506) );
  MOAI22 U23420 ( .A1(n28716), .A2(n2683), .B1(ram[10266]), .B2(n2684), 
        .ZN(n14507) );
  MOAI22 U23421 ( .A1(n28481), .A2(n2683), .B1(ram[10267]), .B2(n2684), 
        .ZN(n14508) );
  MOAI22 U23422 ( .A1(n28246), .A2(n2683), .B1(ram[10268]), .B2(n2684), 
        .ZN(n14509) );
  MOAI22 U23423 ( .A1(n28011), .A2(n2683), .B1(ram[10269]), .B2(n2684), 
        .ZN(n14510) );
  MOAI22 U23424 ( .A1(n27776), .A2(n2683), .B1(ram[10270]), .B2(n2684), 
        .ZN(n14511) );
  MOAI22 U23425 ( .A1(n27541), .A2(n2683), .B1(ram[10271]), .B2(n2684), 
        .ZN(n14512) );
  MOAI22 U23426 ( .A1(n29186), .A2(n2685), .B1(ram[10272]), .B2(n2686), 
        .ZN(n14513) );
  MOAI22 U23427 ( .A1(n28951), .A2(n2685), .B1(ram[10273]), .B2(n2686), 
        .ZN(n14514) );
  MOAI22 U23428 ( .A1(n28716), .A2(n2685), .B1(ram[10274]), .B2(n2686), 
        .ZN(n14515) );
  MOAI22 U23429 ( .A1(n28481), .A2(n2685), .B1(ram[10275]), .B2(n2686), 
        .ZN(n14516) );
  MOAI22 U23430 ( .A1(n28246), .A2(n2685), .B1(ram[10276]), .B2(n2686), 
        .ZN(n14517) );
  MOAI22 U23431 ( .A1(n28011), .A2(n2685), .B1(ram[10277]), .B2(n2686), 
        .ZN(n14518) );
  MOAI22 U23432 ( .A1(n27776), .A2(n2685), .B1(ram[10278]), .B2(n2686), 
        .ZN(n14519) );
  MOAI22 U23433 ( .A1(n27541), .A2(n2685), .B1(ram[10279]), .B2(n2686), 
        .ZN(n14520) );
  MOAI22 U23434 ( .A1(n29186), .A2(n2687), .B1(ram[10280]), .B2(n2688), 
        .ZN(n14521) );
  MOAI22 U23435 ( .A1(n28951), .A2(n2687), .B1(ram[10281]), .B2(n2688), 
        .ZN(n14522) );
  MOAI22 U23436 ( .A1(n28716), .A2(n2687), .B1(ram[10282]), .B2(n2688), 
        .ZN(n14523) );
  MOAI22 U23437 ( .A1(n28481), .A2(n2687), .B1(ram[10283]), .B2(n2688), 
        .ZN(n14524) );
  MOAI22 U23438 ( .A1(n28246), .A2(n2687), .B1(ram[10284]), .B2(n2688), 
        .ZN(n14525) );
  MOAI22 U23439 ( .A1(n28011), .A2(n2687), .B1(ram[10285]), .B2(n2688), 
        .ZN(n14526) );
  MOAI22 U23440 ( .A1(n27776), .A2(n2687), .B1(ram[10286]), .B2(n2688), 
        .ZN(n14527) );
  MOAI22 U23441 ( .A1(n27541), .A2(n2687), .B1(ram[10287]), .B2(n2688), 
        .ZN(n14528) );
  MOAI22 U23442 ( .A1(n29186), .A2(n2689), .B1(ram[10288]), .B2(n2690), 
        .ZN(n14529) );
  MOAI22 U23443 ( .A1(n28951), .A2(n2689), .B1(ram[10289]), .B2(n2690), 
        .ZN(n14530) );
  MOAI22 U23444 ( .A1(n28716), .A2(n2689), .B1(ram[10290]), .B2(n2690), 
        .ZN(n14531) );
  MOAI22 U23445 ( .A1(n28481), .A2(n2689), .B1(ram[10291]), .B2(n2690), 
        .ZN(n14532) );
  MOAI22 U23446 ( .A1(n28246), .A2(n2689), .B1(ram[10292]), .B2(n2690), 
        .ZN(n14533) );
  MOAI22 U23447 ( .A1(n28011), .A2(n2689), .B1(ram[10293]), .B2(n2690), 
        .ZN(n14534) );
  MOAI22 U23448 ( .A1(n27776), .A2(n2689), .B1(ram[10294]), .B2(n2690), 
        .ZN(n14535) );
  MOAI22 U23449 ( .A1(n27541), .A2(n2689), .B1(ram[10295]), .B2(n2690), 
        .ZN(n14536) );
  MOAI22 U23450 ( .A1(n29187), .A2(n2691), .B1(ram[10296]), .B2(n2692), 
        .ZN(n14537) );
  MOAI22 U23451 ( .A1(n28952), .A2(n2691), .B1(ram[10297]), .B2(n2692), 
        .ZN(n14538) );
  MOAI22 U23452 ( .A1(n28717), .A2(n2691), .B1(ram[10298]), .B2(n2692), 
        .ZN(n14539) );
  MOAI22 U23453 ( .A1(n28482), .A2(n2691), .B1(ram[10299]), .B2(n2692), 
        .ZN(n14540) );
  MOAI22 U23454 ( .A1(n28247), .A2(n2691), .B1(ram[10300]), .B2(n2692), 
        .ZN(n14541) );
  MOAI22 U23455 ( .A1(n28012), .A2(n2691), .B1(ram[10301]), .B2(n2692), 
        .ZN(n14542) );
  MOAI22 U23456 ( .A1(n27777), .A2(n2691), .B1(ram[10302]), .B2(n2692), 
        .ZN(n14543) );
  MOAI22 U23457 ( .A1(n27542), .A2(n2691), .B1(ram[10303]), .B2(n2692), 
        .ZN(n14544) );
  MOAI22 U23458 ( .A1(n29187), .A2(n2693), .B1(ram[10304]), .B2(n2694), 
        .ZN(n14545) );
  MOAI22 U23459 ( .A1(n28952), .A2(n2693), .B1(ram[10305]), .B2(n2694), 
        .ZN(n14546) );
  MOAI22 U23460 ( .A1(n28717), .A2(n2693), .B1(ram[10306]), .B2(n2694), 
        .ZN(n14547) );
  MOAI22 U23461 ( .A1(n28482), .A2(n2693), .B1(ram[10307]), .B2(n2694), 
        .ZN(n14548) );
  MOAI22 U23462 ( .A1(n28247), .A2(n2693), .B1(ram[10308]), .B2(n2694), 
        .ZN(n14549) );
  MOAI22 U23463 ( .A1(n28012), .A2(n2693), .B1(ram[10309]), .B2(n2694), 
        .ZN(n14550) );
  MOAI22 U23464 ( .A1(n27777), .A2(n2693), .B1(ram[10310]), .B2(n2694), 
        .ZN(n14551) );
  MOAI22 U23465 ( .A1(n27542), .A2(n2693), .B1(ram[10311]), .B2(n2694), 
        .ZN(n14552) );
  MOAI22 U23466 ( .A1(n29187), .A2(n2695), .B1(ram[10312]), .B2(n2696), 
        .ZN(n14553) );
  MOAI22 U23467 ( .A1(n28952), .A2(n2695), .B1(ram[10313]), .B2(n2696), 
        .ZN(n14554) );
  MOAI22 U23468 ( .A1(n28717), .A2(n2695), .B1(ram[10314]), .B2(n2696), 
        .ZN(n14555) );
  MOAI22 U23469 ( .A1(n28482), .A2(n2695), .B1(ram[10315]), .B2(n2696), 
        .ZN(n14556) );
  MOAI22 U23470 ( .A1(n28247), .A2(n2695), .B1(ram[10316]), .B2(n2696), 
        .ZN(n14557) );
  MOAI22 U23471 ( .A1(n28012), .A2(n2695), .B1(ram[10317]), .B2(n2696), 
        .ZN(n14558) );
  MOAI22 U23472 ( .A1(n27777), .A2(n2695), .B1(ram[10318]), .B2(n2696), 
        .ZN(n14559) );
  MOAI22 U23473 ( .A1(n27542), .A2(n2695), .B1(ram[10319]), .B2(n2696), 
        .ZN(n14560) );
  MOAI22 U23474 ( .A1(n29187), .A2(n2697), .B1(ram[10320]), .B2(n2698), 
        .ZN(n14561) );
  MOAI22 U23475 ( .A1(n28952), .A2(n2697), .B1(ram[10321]), .B2(n2698), 
        .ZN(n14562) );
  MOAI22 U23476 ( .A1(n28717), .A2(n2697), .B1(ram[10322]), .B2(n2698), 
        .ZN(n14563) );
  MOAI22 U23477 ( .A1(n28482), .A2(n2697), .B1(ram[10323]), .B2(n2698), 
        .ZN(n14564) );
  MOAI22 U23478 ( .A1(n28247), .A2(n2697), .B1(ram[10324]), .B2(n2698), 
        .ZN(n14565) );
  MOAI22 U23479 ( .A1(n28012), .A2(n2697), .B1(ram[10325]), .B2(n2698), 
        .ZN(n14566) );
  MOAI22 U23480 ( .A1(n27777), .A2(n2697), .B1(ram[10326]), .B2(n2698), 
        .ZN(n14567) );
  MOAI22 U23481 ( .A1(n27542), .A2(n2697), .B1(ram[10327]), .B2(n2698), 
        .ZN(n14568) );
  MOAI22 U23482 ( .A1(n29187), .A2(n2699), .B1(ram[10328]), .B2(n2700), 
        .ZN(n14569) );
  MOAI22 U23483 ( .A1(n28952), .A2(n2699), .B1(ram[10329]), .B2(n2700), 
        .ZN(n14570) );
  MOAI22 U23484 ( .A1(n28717), .A2(n2699), .B1(ram[10330]), .B2(n2700), 
        .ZN(n14571) );
  MOAI22 U23485 ( .A1(n28482), .A2(n2699), .B1(ram[10331]), .B2(n2700), 
        .ZN(n14572) );
  MOAI22 U23486 ( .A1(n28247), .A2(n2699), .B1(ram[10332]), .B2(n2700), 
        .ZN(n14573) );
  MOAI22 U23487 ( .A1(n28012), .A2(n2699), .B1(ram[10333]), .B2(n2700), 
        .ZN(n14574) );
  MOAI22 U23488 ( .A1(n27777), .A2(n2699), .B1(ram[10334]), .B2(n2700), 
        .ZN(n14575) );
  MOAI22 U23489 ( .A1(n27542), .A2(n2699), .B1(ram[10335]), .B2(n2700), 
        .ZN(n14576) );
  MOAI22 U23490 ( .A1(n29187), .A2(n2701), .B1(ram[10336]), .B2(n2702), 
        .ZN(n14577) );
  MOAI22 U23491 ( .A1(n28952), .A2(n2701), .B1(ram[10337]), .B2(n2702), 
        .ZN(n14578) );
  MOAI22 U23492 ( .A1(n28717), .A2(n2701), .B1(ram[10338]), .B2(n2702), 
        .ZN(n14579) );
  MOAI22 U23493 ( .A1(n28482), .A2(n2701), .B1(ram[10339]), .B2(n2702), 
        .ZN(n14580) );
  MOAI22 U23494 ( .A1(n28247), .A2(n2701), .B1(ram[10340]), .B2(n2702), 
        .ZN(n14581) );
  MOAI22 U23495 ( .A1(n28012), .A2(n2701), .B1(ram[10341]), .B2(n2702), 
        .ZN(n14582) );
  MOAI22 U23496 ( .A1(n27777), .A2(n2701), .B1(ram[10342]), .B2(n2702), 
        .ZN(n14583) );
  MOAI22 U23497 ( .A1(n27542), .A2(n2701), .B1(ram[10343]), .B2(n2702), 
        .ZN(n14584) );
  MOAI22 U23498 ( .A1(n29187), .A2(n2703), .B1(ram[10344]), .B2(n2704), 
        .ZN(n14585) );
  MOAI22 U23499 ( .A1(n28952), .A2(n2703), .B1(ram[10345]), .B2(n2704), 
        .ZN(n14586) );
  MOAI22 U23500 ( .A1(n28717), .A2(n2703), .B1(ram[10346]), .B2(n2704), 
        .ZN(n14587) );
  MOAI22 U23501 ( .A1(n28482), .A2(n2703), .B1(ram[10347]), .B2(n2704), 
        .ZN(n14588) );
  MOAI22 U23502 ( .A1(n28247), .A2(n2703), .B1(ram[10348]), .B2(n2704), 
        .ZN(n14589) );
  MOAI22 U23503 ( .A1(n28012), .A2(n2703), .B1(ram[10349]), .B2(n2704), 
        .ZN(n14590) );
  MOAI22 U23504 ( .A1(n27777), .A2(n2703), .B1(ram[10350]), .B2(n2704), 
        .ZN(n14591) );
  MOAI22 U23505 ( .A1(n27542), .A2(n2703), .B1(ram[10351]), .B2(n2704), 
        .ZN(n14592) );
  MOAI22 U23506 ( .A1(n29187), .A2(n2705), .B1(ram[10352]), .B2(n2706), 
        .ZN(n14593) );
  MOAI22 U23507 ( .A1(n28952), .A2(n2705), .B1(ram[10353]), .B2(n2706), 
        .ZN(n14594) );
  MOAI22 U23508 ( .A1(n28717), .A2(n2705), .B1(ram[10354]), .B2(n2706), 
        .ZN(n14595) );
  MOAI22 U23509 ( .A1(n28482), .A2(n2705), .B1(ram[10355]), .B2(n2706), 
        .ZN(n14596) );
  MOAI22 U23510 ( .A1(n28247), .A2(n2705), .B1(ram[10356]), .B2(n2706), 
        .ZN(n14597) );
  MOAI22 U23511 ( .A1(n28012), .A2(n2705), .B1(ram[10357]), .B2(n2706), 
        .ZN(n14598) );
  MOAI22 U23512 ( .A1(n27777), .A2(n2705), .B1(ram[10358]), .B2(n2706), 
        .ZN(n14599) );
  MOAI22 U23513 ( .A1(n27542), .A2(n2705), .B1(ram[10359]), .B2(n2706), 
        .ZN(n14600) );
  MOAI22 U23514 ( .A1(n29187), .A2(n2707), .B1(ram[10360]), .B2(n2708), 
        .ZN(n14601) );
  MOAI22 U23515 ( .A1(n28952), .A2(n2707), .B1(ram[10361]), .B2(n2708), 
        .ZN(n14602) );
  MOAI22 U23516 ( .A1(n28717), .A2(n2707), .B1(ram[10362]), .B2(n2708), 
        .ZN(n14603) );
  MOAI22 U23517 ( .A1(n28482), .A2(n2707), .B1(ram[10363]), .B2(n2708), 
        .ZN(n14604) );
  MOAI22 U23518 ( .A1(n28247), .A2(n2707), .B1(ram[10364]), .B2(n2708), 
        .ZN(n14605) );
  MOAI22 U23519 ( .A1(n28012), .A2(n2707), .B1(ram[10365]), .B2(n2708), 
        .ZN(n14606) );
  MOAI22 U23520 ( .A1(n27777), .A2(n2707), .B1(ram[10366]), .B2(n2708), 
        .ZN(n14607) );
  MOAI22 U23521 ( .A1(n27542), .A2(n2707), .B1(ram[10367]), .B2(n2708), 
        .ZN(n14608) );
  MOAI22 U23522 ( .A1(n29187), .A2(n2709), .B1(ram[10368]), .B2(n2710), 
        .ZN(n14609) );
  MOAI22 U23523 ( .A1(n28952), .A2(n2709), .B1(ram[10369]), .B2(n2710), 
        .ZN(n14610) );
  MOAI22 U23524 ( .A1(n28717), .A2(n2709), .B1(ram[10370]), .B2(n2710), 
        .ZN(n14611) );
  MOAI22 U23525 ( .A1(n28482), .A2(n2709), .B1(ram[10371]), .B2(n2710), 
        .ZN(n14612) );
  MOAI22 U23526 ( .A1(n28247), .A2(n2709), .B1(ram[10372]), .B2(n2710), 
        .ZN(n14613) );
  MOAI22 U23527 ( .A1(n28012), .A2(n2709), .B1(ram[10373]), .B2(n2710), 
        .ZN(n14614) );
  MOAI22 U23528 ( .A1(n27777), .A2(n2709), .B1(ram[10374]), .B2(n2710), 
        .ZN(n14615) );
  MOAI22 U23529 ( .A1(n27542), .A2(n2709), .B1(ram[10375]), .B2(n2710), 
        .ZN(n14616) );
  MOAI22 U23530 ( .A1(n29187), .A2(n2711), .B1(ram[10376]), .B2(n2712), 
        .ZN(n14617) );
  MOAI22 U23531 ( .A1(n28952), .A2(n2711), .B1(ram[10377]), .B2(n2712), 
        .ZN(n14618) );
  MOAI22 U23532 ( .A1(n28717), .A2(n2711), .B1(ram[10378]), .B2(n2712), 
        .ZN(n14619) );
  MOAI22 U23533 ( .A1(n28482), .A2(n2711), .B1(ram[10379]), .B2(n2712), 
        .ZN(n14620) );
  MOAI22 U23534 ( .A1(n28247), .A2(n2711), .B1(ram[10380]), .B2(n2712), 
        .ZN(n14621) );
  MOAI22 U23535 ( .A1(n28012), .A2(n2711), .B1(ram[10381]), .B2(n2712), 
        .ZN(n14622) );
  MOAI22 U23536 ( .A1(n27777), .A2(n2711), .B1(ram[10382]), .B2(n2712), 
        .ZN(n14623) );
  MOAI22 U23537 ( .A1(n27542), .A2(n2711), .B1(ram[10383]), .B2(n2712), 
        .ZN(n14624) );
  MOAI22 U23538 ( .A1(n29187), .A2(n2713), .B1(ram[10384]), .B2(n2714), 
        .ZN(n14625) );
  MOAI22 U23539 ( .A1(n28952), .A2(n2713), .B1(ram[10385]), .B2(n2714), 
        .ZN(n14626) );
  MOAI22 U23540 ( .A1(n28717), .A2(n2713), .B1(ram[10386]), .B2(n2714), 
        .ZN(n14627) );
  MOAI22 U23541 ( .A1(n28482), .A2(n2713), .B1(ram[10387]), .B2(n2714), 
        .ZN(n14628) );
  MOAI22 U23542 ( .A1(n28247), .A2(n2713), .B1(ram[10388]), .B2(n2714), 
        .ZN(n14629) );
  MOAI22 U23543 ( .A1(n28012), .A2(n2713), .B1(ram[10389]), .B2(n2714), 
        .ZN(n14630) );
  MOAI22 U23544 ( .A1(n27777), .A2(n2713), .B1(ram[10390]), .B2(n2714), 
        .ZN(n14631) );
  MOAI22 U23545 ( .A1(n27542), .A2(n2713), .B1(ram[10391]), .B2(n2714), 
        .ZN(n14632) );
  MOAI22 U23546 ( .A1(n29187), .A2(n2715), .B1(ram[10392]), .B2(n2716), 
        .ZN(n14633) );
  MOAI22 U23547 ( .A1(n28952), .A2(n2715), .B1(ram[10393]), .B2(n2716), 
        .ZN(n14634) );
  MOAI22 U23548 ( .A1(n28717), .A2(n2715), .B1(ram[10394]), .B2(n2716), 
        .ZN(n14635) );
  MOAI22 U23549 ( .A1(n28482), .A2(n2715), .B1(ram[10395]), .B2(n2716), 
        .ZN(n14636) );
  MOAI22 U23550 ( .A1(n28247), .A2(n2715), .B1(ram[10396]), .B2(n2716), 
        .ZN(n14637) );
  MOAI22 U23551 ( .A1(n28012), .A2(n2715), .B1(ram[10397]), .B2(n2716), 
        .ZN(n14638) );
  MOAI22 U23552 ( .A1(n27777), .A2(n2715), .B1(ram[10398]), .B2(n2716), 
        .ZN(n14639) );
  MOAI22 U23553 ( .A1(n27542), .A2(n2715), .B1(ram[10399]), .B2(n2716), 
        .ZN(n14640) );
  MOAI22 U23554 ( .A1(n29188), .A2(n2717), .B1(ram[10400]), .B2(n2718), 
        .ZN(n14641) );
  MOAI22 U23555 ( .A1(n28953), .A2(n2717), .B1(ram[10401]), .B2(n2718), 
        .ZN(n14642) );
  MOAI22 U23556 ( .A1(n28718), .A2(n2717), .B1(ram[10402]), .B2(n2718), 
        .ZN(n14643) );
  MOAI22 U23557 ( .A1(n28483), .A2(n2717), .B1(ram[10403]), .B2(n2718), 
        .ZN(n14644) );
  MOAI22 U23558 ( .A1(n28248), .A2(n2717), .B1(ram[10404]), .B2(n2718), 
        .ZN(n14645) );
  MOAI22 U23559 ( .A1(n28013), .A2(n2717), .B1(ram[10405]), .B2(n2718), 
        .ZN(n14646) );
  MOAI22 U23560 ( .A1(n27778), .A2(n2717), .B1(ram[10406]), .B2(n2718), 
        .ZN(n14647) );
  MOAI22 U23561 ( .A1(n27543), .A2(n2717), .B1(ram[10407]), .B2(n2718), 
        .ZN(n14648) );
  MOAI22 U23562 ( .A1(n29188), .A2(n2719), .B1(ram[10408]), .B2(n2720), 
        .ZN(n14649) );
  MOAI22 U23563 ( .A1(n28953), .A2(n2719), .B1(ram[10409]), .B2(n2720), 
        .ZN(n14650) );
  MOAI22 U23564 ( .A1(n28718), .A2(n2719), .B1(ram[10410]), .B2(n2720), 
        .ZN(n14651) );
  MOAI22 U23565 ( .A1(n28483), .A2(n2719), .B1(ram[10411]), .B2(n2720), 
        .ZN(n14652) );
  MOAI22 U23566 ( .A1(n28248), .A2(n2719), .B1(ram[10412]), .B2(n2720), 
        .ZN(n14653) );
  MOAI22 U23567 ( .A1(n28013), .A2(n2719), .B1(ram[10413]), .B2(n2720), 
        .ZN(n14654) );
  MOAI22 U23568 ( .A1(n27778), .A2(n2719), .B1(ram[10414]), .B2(n2720), 
        .ZN(n14655) );
  MOAI22 U23569 ( .A1(n27543), .A2(n2719), .B1(ram[10415]), .B2(n2720), 
        .ZN(n14656) );
  MOAI22 U23570 ( .A1(n29188), .A2(n2721), .B1(ram[10416]), .B2(n2722), 
        .ZN(n14657) );
  MOAI22 U23571 ( .A1(n28953), .A2(n2721), .B1(ram[10417]), .B2(n2722), 
        .ZN(n14658) );
  MOAI22 U23572 ( .A1(n28718), .A2(n2721), .B1(ram[10418]), .B2(n2722), 
        .ZN(n14659) );
  MOAI22 U23573 ( .A1(n28483), .A2(n2721), .B1(ram[10419]), .B2(n2722), 
        .ZN(n14660) );
  MOAI22 U23574 ( .A1(n28248), .A2(n2721), .B1(ram[10420]), .B2(n2722), 
        .ZN(n14661) );
  MOAI22 U23575 ( .A1(n28013), .A2(n2721), .B1(ram[10421]), .B2(n2722), 
        .ZN(n14662) );
  MOAI22 U23576 ( .A1(n27778), .A2(n2721), .B1(ram[10422]), .B2(n2722), 
        .ZN(n14663) );
  MOAI22 U23577 ( .A1(n27543), .A2(n2721), .B1(ram[10423]), .B2(n2722), 
        .ZN(n14664) );
  MOAI22 U23578 ( .A1(n29188), .A2(n2723), .B1(ram[10424]), .B2(n2724), 
        .ZN(n14665) );
  MOAI22 U23579 ( .A1(n28953), .A2(n2723), .B1(ram[10425]), .B2(n2724), 
        .ZN(n14666) );
  MOAI22 U23580 ( .A1(n28718), .A2(n2723), .B1(ram[10426]), .B2(n2724), 
        .ZN(n14667) );
  MOAI22 U23581 ( .A1(n28483), .A2(n2723), .B1(ram[10427]), .B2(n2724), 
        .ZN(n14668) );
  MOAI22 U23582 ( .A1(n28248), .A2(n2723), .B1(ram[10428]), .B2(n2724), 
        .ZN(n14669) );
  MOAI22 U23583 ( .A1(n28013), .A2(n2723), .B1(ram[10429]), .B2(n2724), 
        .ZN(n14670) );
  MOAI22 U23584 ( .A1(n27778), .A2(n2723), .B1(ram[10430]), .B2(n2724), 
        .ZN(n14671) );
  MOAI22 U23585 ( .A1(n27543), .A2(n2723), .B1(ram[10431]), .B2(n2724), 
        .ZN(n14672) );
  MOAI22 U23586 ( .A1(n29188), .A2(n2725), .B1(ram[10432]), .B2(n2726), 
        .ZN(n14673) );
  MOAI22 U23587 ( .A1(n28953), .A2(n2725), .B1(ram[10433]), .B2(n2726), 
        .ZN(n14674) );
  MOAI22 U23588 ( .A1(n28718), .A2(n2725), .B1(ram[10434]), .B2(n2726), 
        .ZN(n14675) );
  MOAI22 U23589 ( .A1(n28483), .A2(n2725), .B1(ram[10435]), .B2(n2726), 
        .ZN(n14676) );
  MOAI22 U23590 ( .A1(n28248), .A2(n2725), .B1(ram[10436]), .B2(n2726), 
        .ZN(n14677) );
  MOAI22 U23591 ( .A1(n28013), .A2(n2725), .B1(ram[10437]), .B2(n2726), 
        .ZN(n14678) );
  MOAI22 U23592 ( .A1(n27778), .A2(n2725), .B1(ram[10438]), .B2(n2726), 
        .ZN(n14679) );
  MOAI22 U23593 ( .A1(n27543), .A2(n2725), .B1(ram[10439]), .B2(n2726), 
        .ZN(n14680) );
  MOAI22 U23594 ( .A1(n29188), .A2(n2727), .B1(ram[10440]), .B2(n2728), 
        .ZN(n14681) );
  MOAI22 U23595 ( .A1(n28953), .A2(n2727), .B1(ram[10441]), .B2(n2728), 
        .ZN(n14682) );
  MOAI22 U23596 ( .A1(n28718), .A2(n2727), .B1(ram[10442]), .B2(n2728), 
        .ZN(n14683) );
  MOAI22 U23597 ( .A1(n28483), .A2(n2727), .B1(ram[10443]), .B2(n2728), 
        .ZN(n14684) );
  MOAI22 U23598 ( .A1(n28248), .A2(n2727), .B1(ram[10444]), .B2(n2728), 
        .ZN(n14685) );
  MOAI22 U23599 ( .A1(n28013), .A2(n2727), .B1(ram[10445]), .B2(n2728), 
        .ZN(n14686) );
  MOAI22 U23600 ( .A1(n27778), .A2(n2727), .B1(ram[10446]), .B2(n2728), 
        .ZN(n14687) );
  MOAI22 U23601 ( .A1(n27543), .A2(n2727), .B1(ram[10447]), .B2(n2728), 
        .ZN(n14688) );
  MOAI22 U23602 ( .A1(n29188), .A2(n2729), .B1(ram[10448]), .B2(n2730), 
        .ZN(n14689) );
  MOAI22 U23603 ( .A1(n28953), .A2(n2729), .B1(ram[10449]), .B2(n2730), 
        .ZN(n14690) );
  MOAI22 U23604 ( .A1(n28718), .A2(n2729), .B1(ram[10450]), .B2(n2730), 
        .ZN(n14691) );
  MOAI22 U23605 ( .A1(n28483), .A2(n2729), .B1(ram[10451]), .B2(n2730), 
        .ZN(n14692) );
  MOAI22 U23606 ( .A1(n28248), .A2(n2729), .B1(ram[10452]), .B2(n2730), 
        .ZN(n14693) );
  MOAI22 U23607 ( .A1(n28013), .A2(n2729), .B1(ram[10453]), .B2(n2730), 
        .ZN(n14694) );
  MOAI22 U23608 ( .A1(n27778), .A2(n2729), .B1(ram[10454]), .B2(n2730), 
        .ZN(n14695) );
  MOAI22 U23609 ( .A1(n27543), .A2(n2729), .B1(ram[10455]), .B2(n2730), 
        .ZN(n14696) );
  MOAI22 U23610 ( .A1(n29188), .A2(n2731), .B1(ram[10456]), .B2(n2732), 
        .ZN(n14697) );
  MOAI22 U23611 ( .A1(n28953), .A2(n2731), .B1(ram[10457]), .B2(n2732), 
        .ZN(n14698) );
  MOAI22 U23612 ( .A1(n28718), .A2(n2731), .B1(ram[10458]), .B2(n2732), 
        .ZN(n14699) );
  MOAI22 U23613 ( .A1(n28483), .A2(n2731), .B1(ram[10459]), .B2(n2732), 
        .ZN(n14700) );
  MOAI22 U23614 ( .A1(n28248), .A2(n2731), .B1(ram[10460]), .B2(n2732), 
        .ZN(n14701) );
  MOAI22 U23615 ( .A1(n28013), .A2(n2731), .B1(ram[10461]), .B2(n2732), 
        .ZN(n14702) );
  MOAI22 U23616 ( .A1(n27778), .A2(n2731), .B1(ram[10462]), .B2(n2732), 
        .ZN(n14703) );
  MOAI22 U23617 ( .A1(n27543), .A2(n2731), .B1(ram[10463]), .B2(n2732), 
        .ZN(n14704) );
  MOAI22 U23618 ( .A1(n29188), .A2(n2733), .B1(ram[10464]), .B2(n2734), 
        .ZN(n14705) );
  MOAI22 U23619 ( .A1(n28953), .A2(n2733), .B1(ram[10465]), .B2(n2734), 
        .ZN(n14706) );
  MOAI22 U23620 ( .A1(n28718), .A2(n2733), .B1(ram[10466]), .B2(n2734), 
        .ZN(n14707) );
  MOAI22 U23621 ( .A1(n28483), .A2(n2733), .B1(ram[10467]), .B2(n2734), 
        .ZN(n14708) );
  MOAI22 U23622 ( .A1(n28248), .A2(n2733), .B1(ram[10468]), .B2(n2734), 
        .ZN(n14709) );
  MOAI22 U23623 ( .A1(n28013), .A2(n2733), .B1(ram[10469]), .B2(n2734), 
        .ZN(n14710) );
  MOAI22 U23624 ( .A1(n27778), .A2(n2733), .B1(ram[10470]), .B2(n2734), 
        .ZN(n14711) );
  MOAI22 U23625 ( .A1(n27543), .A2(n2733), .B1(ram[10471]), .B2(n2734), 
        .ZN(n14712) );
  MOAI22 U23626 ( .A1(n29188), .A2(n2735), .B1(ram[10472]), .B2(n2736), 
        .ZN(n14713) );
  MOAI22 U23627 ( .A1(n28953), .A2(n2735), .B1(ram[10473]), .B2(n2736), 
        .ZN(n14714) );
  MOAI22 U23628 ( .A1(n28718), .A2(n2735), .B1(ram[10474]), .B2(n2736), 
        .ZN(n14715) );
  MOAI22 U23629 ( .A1(n28483), .A2(n2735), .B1(ram[10475]), .B2(n2736), 
        .ZN(n14716) );
  MOAI22 U23630 ( .A1(n28248), .A2(n2735), .B1(ram[10476]), .B2(n2736), 
        .ZN(n14717) );
  MOAI22 U23631 ( .A1(n28013), .A2(n2735), .B1(ram[10477]), .B2(n2736), 
        .ZN(n14718) );
  MOAI22 U23632 ( .A1(n27778), .A2(n2735), .B1(ram[10478]), .B2(n2736), 
        .ZN(n14719) );
  MOAI22 U23633 ( .A1(n27543), .A2(n2735), .B1(ram[10479]), .B2(n2736), 
        .ZN(n14720) );
  MOAI22 U23634 ( .A1(n29188), .A2(n2737), .B1(ram[10480]), .B2(n2738), 
        .ZN(n14721) );
  MOAI22 U23635 ( .A1(n28953), .A2(n2737), .B1(ram[10481]), .B2(n2738), 
        .ZN(n14722) );
  MOAI22 U23636 ( .A1(n28718), .A2(n2737), .B1(ram[10482]), .B2(n2738), 
        .ZN(n14723) );
  MOAI22 U23637 ( .A1(n28483), .A2(n2737), .B1(ram[10483]), .B2(n2738), 
        .ZN(n14724) );
  MOAI22 U23638 ( .A1(n28248), .A2(n2737), .B1(ram[10484]), .B2(n2738), 
        .ZN(n14725) );
  MOAI22 U23639 ( .A1(n28013), .A2(n2737), .B1(ram[10485]), .B2(n2738), 
        .ZN(n14726) );
  MOAI22 U23640 ( .A1(n27778), .A2(n2737), .B1(ram[10486]), .B2(n2738), 
        .ZN(n14727) );
  MOAI22 U23641 ( .A1(n27543), .A2(n2737), .B1(ram[10487]), .B2(n2738), 
        .ZN(n14728) );
  MOAI22 U23642 ( .A1(n29188), .A2(n2739), .B1(ram[10488]), .B2(n2740), 
        .ZN(n14729) );
  MOAI22 U23643 ( .A1(n28953), .A2(n2739), .B1(ram[10489]), .B2(n2740), 
        .ZN(n14730) );
  MOAI22 U23644 ( .A1(n28718), .A2(n2739), .B1(ram[10490]), .B2(n2740), 
        .ZN(n14731) );
  MOAI22 U23645 ( .A1(n28483), .A2(n2739), .B1(ram[10491]), .B2(n2740), 
        .ZN(n14732) );
  MOAI22 U23646 ( .A1(n28248), .A2(n2739), .B1(ram[10492]), .B2(n2740), 
        .ZN(n14733) );
  MOAI22 U23647 ( .A1(n28013), .A2(n2739), .B1(ram[10493]), .B2(n2740), 
        .ZN(n14734) );
  MOAI22 U23648 ( .A1(n27778), .A2(n2739), .B1(ram[10494]), .B2(n2740), 
        .ZN(n14735) );
  MOAI22 U23649 ( .A1(n27543), .A2(n2739), .B1(ram[10495]), .B2(n2740), 
        .ZN(n14736) );
  MOAI22 U23650 ( .A1(n29188), .A2(n2741), .B1(ram[10496]), .B2(n2742), 
        .ZN(n14737) );
  MOAI22 U23651 ( .A1(n28953), .A2(n2741), .B1(ram[10497]), .B2(n2742), 
        .ZN(n14738) );
  MOAI22 U23652 ( .A1(n28718), .A2(n2741), .B1(ram[10498]), .B2(n2742), 
        .ZN(n14739) );
  MOAI22 U23653 ( .A1(n28483), .A2(n2741), .B1(ram[10499]), .B2(n2742), 
        .ZN(n14740) );
  MOAI22 U23654 ( .A1(n28248), .A2(n2741), .B1(ram[10500]), .B2(n2742), 
        .ZN(n14741) );
  MOAI22 U23655 ( .A1(n28013), .A2(n2741), .B1(ram[10501]), .B2(n2742), 
        .ZN(n14742) );
  MOAI22 U23656 ( .A1(n27778), .A2(n2741), .B1(ram[10502]), .B2(n2742), 
        .ZN(n14743) );
  MOAI22 U23657 ( .A1(n27543), .A2(n2741), .B1(ram[10503]), .B2(n2742), 
        .ZN(n14744) );
  MOAI22 U23658 ( .A1(n29189), .A2(n2743), .B1(ram[10504]), .B2(n2744), 
        .ZN(n14745) );
  MOAI22 U23659 ( .A1(n28954), .A2(n2743), .B1(ram[10505]), .B2(n2744), 
        .ZN(n14746) );
  MOAI22 U23660 ( .A1(n28719), .A2(n2743), .B1(ram[10506]), .B2(n2744), 
        .ZN(n14747) );
  MOAI22 U23661 ( .A1(n28484), .A2(n2743), .B1(ram[10507]), .B2(n2744), 
        .ZN(n14748) );
  MOAI22 U23662 ( .A1(n28249), .A2(n2743), .B1(ram[10508]), .B2(n2744), 
        .ZN(n14749) );
  MOAI22 U23663 ( .A1(n28014), .A2(n2743), .B1(ram[10509]), .B2(n2744), 
        .ZN(n14750) );
  MOAI22 U23664 ( .A1(n27779), .A2(n2743), .B1(ram[10510]), .B2(n2744), 
        .ZN(n14751) );
  MOAI22 U23665 ( .A1(n27544), .A2(n2743), .B1(ram[10511]), .B2(n2744), 
        .ZN(n14752) );
  MOAI22 U23666 ( .A1(n29189), .A2(n2745), .B1(ram[10512]), .B2(n2746), 
        .ZN(n14753) );
  MOAI22 U23667 ( .A1(n28954), .A2(n2745), .B1(ram[10513]), .B2(n2746), 
        .ZN(n14754) );
  MOAI22 U23668 ( .A1(n28719), .A2(n2745), .B1(ram[10514]), .B2(n2746), 
        .ZN(n14755) );
  MOAI22 U23669 ( .A1(n28484), .A2(n2745), .B1(ram[10515]), .B2(n2746), 
        .ZN(n14756) );
  MOAI22 U23670 ( .A1(n28249), .A2(n2745), .B1(ram[10516]), .B2(n2746), 
        .ZN(n14757) );
  MOAI22 U23671 ( .A1(n28014), .A2(n2745), .B1(ram[10517]), .B2(n2746), 
        .ZN(n14758) );
  MOAI22 U23672 ( .A1(n27779), .A2(n2745), .B1(ram[10518]), .B2(n2746), 
        .ZN(n14759) );
  MOAI22 U23673 ( .A1(n27544), .A2(n2745), .B1(ram[10519]), .B2(n2746), 
        .ZN(n14760) );
  MOAI22 U23674 ( .A1(n29189), .A2(n2747), .B1(ram[10520]), .B2(n2748), 
        .ZN(n14761) );
  MOAI22 U23675 ( .A1(n28954), .A2(n2747), .B1(ram[10521]), .B2(n2748), 
        .ZN(n14762) );
  MOAI22 U23676 ( .A1(n28719), .A2(n2747), .B1(ram[10522]), .B2(n2748), 
        .ZN(n14763) );
  MOAI22 U23677 ( .A1(n28484), .A2(n2747), .B1(ram[10523]), .B2(n2748), 
        .ZN(n14764) );
  MOAI22 U23678 ( .A1(n28249), .A2(n2747), .B1(ram[10524]), .B2(n2748), 
        .ZN(n14765) );
  MOAI22 U23679 ( .A1(n28014), .A2(n2747), .B1(ram[10525]), .B2(n2748), 
        .ZN(n14766) );
  MOAI22 U23680 ( .A1(n27779), .A2(n2747), .B1(ram[10526]), .B2(n2748), 
        .ZN(n14767) );
  MOAI22 U23681 ( .A1(n27544), .A2(n2747), .B1(ram[10527]), .B2(n2748), 
        .ZN(n14768) );
  MOAI22 U23682 ( .A1(n29189), .A2(n2749), .B1(ram[10528]), .B2(n2750), 
        .ZN(n14769) );
  MOAI22 U23683 ( .A1(n28954), .A2(n2749), .B1(ram[10529]), .B2(n2750), 
        .ZN(n14770) );
  MOAI22 U23684 ( .A1(n28719), .A2(n2749), .B1(ram[10530]), .B2(n2750), 
        .ZN(n14771) );
  MOAI22 U23685 ( .A1(n28484), .A2(n2749), .B1(ram[10531]), .B2(n2750), 
        .ZN(n14772) );
  MOAI22 U23686 ( .A1(n28249), .A2(n2749), .B1(ram[10532]), .B2(n2750), 
        .ZN(n14773) );
  MOAI22 U23687 ( .A1(n28014), .A2(n2749), .B1(ram[10533]), .B2(n2750), 
        .ZN(n14774) );
  MOAI22 U23688 ( .A1(n27779), .A2(n2749), .B1(ram[10534]), .B2(n2750), 
        .ZN(n14775) );
  MOAI22 U23689 ( .A1(n27544), .A2(n2749), .B1(ram[10535]), .B2(n2750), 
        .ZN(n14776) );
  MOAI22 U23690 ( .A1(n29189), .A2(n2751), .B1(ram[10536]), .B2(n2752), 
        .ZN(n14777) );
  MOAI22 U23691 ( .A1(n28954), .A2(n2751), .B1(ram[10537]), .B2(n2752), 
        .ZN(n14778) );
  MOAI22 U23692 ( .A1(n28719), .A2(n2751), .B1(ram[10538]), .B2(n2752), 
        .ZN(n14779) );
  MOAI22 U23693 ( .A1(n28484), .A2(n2751), .B1(ram[10539]), .B2(n2752), 
        .ZN(n14780) );
  MOAI22 U23694 ( .A1(n28249), .A2(n2751), .B1(ram[10540]), .B2(n2752), 
        .ZN(n14781) );
  MOAI22 U23695 ( .A1(n28014), .A2(n2751), .B1(ram[10541]), .B2(n2752), 
        .ZN(n14782) );
  MOAI22 U23696 ( .A1(n27779), .A2(n2751), .B1(ram[10542]), .B2(n2752), 
        .ZN(n14783) );
  MOAI22 U23697 ( .A1(n27544), .A2(n2751), .B1(ram[10543]), .B2(n2752), 
        .ZN(n14784) );
  MOAI22 U23698 ( .A1(n29189), .A2(n2753), .B1(ram[10544]), .B2(n2754), 
        .ZN(n14785) );
  MOAI22 U23699 ( .A1(n28954), .A2(n2753), .B1(ram[10545]), .B2(n2754), 
        .ZN(n14786) );
  MOAI22 U23700 ( .A1(n28719), .A2(n2753), .B1(ram[10546]), .B2(n2754), 
        .ZN(n14787) );
  MOAI22 U23701 ( .A1(n28484), .A2(n2753), .B1(ram[10547]), .B2(n2754), 
        .ZN(n14788) );
  MOAI22 U23702 ( .A1(n28249), .A2(n2753), .B1(ram[10548]), .B2(n2754), 
        .ZN(n14789) );
  MOAI22 U23703 ( .A1(n28014), .A2(n2753), .B1(ram[10549]), .B2(n2754), 
        .ZN(n14790) );
  MOAI22 U23704 ( .A1(n27779), .A2(n2753), .B1(ram[10550]), .B2(n2754), 
        .ZN(n14791) );
  MOAI22 U23705 ( .A1(n27544), .A2(n2753), .B1(ram[10551]), .B2(n2754), 
        .ZN(n14792) );
  MOAI22 U23706 ( .A1(n29189), .A2(n2755), .B1(ram[10552]), .B2(n2756), 
        .ZN(n14793) );
  MOAI22 U23707 ( .A1(n28954), .A2(n2755), .B1(ram[10553]), .B2(n2756), 
        .ZN(n14794) );
  MOAI22 U23708 ( .A1(n28719), .A2(n2755), .B1(ram[10554]), .B2(n2756), 
        .ZN(n14795) );
  MOAI22 U23709 ( .A1(n28484), .A2(n2755), .B1(ram[10555]), .B2(n2756), 
        .ZN(n14796) );
  MOAI22 U23710 ( .A1(n28249), .A2(n2755), .B1(ram[10556]), .B2(n2756), 
        .ZN(n14797) );
  MOAI22 U23711 ( .A1(n28014), .A2(n2755), .B1(ram[10557]), .B2(n2756), 
        .ZN(n14798) );
  MOAI22 U23712 ( .A1(n27779), .A2(n2755), .B1(ram[10558]), .B2(n2756), 
        .ZN(n14799) );
  MOAI22 U23713 ( .A1(n27544), .A2(n2755), .B1(ram[10559]), .B2(n2756), 
        .ZN(n14800) );
  MOAI22 U23714 ( .A1(n29189), .A2(n2757), .B1(ram[10560]), .B2(n2758), 
        .ZN(n14801) );
  MOAI22 U23715 ( .A1(n28954), .A2(n2757), .B1(ram[10561]), .B2(n2758), 
        .ZN(n14802) );
  MOAI22 U23716 ( .A1(n28719), .A2(n2757), .B1(ram[10562]), .B2(n2758), 
        .ZN(n14803) );
  MOAI22 U23717 ( .A1(n28484), .A2(n2757), .B1(ram[10563]), .B2(n2758), 
        .ZN(n14804) );
  MOAI22 U23718 ( .A1(n28249), .A2(n2757), .B1(ram[10564]), .B2(n2758), 
        .ZN(n14805) );
  MOAI22 U23719 ( .A1(n28014), .A2(n2757), .B1(ram[10565]), .B2(n2758), 
        .ZN(n14806) );
  MOAI22 U23720 ( .A1(n27779), .A2(n2757), .B1(ram[10566]), .B2(n2758), 
        .ZN(n14807) );
  MOAI22 U23721 ( .A1(n27544), .A2(n2757), .B1(ram[10567]), .B2(n2758), 
        .ZN(n14808) );
  MOAI22 U23722 ( .A1(n29189), .A2(n2759), .B1(ram[10568]), .B2(n2760), 
        .ZN(n14809) );
  MOAI22 U23723 ( .A1(n28954), .A2(n2759), .B1(ram[10569]), .B2(n2760), 
        .ZN(n14810) );
  MOAI22 U23724 ( .A1(n28719), .A2(n2759), .B1(ram[10570]), .B2(n2760), 
        .ZN(n14811) );
  MOAI22 U23725 ( .A1(n28484), .A2(n2759), .B1(ram[10571]), .B2(n2760), 
        .ZN(n14812) );
  MOAI22 U23726 ( .A1(n28249), .A2(n2759), .B1(ram[10572]), .B2(n2760), 
        .ZN(n14813) );
  MOAI22 U23727 ( .A1(n28014), .A2(n2759), .B1(ram[10573]), .B2(n2760), 
        .ZN(n14814) );
  MOAI22 U23728 ( .A1(n27779), .A2(n2759), .B1(ram[10574]), .B2(n2760), 
        .ZN(n14815) );
  MOAI22 U23729 ( .A1(n27544), .A2(n2759), .B1(ram[10575]), .B2(n2760), 
        .ZN(n14816) );
  MOAI22 U23730 ( .A1(n29189), .A2(n2761), .B1(ram[10576]), .B2(n2762), 
        .ZN(n14817) );
  MOAI22 U23731 ( .A1(n28954), .A2(n2761), .B1(ram[10577]), .B2(n2762), 
        .ZN(n14818) );
  MOAI22 U23732 ( .A1(n28719), .A2(n2761), .B1(ram[10578]), .B2(n2762), 
        .ZN(n14819) );
  MOAI22 U23733 ( .A1(n28484), .A2(n2761), .B1(ram[10579]), .B2(n2762), 
        .ZN(n14820) );
  MOAI22 U23734 ( .A1(n28249), .A2(n2761), .B1(ram[10580]), .B2(n2762), 
        .ZN(n14821) );
  MOAI22 U23735 ( .A1(n28014), .A2(n2761), .B1(ram[10581]), .B2(n2762), 
        .ZN(n14822) );
  MOAI22 U23736 ( .A1(n27779), .A2(n2761), .B1(ram[10582]), .B2(n2762), 
        .ZN(n14823) );
  MOAI22 U23737 ( .A1(n27544), .A2(n2761), .B1(ram[10583]), .B2(n2762), 
        .ZN(n14824) );
  MOAI22 U23738 ( .A1(n29189), .A2(n2763), .B1(ram[10584]), .B2(n2764), 
        .ZN(n14825) );
  MOAI22 U23739 ( .A1(n28954), .A2(n2763), .B1(ram[10585]), .B2(n2764), 
        .ZN(n14826) );
  MOAI22 U23740 ( .A1(n28719), .A2(n2763), .B1(ram[10586]), .B2(n2764), 
        .ZN(n14827) );
  MOAI22 U23741 ( .A1(n28484), .A2(n2763), .B1(ram[10587]), .B2(n2764), 
        .ZN(n14828) );
  MOAI22 U23742 ( .A1(n28249), .A2(n2763), .B1(ram[10588]), .B2(n2764), 
        .ZN(n14829) );
  MOAI22 U23743 ( .A1(n28014), .A2(n2763), .B1(ram[10589]), .B2(n2764), 
        .ZN(n14830) );
  MOAI22 U23744 ( .A1(n27779), .A2(n2763), .B1(ram[10590]), .B2(n2764), 
        .ZN(n14831) );
  MOAI22 U23745 ( .A1(n27544), .A2(n2763), .B1(ram[10591]), .B2(n2764), 
        .ZN(n14832) );
  MOAI22 U23746 ( .A1(n29189), .A2(n2765), .B1(ram[10592]), .B2(n2766), 
        .ZN(n14833) );
  MOAI22 U23747 ( .A1(n28954), .A2(n2765), .B1(ram[10593]), .B2(n2766), 
        .ZN(n14834) );
  MOAI22 U23748 ( .A1(n28719), .A2(n2765), .B1(ram[10594]), .B2(n2766), 
        .ZN(n14835) );
  MOAI22 U23749 ( .A1(n28484), .A2(n2765), .B1(ram[10595]), .B2(n2766), 
        .ZN(n14836) );
  MOAI22 U23750 ( .A1(n28249), .A2(n2765), .B1(ram[10596]), .B2(n2766), 
        .ZN(n14837) );
  MOAI22 U23751 ( .A1(n28014), .A2(n2765), .B1(ram[10597]), .B2(n2766), 
        .ZN(n14838) );
  MOAI22 U23752 ( .A1(n27779), .A2(n2765), .B1(ram[10598]), .B2(n2766), 
        .ZN(n14839) );
  MOAI22 U23753 ( .A1(n27544), .A2(n2765), .B1(ram[10599]), .B2(n2766), 
        .ZN(n14840) );
  MOAI22 U23754 ( .A1(n29189), .A2(n2767), .B1(ram[10600]), .B2(n2768), 
        .ZN(n14841) );
  MOAI22 U23755 ( .A1(n28954), .A2(n2767), .B1(ram[10601]), .B2(n2768), 
        .ZN(n14842) );
  MOAI22 U23756 ( .A1(n28719), .A2(n2767), .B1(ram[10602]), .B2(n2768), 
        .ZN(n14843) );
  MOAI22 U23757 ( .A1(n28484), .A2(n2767), .B1(ram[10603]), .B2(n2768), 
        .ZN(n14844) );
  MOAI22 U23758 ( .A1(n28249), .A2(n2767), .B1(ram[10604]), .B2(n2768), 
        .ZN(n14845) );
  MOAI22 U23759 ( .A1(n28014), .A2(n2767), .B1(ram[10605]), .B2(n2768), 
        .ZN(n14846) );
  MOAI22 U23760 ( .A1(n27779), .A2(n2767), .B1(ram[10606]), .B2(n2768), 
        .ZN(n14847) );
  MOAI22 U23761 ( .A1(n27544), .A2(n2767), .B1(ram[10607]), .B2(n2768), 
        .ZN(n14848) );
  MOAI22 U23762 ( .A1(n29190), .A2(n2769), .B1(ram[10608]), .B2(n2770), 
        .ZN(n14849) );
  MOAI22 U23763 ( .A1(n28955), .A2(n2769), .B1(ram[10609]), .B2(n2770), 
        .ZN(n14850) );
  MOAI22 U23764 ( .A1(n28720), .A2(n2769), .B1(ram[10610]), .B2(n2770), 
        .ZN(n14851) );
  MOAI22 U23765 ( .A1(n28485), .A2(n2769), .B1(ram[10611]), .B2(n2770), 
        .ZN(n14852) );
  MOAI22 U23766 ( .A1(n28250), .A2(n2769), .B1(ram[10612]), .B2(n2770), 
        .ZN(n14853) );
  MOAI22 U23767 ( .A1(n28015), .A2(n2769), .B1(ram[10613]), .B2(n2770), 
        .ZN(n14854) );
  MOAI22 U23768 ( .A1(n27780), .A2(n2769), .B1(ram[10614]), .B2(n2770), 
        .ZN(n14855) );
  MOAI22 U23769 ( .A1(n27545), .A2(n2769), .B1(ram[10615]), .B2(n2770), 
        .ZN(n14856) );
  MOAI22 U23770 ( .A1(n29190), .A2(n2771), .B1(ram[10616]), .B2(n2772), 
        .ZN(n14857) );
  MOAI22 U23771 ( .A1(n28955), .A2(n2771), .B1(ram[10617]), .B2(n2772), 
        .ZN(n14858) );
  MOAI22 U23772 ( .A1(n28720), .A2(n2771), .B1(ram[10618]), .B2(n2772), 
        .ZN(n14859) );
  MOAI22 U23773 ( .A1(n28485), .A2(n2771), .B1(ram[10619]), .B2(n2772), 
        .ZN(n14860) );
  MOAI22 U23774 ( .A1(n28250), .A2(n2771), .B1(ram[10620]), .B2(n2772), 
        .ZN(n14861) );
  MOAI22 U23775 ( .A1(n28015), .A2(n2771), .B1(ram[10621]), .B2(n2772), 
        .ZN(n14862) );
  MOAI22 U23776 ( .A1(n27780), .A2(n2771), .B1(ram[10622]), .B2(n2772), 
        .ZN(n14863) );
  MOAI22 U23777 ( .A1(n27545), .A2(n2771), .B1(ram[10623]), .B2(n2772), 
        .ZN(n14864) );
  MOAI22 U23778 ( .A1(n29190), .A2(n2773), .B1(ram[10624]), .B2(n2774), 
        .ZN(n14865) );
  MOAI22 U23779 ( .A1(n28955), .A2(n2773), .B1(ram[10625]), .B2(n2774), 
        .ZN(n14866) );
  MOAI22 U23780 ( .A1(n28720), .A2(n2773), .B1(ram[10626]), .B2(n2774), 
        .ZN(n14867) );
  MOAI22 U23781 ( .A1(n28485), .A2(n2773), .B1(ram[10627]), .B2(n2774), 
        .ZN(n14868) );
  MOAI22 U23782 ( .A1(n28250), .A2(n2773), .B1(ram[10628]), .B2(n2774), 
        .ZN(n14869) );
  MOAI22 U23783 ( .A1(n28015), .A2(n2773), .B1(ram[10629]), .B2(n2774), 
        .ZN(n14870) );
  MOAI22 U23784 ( .A1(n27780), .A2(n2773), .B1(ram[10630]), .B2(n2774), 
        .ZN(n14871) );
  MOAI22 U23785 ( .A1(n27545), .A2(n2773), .B1(ram[10631]), .B2(n2774), 
        .ZN(n14872) );
  MOAI22 U23786 ( .A1(n29190), .A2(n2775), .B1(ram[10632]), .B2(n2776), 
        .ZN(n14873) );
  MOAI22 U23787 ( .A1(n28955), .A2(n2775), .B1(ram[10633]), .B2(n2776), 
        .ZN(n14874) );
  MOAI22 U23788 ( .A1(n28720), .A2(n2775), .B1(ram[10634]), .B2(n2776), 
        .ZN(n14875) );
  MOAI22 U23789 ( .A1(n28485), .A2(n2775), .B1(ram[10635]), .B2(n2776), 
        .ZN(n14876) );
  MOAI22 U23790 ( .A1(n28250), .A2(n2775), .B1(ram[10636]), .B2(n2776), 
        .ZN(n14877) );
  MOAI22 U23791 ( .A1(n28015), .A2(n2775), .B1(ram[10637]), .B2(n2776), 
        .ZN(n14878) );
  MOAI22 U23792 ( .A1(n27780), .A2(n2775), .B1(ram[10638]), .B2(n2776), 
        .ZN(n14879) );
  MOAI22 U23793 ( .A1(n27545), .A2(n2775), .B1(ram[10639]), .B2(n2776), 
        .ZN(n14880) );
  MOAI22 U23794 ( .A1(n29190), .A2(n2777), .B1(ram[10640]), .B2(n2778), 
        .ZN(n14881) );
  MOAI22 U23795 ( .A1(n28955), .A2(n2777), .B1(ram[10641]), .B2(n2778), 
        .ZN(n14882) );
  MOAI22 U23796 ( .A1(n28720), .A2(n2777), .B1(ram[10642]), .B2(n2778), 
        .ZN(n14883) );
  MOAI22 U23797 ( .A1(n28485), .A2(n2777), .B1(ram[10643]), .B2(n2778), 
        .ZN(n14884) );
  MOAI22 U23798 ( .A1(n28250), .A2(n2777), .B1(ram[10644]), .B2(n2778), 
        .ZN(n14885) );
  MOAI22 U23799 ( .A1(n28015), .A2(n2777), .B1(ram[10645]), .B2(n2778), 
        .ZN(n14886) );
  MOAI22 U23800 ( .A1(n27780), .A2(n2777), .B1(ram[10646]), .B2(n2778), 
        .ZN(n14887) );
  MOAI22 U23801 ( .A1(n27545), .A2(n2777), .B1(ram[10647]), .B2(n2778), 
        .ZN(n14888) );
  MOAI22 U23802 ( .A1(n29190), .A2(n2779), .B1(ram[10648]), .B2(n2780), 
        .ZN(n14889) );
  MOAI22 U23803 ( .A1(n28955), .A2(n2779), .B1(ram[10649]), .B2(n2780), 
        .ZN(n14890) );
  MOAI22 U23804 ( .A1(n28720), .A2(n2779), .B1(ram[10650]), .B2(n2780), 
        .ZN(n14891) );
  MOAI22 U23805 ( .A1(n28485), .A2(n2779), .B1(ram[10651]), .B2(n2780), 
        .ZN(n14892) );
  MOAI22 U23806 ( .A1(n28250), .A2(n2779), .B1(ram[10652]), .B2(n2780), 
        .ZN(n14893) );
  MOAI22 U23807 ( .A1(n28015), .A2(n2779), .B1(ram[10653]), .B2(n2780), 
        .ZN(n14894) );
  MOAI22 U23808 ( .A1(n27780), .A2(n2779), .B1(ram[10654]), .B2(n2780), 
        .ZN(n14895) );
  MOAI22 U23809 ( .A1(n27545), .A2(n2779), .B1(ram[10655]), .B2(n2780), 
        .ZN(n14896) );
  MOAI22 U23810 ( .A1(n29190), .A2(n2781), .B1(ram[10656]), .B2(n2782), 
        .ZN(n14897) );
  MOAI22 U23811 ( .A1(n28955), .A2(n2781), .B1(ram[10657]), .B2(n2782), 
        .ZN(n14898) );
  MOAI22 U23812 ( .A1(n28720), .A2(n2781), .B1(ram[10658]), .B2(n2782), 
        .ZN(n14899) );
  MOAI22 U23813 ( .A1(n28485), .A2(n2781), .B1(ram[10659]), .B2(n2782), 
        .ZN(n14900) );
  MOAI22 U23814 ( .A1(n28250), .A2(n2781), .B1(ram[10660]), .B2(n2782), 
        .ZN(n14901) );
  MOAI22 U23815 ( .A1(n28015), .A2(n2781), .B1(ram[10661]), .B2(n2782), 
        .ZN(n14902) );
  MOAI22 U23816 ( .A1(n27780), .A2(n2781), .B1(ram[10662]), .B2(n2782), 
        .ZN(n14903) );
  MOAI22 U23817 ( .A1(n27545), .A2(n2781), .B1(ram[10663]), .B2(n2782), 
        .ZN(n14904) );
  MOAI22 U23818 ( .A1(n29190), .A2(n2783), .B1(ram[10664]), .B2(n2784), 
        .ZN(n14905) );
  MOAI22 U23819 ( .A1(n28955), .A2(n2783), .B1(ram[10665]), .B2(n2784), 
        .ZN(n14906) );
  MOAI22 U23820 ( .A1(n28720), .A2(n2783), .B1(ram[10666]), .B2(n2784), 
        .ZN(n14907) );
  MOAI22 U23821 ( .A1(n28485), .A2(n2783), .B1(ram[10667]), .B2(n2784), 
        .ZN(n14908) );
  MOAI22 U23822 ( .A1(n28250), .A2(n2783), .B1(ram[10668]), .B2(n2784), 
        .ZN(n14909) );
  MOAI22 U23823 ( .A1(n28015), .A2(n2783), .B1(ram[10669]), .B2(n2784), 
        .ZN(n14910) );
  MOAI22 U23824 ( .A1(n27780), .A2(n2783), .B1(ram[10670]), .B2(n2784), 
        .ZN(n14911) );
  MOAI22 U23825 ( .A1(n27545), .A2(n2783), .B1(ram[10671]), .B2(n2784), 
        .ZN(n14912) );
  MOAI22 U23826 ( .A1(n29190), .A2(n2785), .B1(ram[10672]), .B2(n2786), 
        .ZN(n14913) );
  MOAI22 U23827 ( .A1(n28955), .A2(n2785), .B1(ram[10673]), .B2(n2786), 
        .ZN(n14914) );
  MOAI22 U23828 ( .A1(n28720), .A2(n2785), .B1(ram[10674]), .B2(n2786), 
        .ZN(n14915) );
  MOAI22 U23829 ( .A1(n28485), .A2(n2785), .B1(ram[10675]), .B2(n2786), 
        .ZN(n14916) );
  MOAI22 U23830 ( .A1(n28250), .A2(n2785), .B1(ram[10676]), .B2(n2786), 
        .ZN(n14917) );
  MOAI22 U23831 ( .A1(n28015), .A2(n2785), .B1(ram[10677]), .B2(n2786), 
        .ZN(n14918) );
  MOAI22 U23832 ( .A1(n27780), .A2(n2785), .B1(ram[10678]), .B2(n2786), 
        .ZN(n14919) );
  MOAI22 U23833 ( .A1(n27545), .A2(n2785), .B1(ram[10679]), .B2(n2786), 
        .ZN(n14920) );
  MOAI22 U23834 ( .A1(n29190), .A2(n2787), .B1(ram[10680]), .B2(n2788), 
        .ZN(n14921) );
  MOAI22 U23835 ( .A1(n28955), .A2(n2787), .B1(ram[10681]), .B2(n2788), 
        .ZN(n14922) );
  MOAI22 U23836 ( .A1(n28720), .A2(n2787), .B1(ram[10682]), .B2(n2788), 
        .ZN(n14923) );
  MOAI22 U23837 ( .A1(n28485), .A2(n2787), .B1(ram[10683]), .B2(n2788), 
        .ZN(n14924) );
  MOAI22 U23838 ( .A1(n28250), .A2(n2787), .B1(ram[10684]), .B2(n2788), 
        .ZN(n14925) );
  MOAI22 U23839 ( .A1(n28015), .A2(n2787), .B1(ram[10685]), .B2(n2788), 
        .ZN(n14926) );
  MOAI22 U23840 ( .A1(n27780), .A2(n2787), .B1(ram[10686]), .B2(n2788), 
        .ZN(n14927) );
  MOAI22 U23841 ( .A1(n27545), .A2(n2787), .B1(ram[10687]), .B2(n2788), 
        .ZN(n14928) );
  MOAI22 U23842 ( .A1(n29190), .A2(n2789), .B1(ram[10688]), .B2(n2790), 
        .ZN(n14929) );
  MOAI22 U23843 ( .A1(n28955), .A2(n2789), .B1(ram[10689]), .B2(n2790), 
        .ZN(n14930) );
  MOAI22 U23844 ( .A1(n28720), .A2(n2789), .B1(ram[10690]), .B2(n2790), 
        .ZN(n14931) );
  MOAI22 U23845 ( .A1(n28485), .A2(n2789), .B1(ram[10691]), .B2(n2790), 
        .ZN(n14932) );
  MOAI22 U23846 ( .A1(n28250), .A2(n2789), .B1(ram[10692]), .B2(n2790), 
        .ZN(n14933) );
  MOAI22 U23847 ( .A1(n28015), .A2(n2789), .B1(ram[10693]), .B2(n2790), 
        .ZN(n14934) );
  MOAI22 U23848 ( .A1(n27780), .A2(n2789), .B1(ram[10694]), .B2(n2790), 
        .ZN(n14935) );
  MOAI22 U23849 ( .A1(n27545), .A2(n2789), .B1(ram[10695]), .B2(n2790), 
        .ZN(n14936) );
  MOAI22 U23850 ( .A1(n29190), .A2(n2791), .B1(ram[10696]), .B2(n2792), 
        .ZN(n14937) );
  MOAI22 U23851 ( .A1(n28955), .A2(n2791), .B1(ram[10697]), .B2(n2792), 
        .ZN(n14938) );
  MOAI22 U23852 ( .A1(n28720), .A2(n2791), .B1(ram[10698]), .B2(n2792), 
        .ZN(n14939) );
  MOAI22 U23853 ( .A1(n28485), .A2(n2791), .B1(ram[10699]), .B2(n2792), 
        .ZN(n14940) );
  MOAI22 U23854 ( .A1(n28250), .A2(n2791), .B1(ram[10700]), .B2(n2792), 
        .ZN(n14941) );
  MOAI22 U23855 ( .A1(n28015), .A2(n2791), .B1(ram[10701]), .B2(n2792), 
        .ZN(n14942) );
  MOAI22 U23856 ( .A1(n27780), .A2(n2791), .B1(ram[10702]), .B2(n2792), 
        .ZN(n14943) );
  MOAI22 U23857 ( .A1(n27545), .A2(n2791), .B1(ram[10703]), .B2(n2792), 
        .ZN(n14944) );
  MOAI22 U23858 ( .A1(n29190), .A2(n2793), .B1(ram[10704]), .B2(n2794), 
        .ZN(n14945) );
  MOAI22 U23859 ( .A1(n28955), .A2(n2793), .B1(ram[10705]), .B2(n2794), 
        .ZN(n14946) );
  MOAI22 U23860 ( .A1(n28720), .A2(n2793), .B1(ram[10706]), .B2(n2794), 
        .ZN(n14947) );
  MOAI22 U23861 ( .A1(n28485), .A2(n2793), .B1(ram[10707]), .B2(n2794), 
        .ZN(n14948) );
  MOAI22 U23862 ( .A1(n28250), .A2(n2793), .B1(ram[10708]), .B2(n2794), 
        .ZN(n14949) );
  MOAI22 U23863 ( .A1(n28015), .A2(n2793), .B1(ram[10709]), .B2(n2794), 
        .ZN(n14950) );
  MOAI22 U23864 ( .A1(n27780), .A2(n2793), .B1(ram[10710]), .B2(n2794), 
        .ZN(n14951) );
  MOAI22 U23865 ( .A1(n27545), .A2(n2793), .B1(ram[10711]), .B2(n2794), 
        .ZN(n14952) );
  MOAI22 U23866 ( .A1(n29191), .A2(n2795), .B1(ram[10712]), .B2(n2796), 
        .ZN(n14953) );
  MOAI22 U23867 ( .A1(n28956), .A2(n2795), .B1(ram[10713]), .B2(n2796), 
        .ZN(n14954) );
  MOAI22 U23868 ( .A1(n28721), .A2(n2795), .B1(ram[10714]), .B2(n2796), 
        .ZN(n14955) );
  MOAI22 U23869 ( .A1(n28486), .A2(n2795), .B1(ram[10715]), .B2(n2796), 
        .ZN(n14956) );
  MOAI22 U23870 ( .A1(n28251), .A2(n2795), .B1(ram[10716]), .B2(n2796), 
        .ZN(n14957) );
  MOAI22 U23871 ( .A1(n28016), .A2(n2795), .B1(ram[10717]), .B2(n2796), 
        .ZN(n14958) );
  MOAI22 U23872 ( .A1(n27781), .A2(n2795), .B1(ram[10718]), .B2(n2796), 
        .ZN(n14959) );
  MOAI22 U23873 ( .A1(n27546), .A2(n2795), .B1(ram[10719]), .B2(n2796), 
        .ZN(n14960) );
  MOAI22 U23874 ( .A1(n29191), .A2(n2797), .B1(ram[10720]), .B2(n2798), 
        .ZN(n14961) );
  MOAI22 U23875 ( .A1(n28956), .A2(n2797), .B1(ram[10721]), .B2(n2798), 
        .ZN(n14962) );
  MOAI22 U23876 ( .A1(n28721), .A2(n2797), .B1(ram[10722]), .B2(n2798), 
        .ZN(n14963) );
  MOAI22 U23877 ( .A1(n28486), .A2(n2797), .B1(ram[10723]), .B2(n2798), 
        .ZN(n14964) );
  MOAI22 U23878 ( .A1(n28251), .A2(n2797), .B1(ram[10724]), .B2(n2798), 
        .ZN(n14965) );
  MOAI22 U23879 ( .A1(n28016), .A2(n2797), .B1(ram[10725]), .B2(n2798), 
        .ZN(n14966) );
  MOAI22 U23880 ( .A1(n27781), .A2(n2797), .B1(ram[10726]), .B2(n2798), 
        .ZN(n14967) );
  MOAI22 U23881 ( .A1(n27546), .A2(n2797), .B1(ram[10727]), .B2(n2798), 
        .ZN(n14968) );
  MOAI22 U23882 ( .A1(n29191), .A2(n2799), .B1(ram[10728]), .B2(n2800), 
        .ZN(n14969) );
  MOAI22 U23883 ( .A1(n28956), .A2(n2799), .B1(ram[10729]), .B2(n2800), 
        .ZN(n14970) );
  MOAI22 U23884 ( .A1(n28721), .A2(n2799), .B1(ram[10730]), .B2(n2800), 
        .ZN(n14971) );
  MOAI22 U23885 ( .A1(n28486), .A2(n2799), .B1(ram[10731]), .B2(n2800), 
        .ZN(n14972) );
  MOAI22 U23886 ( .A1(n28251), .A2(n2799), .B1(ram[10732]), .B2(n2800), 
        .ZN(n14973) );
  MOAI22 U23887 ( .A1(n28016), .A2(n2799), .B1(ram[10733]), .B2(n2800), 
        .ZN(n14974) );
  MOAI22 U23888 ( .A1(n27781), .A2(n2799), .B1(ram[10734]), .B2(n2800), 
        .ZN(n14975) );
  MOAI22 U23889 ( .A1(n27546), .A2(n2799), .B1(ram[10735]), .B2(n2800), 
        .ZN(n14976) );
  MOAI22 U23890 ( .A1(n29191), .A2(n2801), .B1(ram[10736]), .B2(n2802), 
        .ZN(n14977) );
  MOAI22 U23891 ( .A1(n28956), .A2(n2801), .B1(ram[10737]), .B2(n2802), 
        .ZN(n14978) );
  MOAI22 U23892 ( .A1(n28721), .A2(n2801), .B1(ram[10738]), .B2(n2802), 
        .ZN(n14979) );
  MOAI22 U23893 ( .A1(n28486), .A2(n2801), .B1(ram[10739]), .B2(n2802), 
        .ZN(n14980) );
  MOAI22 U23894 ( .A1(n28251), .A2(n2801), .B1(ram[10740]), .B2(n2802), 
        .ZN(n14981) );
  MOAI22 U23895 ( .A1(n28016), .A2(n2801), .B1(ram[10741]), .B2(n2802), 
        .ZN(n14982) );
  MOAI22 U23896 ( .A1(n27781), .A2(n2801), .B1(ram[10742]), .B2(n2802), 
        .ZN(n14983) );
  MOAI22 U23897 ( .A1(n27546), .A2(n2801), .B1(ram[10743]), .B2(n2802), 
        .ZN(n14984) );
  MOAI22 U23898 ( .A1(n29191), .A2(n2803), .B1(ram[10744]), .B2(n2804), 
        .ZN(n14985) );
  MOAI22 U23899 ( .A1(n28956), .A2(n2803), .B1(ram[10745]), .B2(n2804), 
        .ZN(n14986) );
  MOAI22 U23900 ( .A1(n28721), .A2(n2803), .B1(ram[10746]), .B2(n2804), 
        .ZN(n14987) );
  MOAI22 U23901 ( .A1(n28486), .A2(n2803), .B1(ram[10747]), .B2(n2804), 
        .ZN(n14988) );
  MOAI22 U23902 ( .A1(n28251), .A2(n2803), .B1(ram[10748]), .B2(n2804), 
        .ZN(n14989) );
  MOAI22 U23903 ( .A1(n28016), .A2(n2803), .B1(ram[10749]), .B2(n2804), 
        .ZN(n14990) );
  MOAI22 U23904 ( .A1(n27781), .A2(n2803), .B1(ram[10750]), .B2(n2804), 
        .ZN(n14991) );
  MOAI22 U23905 ( .A1(n27546), .A2(n2803), .B1(ram[10751]), .B2(n2804), 
        .ZN(n14992) );
  MOAI22 U23906 ( .A1(n29191), .A2(n2805), .B1(ram[10752]), .B2(n2806), 
        .ZN(n14993) );
  MOAI22 U23907 ( .A1(n28956), .A2(n2805), .B1(ram[10753]), .B2(n2806), 
        .ZN(n14994) );
  MOAI22 U23908 ( .A1(n28721), .A2(n2805), .B1(ram[10754]), .B2(n2806), 
        .ZN(n14995) );
  MOAI22 U23909 ( .A1(n28486), .A2(n2805), .B1(ram[10755]), .B2(n2806), 
        .ZN(n14996) );
  MOAI22 U23910 ( .A1(n28251), .A2(n2805), .B1(ram[10756]), .B2(n2806), 
        .ZN(n14997) );
  MOAI22 U23911 ( .A1(n28016), .A2(n2805), .B1(ram[10757]), .B2(n2806), 
        .ZN(n14998) );
  MOAI22 U23912 ( .A1(n27781), .A2(n2805), .B1(ram[10758]), .B2(n2806), 
        .ZN(n14999) );
  MOAI22 U23913 ( .A1(n27546), .A2(n2805), .B1(ram[10759]), .B2(n2806), 
        .ZN(n15000) );
  MOAI22 U23914 ( .A1(n29191), .A2(n2808), .B1(ram[10760]), .B2(n2809), 
        .ZN(n15001) );
  MOAI22 U23915 ( .A1(n28956), .A2(n2808), .B1(ram[10761]), .B2(n2809), 
        .ZN(n15002) );
  MOAI22 U23916 ( .A1(n28721), .A2(n2808), .B1(ram[10762]), .B2(n2809), 
        .ZN(n15003) );
  MOAI22 U23917 ( .A1(n28486), .A2(n2808), .B1(ram[10763]), .B2(n2809), 
        .ZN(n15004) );
  MOAI22 U23918 ( .A1(n28251), .A2(n2808), .B1(ram[10764]), .B2(n2809), 
        .ZN(n15005) );
  MOAI22 U23919 ( .A1(n28016), .A2(n2808), .B1(ram[10765]), .B2(n2809), 
        .ZN(n15006) );
  MOAI22 U23920 ( .A1(n27781), .A2(n2808), .B1(ram[10766]), .B2(n2809), 
        .ZN(n15007) );
  MOAI22 U23921 ( .A1(n27546), .A2(n2808), .B1(ram[10767]), .B2(n2809), 
        .ZN(n15008) );
  MOAI22 U23922 ( .A1(n29191), .A2(n2810), .B1(ram[10768]), .B2(n2811), 
        .ZN(n15009) );
  MOAI22 U23923 ( .A1(n28956), .A2(n2810), .B1(ram[10769]), .B2(n2811), 
        .ZN(n15010) );
  MOAI22 U23924 ( .A1(n28721), .A2(n2810), .B1(ram[10770]), .B2(n2811), 
        .ZN(n15011) );
  MOAI22 U23925 ( .A1(n28486), .A2(n2810), .B1(ram[10771]), .B2(n2811), 
        .ZN(n15012) );
  MOAI22 U23926 ( .A1(n28251), .A2(n2810), .B1(ram[10772]), .B2(n2811), 
        .ZN(n15013) );
  MOAI22 U23927 ( .A1(n28016), .A2(n2810), .B1(ram[10773]), .B2(n2811), 
        .ZN(n15014) );
  MOAI22 U23928 ( .A1(n27781), .A2(n2810), .B1(ram[10774]), .B2(n2811), 
        .ZN(n15015) );
  MOAI22 U23929 ( .A1(n27546), .A2(n2810), .B1(ram[10775]), .B2(n2811), 
        .ZN(n15016) );
  MOAI22 U23930 ( .A1(n29191), .A2(n2812), .B1(ram[10776]), .B2(n2813), 
        .ZN(n15017) );
  MOAI22 U23931 ( .A1(n28956), .A2(n2812), .B1(ram[10777]), .B2(n2813), 
        .ZN(n15018) );
  MOAI22 U23932 ( .A1(n28721), .A2(n2812), .B1(ram[10778]), .B2(n2813), 
        .ZN(n15019) );
  MOAI22 U23933 ( .A1(n28486), .A2(n2812), .B1(ram[10779]), .B2(n2813), 
        .ZN(n15020) );
  MOAI22 U23934 ( .A1(n28251), .A2(n2812), .B1(ram[10780]), .B2(n2813), 
        .ZN(n15021) );
  MOAI22 U23935 ( .A1(n28016), .A2(n2812), .B1(ram[10781]), .B2(n2813), 
        .ZN(n15022) );
  MOAI22 U23936 ( .A1(n27781), .A2(n2812), .B1(ram[10782]), .B2(n2813), 
        .ZN(n15023) );
  MOAI22 U23937 ( .A1(n27546), .A2(n2812), .B1(ram[10783]), .B2(n2813), 
        .ZN(n15024) );
  MOAI22 U23938 ( .A1(n29191), .A2(n2814), .B1(ram[10784]), .B2(n2815), 
        .ZN(n15025) );
  MOAI22 U23939 ( .A1(n28956), .A2(n2814), .B1(ram[10785]), .B2(n2815), 
        .ZN(n15026) );
  MOAI22 U23940 ( .A1(n28721), .A2(n2814), .B1(ram[10786]), .B2(n2815), 
        .ZN(n15027) );
  MOAI22 U23941 ( .A1(n28486), .A2(n2814), .B1(ram[10787]), .B2(n2815), 
        .ZN(n15028) );
  MOAI22 U23942 ( .A1(n28251), .A2(n2814), .B1(ram[10788]), .B2(n2815), 
        .ZN(n15029) );
  MOAI22 U23943 ( .A1(n28016), .A2(n2814), .B1(ram[10789]), .B2(n2815), 
        .ZN(n15030) );
  MOAI22 U23944 ( .A1(n27781), .A2(n2814), .B1(ram[10790]), .B2(n2815), 
        .ZN(n15031) );
  MOAI22 U23945 ( .A1(n27546), .A2(n2814), .B1(ram[10791]), .B2(n2815), 
        .ZN(n15032) );
  MOAI22 U23946 ( .A1(n29191), .A2(n2816), .B1(ram[10792]), .B2(n2817), 
        .ZN(n15033) );
  MOAI22 U23947 ( .A1(n28956), .A2(n2816), .B1(ram[10793]), .B2(n2817), 
        .ZN(n15034) );
  MOAI22 U23948 ( .A1(n28721), .A2(n2816), .B1(ram[10794]), .B2(n2817), 
        .ZN(n15035) );
  MOAI22 U23949 ( .A1(n28486), .A2(n2816), .B1(ram[10795]), .B2(n2817), 
        .ZN(n15036) );
  MOAI22 U23950 ( .A1(n28251), .A2(n2816), .B1(ram[10796]), .B2(n2817), 
        .ZN(n15037) );
  MOAI22 U23951 ( .A1(n28016), .A2(n2816), .B1(ram[10797]), .B2(n2817), 
        .ZN(n15038) );
  MOAI22 U23952 ( .A1(n27781), .A2(n2816), .B1(ram[10798]), .B2(n2817), 
        .ZN(n15039) );
  MOAI22 U23953 ( .A1(n27546), .A2(n2816), .B1(ram[10799]), .B2(n2817), 
        .ZN(n15040) );
  MOAI22 U23954 ( .A1(n29191), .A2(n2818), .B1(ram[10800]), .B2(n2819), 
        .ZN(n15041) );
  MOAI22 U23955 ( .A1(n28956), .A2(n2818), .B1(ram[10801]), .B2(n2819), 
        .ZN(n15042) );
  MOAI22 U23956 ( .A1(n28721), .A2(n2818), .B1(ram[10802]), .B2(n2819), 
        .ZN(n15043) );
  MOAI22 U23957 ( .A1(n28486), .A2(n2818), .B1(ram[10803]), .B2(n2819), 
        .ZN(n15044) );
  MOAI22 U23958 ( .A1(n28251), .A2(n2818), .B1(ram[10804]), .B2(n2819), 
        .ZN(n15045) );
  MOAI22 U23959 ( .A1(n28016), .A2(n2818), .B1(ram[10805]), .B2(n2819), 
        .ZN(n15046) );
  MOAI22 U23960 ( .A1(n27781), .A2(n2818), .B1(ram[10806]), .B2(n2819), 
        .ZN(n15047) );
  MOAI22 U23961 ( .A1(n27546), .A2(n2818), .B1(ram[10807]), .B2(n2819), 
        .ZN(n15048) );
  MOAI22 U23962 ( .A1(n29191), .A2(n2820), .B1(ram[10808]), .B2(n2821), 
        .ZN(n15049) );
  MOAI22 U23963 ( .A1(n28956), .A2(n2820), .B1(ram[10809]), .B2(n2821), 
        .ZN(n15050) );
  MOAI22 U23964 ( .A1(n28721), .A2(n2820), .B1(ram[10810]), .B2(n2821), 
        .ZN(n15051) );
  MOAI22 U23965 ( .A1(n28486), .A2(n2820), .B1(ram[10811]), .B2(n2821), 
        .ZN(n15052) );
  MOAI22 U23966 ( .A1(n28251), .A2(n2820), .B1(ram[10812]), .B2(n2821), 
        .ZN(n15053) );
  MOAI22 U23967 ( .A1(n28016), .A2(n2820), .B1(ram[10813]), .B2(n2821), 
        .ZN(n15054) );
  MOAI22 U23968 ( .A1(n27781), .A2(n2820), .B1(ram[10814]), .B2(n2821), 
        .ZN(n15055) );
  MOAI22 U23969 ( .A1(n27546), .A2(n2820), .B1(ram[10815]), .B2(n2821), 
        .ZN(n15056) );
  MOAI22 U23970 ( .A1(n29192), .A2(n2822), .B1(ram[10816]), .B2(n2823), 
        .ZN(n15057) );
  MOAI22 U23971 ( .A1(n28957), .A2(n2822), .B1(ram[10817]), .B2(n2823), 
        .ZN(n15058) );
  MOAI22 U23972 ( .A1(n28722), .A2(n2822), .B1(ram[10818]), .B2(n2823), 
        .ZN(n15059) );
  MOAI22 U23973 ( .A1(n28487), .A2(n2822), .B1(ram[10819]), .B2(n2823), 
        .ZN(n15060) );
  MOAI22 U23974 ( .A1(n28252), .A2(n2822), .B1(ram[10820]), .B2(n2823), 
        .ZN(n15061) );
  MOAI22 U23975 ( .A1(n28017), .A2(n2822), .B1(ram[10821]), .B2(n2823), 
        .ZN(n15062) );
  MOAI22 U23976 ( .A1(n27782), .A2(n2822), .B1(ram[10822]), .B2(n2823), 
        .ZN(n15063) );
  MOAI22 U23977 ( .A1(n27547), .A2(n2822), .B1(ram[10823]), .B2(n2823), 
        .ZN(n15064) );
  MOAI22 U23978 ( .A1(n29192), .A2(n2824), .B1(ram[10824]), .B2(n2825), 
        .ZN(n15065) );
  MOAI22 U23979 ( .A1(n28957), .A2(n2824), .B1(ram[10825]), .B2(n2825), 
        .ZN(n15066) );
  MOAI22 U23980 ( .A1(n28722), .A2(n2824), .B1(ram[10826]), .B2(n2825), 
        .ZN(n15067) );
  MOAI22 U23981 ( .A1(n28487), .A2(n2824), .B1(ram[10827]), .B2(n2825), 
        .ZN(n15068) );
  MOAI22 U23982 ( .A1(n28252), .A2(n2824), .B1(ram[10828]), .B2(n2825), 
        .ZN(n15069) );
  MOAI22 U23983 ( .A1(n28017), .A2(n2824), .B1(ram[10829]), .B2(n2825), 
        .ZN(n15070) );
  MOAI22 U23984 ( .A1(n27782), .A2(n2824), .B1(ram[10830]), .B2(n2825), 
        .ZN(n15071) );
  MOAI22 U23985 ( .A1(n27547), .A2(n2824), .B1(ram[10831]), .B2(n2825), 
        .ZN(n15072) );
  MOAI22 U23986 ( .A1(n29192), .A2(n2826), .B1(ram[10832]), .B2(n2827), 
        .ZN(n15073) );
  MOAI22 U23987 ( .A1(n28957), .A2(n2826), .B1(ram[10833]), .B2(n2827), 
        .ZN(n15074) );
  MOAI22 U23988 ( .A1(n28722), .A2(n2826), .B1(ram[10834]), .B2(n2827), 
        .ZN(n15075) );
  MOAI22 U23989 ( .A1(n28487), .A2(n2826), .B1(ram[10835]), .B2(n2827), 
        .ZN(n15076) );
  MOAI22 U23990 ( .A1(n28252), .A2(n2826), .B1(ram[10836]), .B2(n2827), 
        .ZN(n15077) );
  MOAI22 U23991 ( .A1(n28017), .A2(n2826), .B1(ram[10837]), .B2(n2827), 
        .ZN(n15078) );
  MOAI22 U23992 ( .A1(n27782), .A2(n2826), .B1(ram[10838]), .B2(n2827), 
        .ZN(n15079) );
  MOAI22 U23993 ( .A1(n27547), .A2(n2826), .B1(ram[10839]), .B2(n2827), 
        .ZN(n15080) );
  MOAI22 U23994 ( .A1(n29192), .A2(n2828), .B1(ram[10840]), .B2(n2829), 
        .ZN(n15081) );
  MOAI22 U23995 ( .A1(n28957), .A2(n2828), .B1(ram[10841]), .B2(n2829), 
        .ZN(n15082) );
  MOAI22 U23996 ( .A1(n28722), .A2(n2828), .B1(ram[10842]), .B2(n2829), 
        .ZN(n15083) );
  MOAI22 U23997 ( .A1(n28487), .A2(n2828), .B1(ram[10843]), .B2(n2829), 
        .ZN(n15084) );
  MOAI22 U23998 ( .A1(n28252), .A2(n2828), .B1(ram[10844]), .B2(n2829), 
        .ZN(n15085) );
  MOAI22 U23999 ( .A1(n28017), .A2(n2828), .B1(ram[10845]), .B2(n2829), 
        .ZN(n15086) );
  MOAI22 U24000 ( .A1(n27782), .A2(n2828), .B1(ram[10846]), .B2(n2829), 
        .ZN(n15087) );
  MOAI22 U24001 ( .A1(n27547), .A2(n2828), .B1(ram[10847]), .B2(n2829), 
        .ZN(n15088) );
  MOAI22 U24002 ( .A1(n29192), .A2(n2830), .B1(ram[10848]), .B2(n2831), 
        .ZN(n15089) );
  MOAI22 U24003 ( .A1(n28957), .A2(n2830), .B1(ram[10849]), .B2(n2831), 
        .ZN(n15090) );
  MOAI22 U24004 ( .A1(n28722), .A2(n2830), .B1(ram[10850]), .B2(n2831), 
        .ZN(n15091) );
  MOAI22 U24005 ( .A1(n28487), .A2(n2830), .B1(ram[10851]), .B2(n2831), 
        .ZN(n15092) );
  MOAI22 U24006 ( .A1(n28252), .A2(n2830), .B1(ram[10852]), .B2(n2831), 
        .ZN(n15093) );
  MOAI22 U24007 ( .A1(n28017), .A2(n2830), .B1(ram[10853]), .B2(n2831), 
        .ZN(n15094) );
  MOAI22 U24008 ( .A1(n27782), .A2(n2830), .B1(ram[10854]), .B2(n2831), 
        .ZN(n15095) );
  MOAI22 U24009 ( .A1(n27547), .A2(n2830), .B1(ram[10855]), .B2(n2831), 
        .ZN(n15096) );
  MOAI22 U24010 ( .A1(n29192), .A2(n2832), .B1(ram[10856]), .B2(n2833), 
        .ZN(n15097) );
  MOAI22 U24011 ( .A1(n28957), .A2(n2832), .B1(ram[10857]), .B2(n2833), 
        .ZN(n15098) );
  MOAI22 U24012 ( .A1(n28722), .A2(n2832), .B1(ram[10858]), .B2(n2833), 
        .ZN(n15099) );
  MOAI22 U24013 ( .A1(n28487), .A2(n2832), .B1(ram[10859]), .B2(n2833), 
        .ZN(n15100) );
  MOAI22 U24014 ( .A1(n28252), .A2(n2832), .B1(ram[10860]), .B2(n2833), 
        .ZN(n15101) );
  MOAI22 U24015 ( .A1(n28017), .A2(n2832), .B1(ram[10861]), .B2(n2833), 
        .ZN(n15102) );
  MOAI22 U24016 ( .A1(n27782), .A2(n2832), .B1(ram[10862]), .B2(n2833), 
        .ZN(n15103) );
  MOAI22 U24017 ( .A1(n27547), .A2(n2832), .B1(ram[10863]), .B2(n2833), 
        .ZN(n15104) );
  MOAI22 U24018 ( .A1(n29192), .A2(n2834), .B1(ram[10864]), .B2(n2835), 
        .ZN(n15105) );
  MOAI22 U24019 ( .A1(n28957), .A2(n2834), .B1(ram[10865]), .B2(n2835), 
        .ZN(n15106) );
  MOAI22 U24020 ( .A1(n28722), .A2(n2834), .B1(ram[10866]), .B2(n2835), 
        .ZN(n15107) );
  MOAI22 U24021 ( .A1(n28487), .A2(n2834), .B1(ram[10867]), .B2(n2835), 
        .ZN(n15108) );
  MOAI22 U24022 ( .A1(n28252), .A2(n2834), .B1(ram[10868]), .B2(n2835), 
        .ZN(n15109) );
  MOAI22 U24023 ( .A1(n28017), .A2(n2834), .B1(ram[10869]), .B2(n2835), 
        .ZN(n15110) );
  MOAI22 U24024 ( .A1(n27782), .A2(n2834), .B1(ram[10870]), .B2(n2835), 
        .ZN(n15111) );
  MOAI22 U24025 ( .A1(n27547), .A2(n2834), .B1(ram[10871]), .B2(n2835), 
        .ZN(n15112) );
  MOAI22 U24026 ( .A1(n29192), .A2(n2836), .B1(ram[10872]), .B2(n2837), 
        .ZN(n15113) );
  MOAI22 U24027 ( .A1(n28957), .A2(n2836), .B1(ram[10873]), .B2(n2837), 
        .ZN(n15114) );
  MOAI22 U24028 ( .A1(n28722), .A2(n2836), .B1(ram[10874]), .B2(n2837), 
        .ZN(n15115) );
  MOAI22 U24029 ( .A1(n28487), .A2(n2836), .B1(ram[10875]), .B2(n2837), 
        .ZN(n15116) );
  MOAI22 U24030 ( .A1(n28252), .A2(n2836), .B1(ram[10876]), .B2(n2837), 
        .ZN(n15117) );
  MOAI22 U24031 ( .A1(n28017), .A2(n2836), .B1(ram[10877]), .B2(n2837), 
        .ZN(n15118) );
  MOAI22 U24032 ( .A1(n27782), .A2(n2836), .B1(ram[10878]), .B2(n2837), 
        .ZN(n15119) );
  MOAI22 U24033 ( .A1(n27547), .A2(n2836), .B1(ram[10879]), .B2(n2837), 
        .ZN(n15120) );
  MOAI22 U24034 ( .A1(n29192), .A2(n2838), .B1(ram[10880]), .B2(n2839), 
        .ZN(n15121) );
  MOAI22 U24035 ( .A1(n28957), .A2(n2838), .B1(ram[10881]), .B2(n2839), 
        .ZN(n15122) );
  MOAI22 U24036 ( .A1(n28722), .A2(n2838), .B1(ram[10882]), .B2(n2839), 
        .ZN(n15123) );
  MOAI22 U24037 ( .A1(n28487), .A2(n2838), .B1(ram[10883]), .B2(n2839), 
        .ZN(n15124) );
  MOAI22 U24038 ( .A1(n28252), .A2(n2838), .B1(ram[10884]), .B2(n2839), 
        .ZN(n15125) );
  MOAI22 U24039 ( .A1(n28017), .A2(n2838), .B1(ram[10885]), .B2(n2839), 
        .ZN(n15126) );
  MOAI22 U24040 ( .A1(n27782), .A2(n2838), .B1(ram[10886]), .B2(n2839), 
        .ZN(n15127) );
  MOAI22 U24041 ( .A1(n27547), .A2(n2838), .B1(ram[10887]), .B2(n2839), 
        .ZN(n15128) );
  MOAI22 U24042 ( .A1(n29192), .A2(n2840), .B1(ram[10888]), .B2(n2841), 
        .ZN(n15129) );
  MOAI22 U24043 ( .A1(n28957), .A2(n2840), .B1(ram[10889]), .B2(n2841), 
        .ZN(n15130) );
  MOAI22 U24044 ( .A1(n28722), .A2(n2840), .B1(ram[10890]), .B2(n2841), 
        .ZN(n15131) );
  MOAI22 U24045 ( .A1(n28487), .A2(n2840), .B1(ram[10891]), .B2(n2841), 
        .ZN(n15132) );
  MOAI22 U24046 ( .A1(n28252), .A2(n2840), .B1(ram[10892]), .B2(n2841), 
        .ZN(n15133) );
  MOAI22 U24047 ( .A1(n28017), .A2(n2840), .B1(ram[10893]), .B2(n2841), 
        .ZN(n15134) );
  MOAI22 U24048 ( .A1(n27782), .A2(n2840), .B1(ram[10894]), .B2(n2841), 
        .ZN(n15135) );
  MOAI22 U24049 ( .A1(n27547), .A2(n2840), .B1(ram[10895]), .B2(n2841), 
        .ZN(n15136) );
  MOAI22 U24050 ( .A1(n29192), .A2(n2842), .B1(ram[10896]), .B2(n2843), 
        .ZN(n15137) );
  MOAI22 U24051 ( .A1(n28957), .A2(n2842), .B1(ram[10897]), .B2(n2843), 
        .ZN(n15138) );
  MOAI22 U24052 ( .A1(n28722), .A2(n2842), .B1(ram[10898]), .B2(n2843), 
        .ZN(n15139) );
  MOAI22 U24053 ( .A1(n28487), .A2(n2842), .B1(ram[10899]), .B2(n2843), 
        .ZN(n15140) );
  MOAI22 U24054 ( .A1(n28252), .A2(n2842), .B1(ram[10900]), .B2(n2843), 
        .ZN(n15141) );
  MOAI22 U24055 ( .A1(n28017), .A2(n2842), .B1(ram[10901]), .B2(n2843), 
        .ZN(n15142) );
  MOAI22 U24056 ( .A1(n27782), .A2(n2842), .B1(ram[10902]), .B2(n2843), 
        .ZN(n15143) );
  MOAI22 U24057 ( .A1(n27547), .A2(n2842), .B1(ram[10903]), .B2(n2843), 
        .ZN(n15144) );
  MOAI22 U24058 ( .A1(n29192), .A2(n2844), .B1(ram[10904]), .B2(n2845), 
        .ZN(n15145) );
  MOAI22 U24059 ( .A1(n28957), .A2(n2844), .B1(ram[10905]), .B2(n2845), 
        .ZN(n15146) );
  MOAI22 U24060 ( .A1(n28722), .A2(n2844), .B1(ram[10906]), .B2(n2845), 
        .ZN(n15147) );
  MOAI22 U24061 ( .A1(n28487), .A2(n2844), .B1(ram[10907]), .B2(n2845), 
        .ZN(n15148) );
  MOAI22 U24062 ( .A1(n28252), .A2(n2844), .B1(ram[10908]), .B2(n2845), 
        .ZN(n15149) );
  MOAI22 U24063 ( .A1(n28017), .A2(n2844), .B1(ram[10909]), .B2(n2845), 
        .ZN(n15150) );
  MOAI22 U24064 ( .A1(n27782), .A2(n2844), .B1(ram[10910]), .B2(n2845), 
        .ZN(n15151) );
  MOAI22 U24065 ( .A1(n27547), .A2(n2844), .B1(ram[10911]), .B2(n2845), 
        .ZN(n15152) );
  MOAI22 U24066 ( .A1(n29192), .A2(n2846), .B1(ram[10912]), .B2(n2847), 
        .ZN(n15153) );
  MOAI22 U24067 ( .A1(n28957), .A2(n2846), .B1(ram[10913]), .B2(n2847), 
        .ZN(n15154) );
  MOAI22 U24068 ( .A1(n28722), .A2(n2846), .B1(ram[10914]), .B2(n2847), 
        .ZN(n15155) );
  MOAI22 U24069 ( .A1(n28487), .A2(n2846), .B1(ram[10915]), .B2(n2847), 
        .ZN(n15156) );
  MOAI22 U24070 ( .A1(n28252), .A2(n2846), .B1(ram[10916]), .B2(n2847), 
        .ZN(n15157) );
  MOAI22 U24071 ( .A1(n28017), .A2(n2846), .B1(ram[10917]), .B2(n2847), 
        .ZN(n15158) );
  MOAI22 U24072 ( .A1(n27782), .A2(n2846), .B1(ram[10918]), .B2(n2847), 
        .ZN(n15159) );
  MOAI22 U24073 ( .A1(n27547), .A2(n2846), .B1(ram[10919]), .B2(n2847), 
        .ZN(n15160) );
  MOAI22 U24074 ( .A1(n29193), .A2(n2848), .B1(ram[10920]), .B2(n2849), 
        .ZN(n15161) );
  MOAI22 U24075 ( .A1(n28958), .A2(n2848), .B1(ram[10921]), .B2(n2849), 
        .ZN(n15162) );
  MOAI22 U24076 ( .A1(n28723), .A2(n2848), .B1(ram[10922]), .B2(n2849), 
        .ZN(n15163) );
  MOAI22 U24077 ( .A1(n28488), .A2(n2848), .B1(ram[10923]), .B2(n2849), 
        .ZN(n15164) );
  MOAI22 U24078 ( .A1(n28253), .A2(n2848), .B1(ram[10924]), .B2(n2849), 
        .ZN(n15165) );
  MOAI22 U24079 ( .A1(n28018), .A2(n2848), .B1(ram[10925]), .B2(n2849), 
        .ZN(n15166) );
  MOAI22 U24080 ( .A1(n27783), .A2(n2848), .B1(ram[10926]), .B2(n2849), 
        .ZN(n15167) );
  MOAI22 U24081 ( .A1(n27548), .A2(n2848), .B1(ram[10927]), .B2(n2849), 
        .ZN(n15168) );
  MOAI22 U24082 ( .A1(n29193), .A2(n2850), .B1(ram[10928]), .B2(n2851), 
        .ZN(n15169) );
  MOAI22 U24083 ( .A1(n28958), .A2(n2850), .B1(ram[10929]), .B2(n2851), 
        .ZN(n15170) );
  MOAI22 U24084 ( .A1(n28723), .A2(n2850), .B1(ram[10930]), .B2(n2851), 
        .ZN(n15171) );
  MOAI22 U24085 ( .A1(n28488), .A2(n2850), .B1(ram[10931]), .B2(n2851), 
        .ZN(n15172) );
  MOAI22 U24086 ( .A1(n28253), .A2(n2850), .B1(ram[10932]), .B2(n2851), 
        .ZN(n15173) );
  MOAI22 U24087 ( .A1(n28018), .A2(n2850), .B1(ram[10933]), .B2(n2851), 
        .ZN(n15174) );
  MOAI22 U24088 ( .A1(n27783), .A2(n2850), .B1(ram[10934]), .B2(n2851), 
        .ZN(n15175) );
  MOAI22 U24089 ( .A1(n27548), .A2(n2850), .B1(ram[10935]), .B2(n2851), 
        .ZN(n15176) );
  MOAI22 U24090 ( .A1(n29193), .A2(n2852), .B1(ram[10936]), .B2(n2853), 
        .ZN(n15177) );
  MOAI22 U24091 ( .A1(n28958), .A2(n2852), .B1(ram[10937]), .B2(n2853), 
        .ZN(n15178) );
  MOAI22 U24092 ( .A1(n28723), .A2(n2852), .B1(ram[10938]), .B2(n2853), 
        .ZN(n15179) );
  MOAI22 U24093 ( .A1(n28488), .A2(n2852), .B1(ram[10939]), .B2(n2853), 
        .ZN(n15180) );
  MOAI22 U24094 ( .A1(n28253), .A2(n2852), .B1(ram[10940]), .B2(n2853), 
        .ZN(n15181) );
  MOAI22 U24095 ( .A1(n28018), .A2(n2852), .B1(ram[10941]), .B2(n2853), 
        .ZN(n15182) );
  MOAI22 U24096 ( .A1(n27783), .A2(n2852), .B1(ram[10942]), .B2(n2853), 
        .ZN(n15183) );
  MOAI22 U24097 ( .A1(n27548), .A2(n2852), .B1(ram[10943]), .B2(n2853), 
        .ZN(n15184) );
  MOAI22 U24098 ( .A1(n29193), .A2(n2854), .B1(ram[10944]), .B2(n2855), 
        .ZN(n15185) );
  MOAI22 U24099 ( .A1(n28958), .A2(n2854), .B1(ram[10945]), .B2(n2855), 
        .ZN(n15186) );
  MOAI22 U24100 ( .A1(n28723), .A2(n2854), .B1(ram[10946]), .B2(n2855), 
        .ZN(n15187) );
  MOAI22 U24101 ( .A1(n28488), .A2(n2854), .B1(ram[10947]), .B2(n2855), 
        .ZN(n15188) );
  MOAI22 U24102 ( .A1(n28253), .A2(n2854), .B1(ram[10948]), .B2(n2855), 
        .ZN(n15189) );
  MOAI22 U24103 ( .A1(n28018), .A2(n2854), .B1(ram[10949]), .B2(n2855), 
        .ZN(n15190) );
  MOAI22 U24104 ( .A1(n27783), .A2(n2854), .B1(ram[10950]), .B2(n2855), 
        .ZN(n15191) );
  MOAI22 U24105 ( .A1(n27548), .A2(n2854), .B1(ram[10951]), .B2(n2855), 
        .ZN(n15192) );
  MOAI22 U24106 ( .A1(n29193), .A2(n2856), .B1(ram[10952]), .B2(n2857), 
        .ZN(n15193) );
  MOAI22 U24107 ( .A1(n28958), .A2(n2856), .B1(ram[10953]), .B2(n2857), 
        .ZN(n15194) );
  MOAI22 U24108 ( .A1(n28723), .A2(n2856), .B1(ram[10954]), .B2(n2857), 
        .ZN(n15195) );
  MOAI22 U24109 ( .A1(n28488), .A2(n2856), .B1(ram[10955]), .B2(n2857), 
        .ZN(n15196) );
  MOAI22 U24110 ( .A1(n28253), .A2(n2856), .B1(ram[10956]), .B2(n2857), 
        .ZN(n15197) );
  MOAI22 U24111 ( .A1(n28018), .A2(n2856), .B1(ram[10957]), .B2(n2857), 
        .ZN(n15198) );
  MOAI22 U24112 ( .A1(n27783), .A2(n2856), .B1(ram[10958]), .B2(n2857), 
        .ZN(n15199) );
  MOAI22 U24113 ( .A1(n27548), .A2(n2856), .B1(ram[10959]), .B2(n2857), 
        .ZN(n15200) );
  MOAI22 U24114 ( .A1(n29193), .A2(n2858), .B1(ram[10960]), .B2(n2859), 
        .ZN(n15201) );
  MOAI22 U24115 ( .A1(n28958), .A2(n2858), .B1(ram[10961]), .B2(n2859), 
        .ZN(n15202) );
  MOAI22 U24116 ( .A1(n28723), .A2(n2858), .B1(ram[10962]), .B2(n2859), 
        .ZN(n15203) );
  MOAI22 U24117 ( .A1(n28488), .A2(n2858), .B1(ram[10963]), .B2(n2859), 
        .ZN(n15204) );
  MOAI22 U24118 ( .A1(n28253), .A2(n2858), .B1(ram[10964]), .B2(n2859), 
        .ZN(n15205) );
  MOAI22 U24119 ( .A1(n28018), .A2(n2858), .B1(ram[10965]), .B2(n2859), 
        .ZN(n15206) );
  MOAI22 U24120 ( .A1(n27783), .A2(n2858), .B1(ram[10966]), .B2(n2859), 
        .ZN(n15207) );
  MOAI22 U24121 ( .A1(n27548), .A2(n2858), .B1(ram[10967]), .B2(n2859), 
        .ZN(n15208) );
  MOAI22 U24122 ( .A1(n29193), .A2(n2860), .B1(ram[10968]), .B2(n2861), 
        .ZN(n15209) );
  MOAI22 U24123 ( .A1(n28958), .A2(n2860), .B1(ram[10969]), .B2(n2861), 
        .ZN(n15210) );
  MOAI22 U24124 ( .A1(n28723), .A2(n2860), .B1(ram[10970]), .B2(n2861), 
        .ZN(n15211) );
  MOAI22 U24125 ( .A1(n28488), .A2(n2860), .B1(ram[10971]), .B2(n2861), 
        .ZN(n15212) );
  MOAI22 U24126 ( .A1(n28253), .A2(n2860), .B1(ram[10972]), .B2(n2861), 
        .ZN(n15213) );
  MOAI22 U24127 ( .A1(n28018), .A2(n2860), .B1(ram[10973]), .B2(n2861), 
        .ZN(n15214) );
  MOAI22 U24128 ( .A1(n27783), .A2(n2860), .B1(ram[10974]), .B2(n2861), 
        .ZN(n15215) );
  MOAI22 U24129 ( .A1(n27548), .A2(n2860), .B1(ram[10975]), .B2(n2861), 
        .ZN(n15216) );
  MOAI22 U24130 ( .A1(n29193), .A2(n2862), .B1(ram[10976]), .B2(n2863), 
        .ZN(n15217) );
  MOAI22 U24131 ( .A1(n28958), .A2(n2862), .B1(ram[10977]), .B2(n2863), 
        .ZN(n15218) );
  MOAI22 U24132 ( .A1(n28723), .A2(n2862), .B1(ram[10978]), .B2(n2863), 
        .ZN(n15219) );
  MOAI22 U24133 ( .A1(n28488), .A2(n2862), .B1(ram[10979]), .B2(n2863), 
        .ZN(n15220) );
  MOAI22 U24134 ( .A1(n28253), .A2(n2862), .B1(ram[10980]), .B2(n2863), 
        .ZN(n15221) );
  MOAI22 U24135 ( .A1(n28018), .A2(n2862), .B1(ram[10981]), .B2(n2863), 
        .ZN(n15222) );
  MOAI22 U24136 ( .A1(n27783), .A2(n2862), .B1(ram[10982]), .B2(n2863), 
        .ZN(n15223) );
  MOAI22 U24137 ( .A1(n27548), .A2(n2862), .B1(ram[10983]), .B2(n2863), 
        .ZN(n15224) );
  MOAI22 U24138 ( .A1(n29193), .A2(n2864), .B1(ram[10984]), .B2(n2865), 
        .ZN(n15225) );
  MOAI22 U24139 ( .A1(n28958), .A2(n2864), .B1(ram[10985]), .B2(n2865), 
        .ZN(n15226) );
  MOAI22 U24140 ( .A1(n28723), .A2(n2864), .B1(ram[10986]), .B2(n2865), 
        .ZN(n15227) );
  MOAI22 U24141 ( .A1(n28488), .A2(n2864), .B1(ram[10987]), .B2(n2865), 
        .ZN(n15228) );
  MOAI22 U24142 ( .A1(n28253), .A2(n2864), .B1(ram[10988]), .B2(n2865), 
        .ZN(n15229) );
  MOAI22 U24143 ( .A1(n28018), .A2(n2864), .B1(ram[10989]), .B2(n2865), 
        .ZN(n15230) );
  MOAI22 U24144 ( .A1(n27783), .A2(n2864), .B1(ram[10990]), .B2(n2865), 
        .ZN(n15231) );
  MOAI22 U24145 ( .A1(n27548), .A2(n2864), .B1(ram[10991]), .B2(n2865), 
        .ZN(n15232) );
  MOAI22 U24146 ( .A1(n29193), .A2(n2866), .B1(ram[10992]), .B2(n2867), 
        .ZN(n15233) );
  MOAI22 U24147 ( .A1(n28958), .A2(n2866), .B1(ram[10993]), .B2(n2867), 
        .ZN(n15234) );
  MOAI22 U24148 ( .A1(n28723), .A2(n2866), .B1(ram[10994]), .B2(n2867), 
        .ZN(n15235) );
  MOAI22 U24149 ( .A1(n28488), .A2(n2866), .B1(ram[10995]), .B2(n2867), 
        .ZN(n15236) );
  MOAI22 U24150 ( .A1(n28253), .A2(n2866), .B1(ram[10996]), .B2(n2867), 
        .ZN(n15237) );
  MOAI22 U24151 ( .A1(n28018), .A2(n2866), .B1(ram[10997]), .B2(n2867), 
        .ZN(n15238) );
  MOAI22 U24152 ( .A1(n27783), .A2(n2866), .B1(ram[10998]), .B2(n2867), 
        .ZN(n15239) );
  MOAI22 U24153 ( .A1(n27548), .A2(n2866), .B1(ram[10999]), .B2(n2867), 
        .ZN(n15240) );
  MOAI22 U24154 ( .A1(n29193), .A2(n2868), .B1(ram[11000]), .B2(n2869), 
        .ZN(n15241) );
  MOAI22 U24155 ( .A1(n28958), .A2(n2868), .B1(ram[11001]), .B2(n2869), 
        .ZN(n15242) );
  MOAI22 U24156 ( .A1(n28723), .A2(n2868), .B1(ram[11002]), .B2(n2869), 
        .ZN(n15243) );
  MOAI22 U24157 ( .A1(n28488), .A2(n2868), .B1(ram[11003]), .B2(n2869), 
        .ZN(n15244) );
  MOAI22 U24158 ( .A1(n28253), .A2(n2868), .B1(ram[11004]), .B2(n2869), 
        .ZN(n15245) );
  MOAI22 U24159 ( .A1(n28018), .A2(n2868), .B1(ram[11005]), .B2(n2869), 
        .ZN(n15246) );
  MOAI22 U24160 ( .A1(n27783), .A2(n2868), .B1(ram[11006]), .B2(n2869), 
        .ZN(n15247) );
  MOAI22 U24161 ( .A1(n27548), .A2(n2868), .B1(ram[11007]), .B2(n2869), 
        .ZN(n15248) );
  MOAI22 U24162 ( .A1(n29193), .A2(n2870), .B1(ram[11008]), .B2(n2871), 
        .ZN(n15249) );
  MOAI22 U24163 ( .A1(n28958), .A2(n2870), .B1(ram[11009]), .B2(n2871), 
        .ZN(n15250) );
  MOAI22 U24164 ( .A1(n28723), .A2(n2870), .B1(ram[11010]), .B2(n2871), 
        .ZN(n15251) );
  MOAI22 U24165 ( .A1(n28488), .A2(n2870), .B1(ram[11011]), .B2(n2871), 
        .ZN(n15252) );
  MOAI22 U24166 ( .A1(n28253), .A2(n2870), .B1(ram[11012]), .B2(n2871), 
        .ZN(n15253) );
  MOAI22 U24167 ( .A1(n28018), .A2(n2870), .B1(ram[11013]), .B2(n2871), 
        .ZN(n15254) );
  MOAI22 U24168 ( .A1(n27783), .A2(n2870), .B1(ram[11014]), .B2(n2871), 
        .ZN(n15255) );
  MOAI22 U24169 ( .A1(n27548), .A2(n2870), .B1(ram[11015]), .B2(n2871), 
        .ZN(n15256) );
  MOAI22 U24170 ( .A1(n29193), .A2(n2872), .B1(ram[11016]), .B2(n2873), 
        .ZN(n15257) );
  MOAI22 U24171 ( .A1(n28958), .A2(n2872), .B1(ram[11017]), .B2(n2873), 
        .ZN(n15258) );
  MOAI22 U24172 ( .A1(n28723), .A2(n2872), .B1(ram[11018]), .B2(n2873), 
        .ZN(n15259) );
  MOAI22 U24173 ( .A1(n28488), .A2(n2872), .B1(ram[11019]), .B2(n2873), 
        .ZN(n15260) );
  MOAI22 U24174 ( .A1(n28253), .A2(n2872), .B1(ram[11020]), .B2(n2873), 
        .ZN(n15261) );
  MOAI22 U24175 ( .A1(n28018), .A2(n2872), .B1(ram[11021]), .B2(n2873), 
        .ZN(n15262) );
  MOAI22 U24176 ( .A1(n27783), .A2(n2872), .B1(ram[11022]), .B2(n2873), 
        .ZN(n15263) );
  MOAI22 U24177 ( .A1(n27548), .A2(n2872), .B1(ram[11023]), .B2(n2873), 
        .ZN(n15264) );
  MOAI22 U24178 ( .A1(n29194), .A2(n2874), .B1(ram[11024]), .B2(n2875), 
        .ZN(n15265) );
  MOAI22 U24179 ( .A1(n28959), .A2(n2874), .B1(ram[11025]), .B2(n2875), 
        .ZN(n15266) );
  MOAI22 U24180 ( .A1(n28724), .A2(n2874), .B1(ram[11026]), .B2(n2875), 
        .ZN(n15267) );
  MOAI22 U24181 ( .A1(n28489), .A2(n2874), .B1(ram[11027]), .B2(n2875), 
        .ZN(n15268) );
  MOAI22 U24182 ( .A1(n28254), .A2(n2874), .B1(ram[11028]), .B2(n2875), 
        .ZN(n15269) );
  MOAI22 U24183 ( .A1(n28019), .A2(n2874), .B1(ram[11029]), .B2(n2875), 
        .ZN(n15270) );
  MOAI22 U24184 ( .A1(n27784), .A2(n2874), .B1(ram[11030]), .B2(n2875), 
        .ZN(n15271) );
  MOAI22 U24185 ( .A1(n27549), .A2(n2874), .B1(ram[11031]), .B2(n2875), 
        .ZN(n15272) );
  MOAI22 U24186 ( .A1(n29194), .A2(n2876), .B1(ram[11032]), .B2(n2877), 
        .ZN(n15273) );
  MOAI22 U24187 ( .A1(n28959), .A2(n2876), .B1(ram[11033]), .B2(n2877), 
        .ZN(n15274) );
  MOAI22 U24188 ( .A1(n28724), .A2(n2876), .B1(ram[11034]), .B2(n2877), 
        .ZN(n15275) );
  MOAI22 U24189 ( .A1(n28489), .A2(n2876), .B1(ram[11035]), .B2(n2877), 
        .ZN(n15276) );
  MOAI22 U24190 ( .A1(n28254), .A2(n2876), .B1(ram[11036]), .B2(n2877), 
        .ZN(n15277) );
  MOAI22 U24191 ( .A1(n28019), .A2(n2876), .B1(ram[11037]), .B2(n2877), 
        .ZN(n15278) );
  MOAI22 U24192 ( .A1(n27784), .A2(n2876), .B1(ram[11038]), .B2(n2877), 
        .ZN(n15279) );
  MOAI22 U24193 ( .A1(n27549), .A2(n2876), .B1(ram[11039]), .B2(n2877), 
        .ZN(n15280) );
  MOAI22 U24194 ( .A1(n29194), .A2(n2878), .B1(ram[11040]), .B2(n2879), 
        .ZN(n15281) );
  MOAI22 U24195 ( .A1(n28959), .A2(n2878), .B1(ram[11041]), .B2(n2879), 
        .ZN(n15282) );
  MOAI22 U24196 ( .A1(n28724), .A2(n2878), .B1(ram[11042]), .B2(n2879), 
        .ZN(n15283) );
  MOAI22 U24197 ( .A1(n28489), .A2(n2878), .B1(ram[11043]), .B2(n2879), 
        .ZN(n15284) );
  MOAI22 U24198 ( .A1(n28254), .A2(n2878), .B1(ram[11044]), .B2(n2879), 
        .ZN(n15285) );
  MOAI22 U24199 ( .A1(n28019), .A2(n2878), .B1(ram[11045]), .B2(n2879), 
        .ZN(n15286) );
  MOAI22 U24200 ( .A1(n27784), .A2(n2878), .B1(ram[11046]), .B2(n2879), 
        .ZN(n15287) );
  MOAI22 U24201 ( .A1(n27549), .A2(n2878), .B1(ram[11047]), .B2(n2879), 
        .ZN(n15288) );
  MOAI22 U24202 ( .A1(n29194), .A2(n2880), .B1(ram[11048]), .B2(n2881), 
        .ZN(n15289) );
  MOAI22 U24203 ( .A1(n28959), .A2(n2880), .B1(ram[11049]), .B2(n2881), 
        .ZN(n15290) );
  MOAI22 U24204 ( .A1(n28724), .A2(n2880), .B1(ram[11050]), .B2(n2881), 
        .ZN(n15291) );
  MOAI22 U24205 ( .A1(n28489), .A2(n2880), .B1(ram[11051]), .B2(n2881), 
        .ZN(n15292) );
  MOAI22 U24206 ( .A1(n28254), .A2(n2880), .B1(ram[11052]), .B2(n2881), 
        .ZN(n15293) );
  MOAI22 U24207 ( .A1(n28019), .A2(n2880), .B1(ram[11053]), .B2(n2881), 
        .ZN(n15294) );
  MOAI22 U24208 ( .A1(n27784), .A2(n2880), .B1(ram[11054]), .B2(n2881), 
        .ZN(n15295) );
  MOAI22 U24209 ( .A1(n27549), .A2(n2880), .B1(ram[11055]), .B2(n2881), 
        .ZN(n15296) );
  MOAI22 U24210 ( .A1(n29194), .A2(n2882), .B1(ram[11056]), .B2(n2883), 
        .ZN(n15297) );
  MOAI22 U24211 ( .A1(n28959), .A2(n2882), .B1(ram[11057]), .B2(n2883), 
        .ZN(n15298) );
  MOAI22 U24212 ( .A1(n28724), .A2(n2882), .B1(ram[11058]), .B2(n2883), 
        .ZN(n15299) );
  MOAI22 U24213 ( .A1(n28489), .A2(n2882), .B1(ram[11059]), .B2(n2883), 
        .ZN(n15300) );
  MOAI22 U24214 ( .A1(n28254), .A2(n2882), .B1(ram[11060]), .B2(n2883), 
        .ZN(n15301) );
  MOAI22 U24215 ( .A1(n28019), .A2(n2882), .B1(ram[11061]), .B2(n2883), 
        .ZN(n15302) );
  MOAI22 U24216 ( .A1(n27784), .A2(n2882), .B1(ram[11062]), .B2(n2883), 
        .ZN(n15303) );
  MOAI22 U24217 ( .A1(n27549), .A2(n2882), .B1(ram[11063]), .B2(n2883), 
        .ZN(n15304) );
  MOAI22 U24218 ( .A1(n29194), .A2(n2884), .B1(ram[11064]), .B2(n2885), 
        .ZN(n15305) );
  MOAI22 U24219 ( .A1(n28959), .A2(n2884), .B1(ram[11065]), .B2(n2885), 
        .ZN(n15306) );
  MOAI22 U24220 ( .A1(n28724), .A2(n2884), .B1(ram[11066]), .B2(n2885), 
        .ZN(n15307) );
  MOAI22 U24221 ( .A1(n28489), .A2(n2884), .B1(ram[11067]), .B2(n2885), 
        .ZN(n15308) );
  MOAI22 U24222 ( .A1(n28254), .A2(n2884), .B1(ram[11068]), .B2(n2885), 
        .ZN(n15309) );
  MOAI22 U24223 ( .A1(n28019), .A2(n2884), .B1(ram[11069]), .B2(n2885), 
        .ZN(n15310) );
  MOAI22 U24224 ( .A1(n27784), .A2(n2884), .B1(ram[11070]), .B2(n2885), 
        .ZN(n15311) );
  MOAI22 U24225 ( .A1(n27549), .A2(n2884), .B1(ram[11071]), .B2(n2885), 
        .ZN(n15312) );
  MOAI22 U24226 ( .A1(n29194), .A2(n2886), .B1(ram[11072]), .B2(n2887), 
        .ZN(n15313) );
  MOAI22 U24227 ( .A1(n28959), .A2(n2886), .B1(ram[11073]), .B2(n2887), 
        .ZN(n15314) );
  MOAI22 U24228 ( .A1(n28724), .A2(n2886), .B1(ram[11074]), .B2(n2887), 
        .ZN(n15315) );
  MOAI22 U24229 ( .A1(n28489), .A2(n2886), .B1(ram[11075]), .B2(n2887), 
        .ZN(n15316) );
  MOAI22 U24230 ( .A1(n28254), .A2(n2886), .B1(ram[11076]), .B2(n2887), 
        .ZN(n15317) );
  MOAI22 U24231 ( .A1(n28019), .A2(n2886), .B1(ram[11077]), .B2(n2887), 
        .ZN(n15318) );
  MOAI22 U24232 ( .A1(n27784), .A2(n2886), .B1(ram[11078]), .B2(n2887), 
        .ZN(n15319) );
  MOAI22 U24233 ( .A1(n27549), .A2(n2886), .B1(ram[11079]), .B2(n2887), 
        .ZN(n15320) );
  MOAI22 U24234 ( .A1(n29194), .A2(n2888), .B1(ram[11080]), .B2(n2889), 
        .ZN(n15321) );
  MOAI22 U24235 ( .A1(n28959), .A2(n2888), .B1(ram[11081]), .B2(n2889), 
        .ZN(n15322) );
  MOAI22 U24236 ( .A1(n28724), .A2(n2888), .B1(ram[11082]), .B2(n2889), 
        .ZN(n15323) );
  MOAI22 U24237 ( .A1(n28489), .A2(n2888), .B1(ram[11083]), .B2(n2889), 
        .ZN(n15324) );
  MOAI22 U24238 ( .A1(n28254), .A2(n2888), .B1(ram[11084]), .B2(n2889), 
        .ZN(n15325) );
  MOAI22 U24239 ( .A1(n28019), .A2(n2888), .B1(ram[11085]), .B2(n2889), 
        .ZN(n15326) );
  MOAI22 U24240 ( .A1(n27784), .A2(n2888), .B1(ram[11086]), .B2(n2889), 
        .ZN(n15327) );
  MOAI22 U24241 ( .A1(n27549), .A2(n2888), .B1(ram[11087]), .B2(n2889), 
        .ZN(n15328) );
  MOAI22 U24242 ( .A1(n29194), .A2(n2890), .B1(ram[11088]), .B2(n2891), 
        .ZN(n15329) );
  MOAI22 U24243 ( .A1(n28959), .A2(n2890), .B1(ram[11089]), .B2(n2891), 
        .ZN(n15330) );
  MOAI22 U24244 ( .A1(n28724), .A2(n2890), .B1(ram[11090]), .B2(n2891), 
        .ZN(n15331) );
  MOAI22 U24245 ( .A1(n28489), .A2(n2890), .B1(ram[11091]), .B2(n2891), 
        .ZN(n15332) );
  MOAI22 U24246 ( .A1(n28254), .A2(n2890), .B1(ram[11092]), .B2(n2891), 
        .ZN(n15333) );
  MOAI22 U24247 ( .A1(n28019), .A2(n2890), .B1(ram[11093]), .B2(n2891), 
        .ZN(n15334) );
  MOAI22 U24248 ( .A1(n27784), .A2(n2890), .B1(ram[11094]), .B2(n2891), 
        .ZN(n15335) );
  MOAI22 U24249 ( .A1(n27549), .A2(n2890), .B1(ram[11095]), .B2(n2891), 
        .ZN(n15336) );
  MOAI22 U24250 ( .A1(n29194), .A2(n2892), .B1(ram[11096]), .B2(n2893), 
        .ZN(n15337) );
  MOAI22 U24251 ( .A1(n28959), .A2(n2892), .B1(ram[11097]), .B2(n2893), 
        .ZN(n15338) );
  MOAI22 U24252 ( .A1(n28724), .A2(n2892), .B1(ram[11098]), .B2(n2893), 
        .ZN(n15339) );
  MOAI22 U24253 ( .A1(n28489), .A2(n2892), .B1(ram[11099]), .B2(n2893), 
        .ZN(n15340) );
  MOAI22 U24254 ( .A1(n28254), .A2(n2892), .B1(ram[11100]), .B2(n2893), 
        .ZN(n15341) );
  MOAI22 U24255 ( .A1(n28019), .A2(n2892), .B1(ram[11101]), .B2(n2893), 
        .ZN(n15342) );
  MOAI22 U24256 ( .A1(n27784), .A2(n2892), .B1(ram[11102]), .B2(n2893), 
        .ZN(n15343) );
  MOAI22 U24257 ( .A1(n27549), .A2(n2892), .B1(ram[11103]), .B2(n2893), 
        .ZN(n15344) );
  MOAI22 U24258 ( .A1(n29194), .A2(n2894), .B1(ram[11104]), .B2(n2895), 
        .ZN(n15345) );
  MOAI22 U24259 ( .A1(n28959), .A2(n2894), .B1(ram[11105]), .B2(n2895), 
        .ZN(n15346) );
  MOAI22 U24260 ( .A1(n28724), .A2(n2894), .B1(ram[11106]), .B2(n2895), 
        .ZN(n15347) );
  MOAI22 U24261 ( .A1(n28489), .A2(n2894), .B1(ram[11107]), .B2(n2895), 
        .ZN(n15348) );
  MOAI22 U24262 ( .A1(n28254), .A2(n2894), .B1(ram[11108]), .B2(n2895), 
        .ZN(n15349) );
  MOAI22 U24263 ( .A1(n28019), .A2(n2894), .B1(ram[11109]), .B2(n2895), 
        .ZN(n15350) );
  MOAI22 U24264 ( .A1(n27784), .A2(n2894), .B1(ram[11110]), .B2(n2895), 
        .ZN(n15351) );
  MOAI22 U24265 ( .A1(n27549), .A2(n2894), .B1(ram[11111]), .B2(n2895), 
        .ZN(n15352) );
  MOAI22 U24266 ( .A1(n29194), .A2(n2896), .B1(ram[11112]), .B2(n2897), 
        .ZN(n15353) );
  MOAI22 U24267 ( .A1(n28959), .A2(n2896), .B1(ram[11113]), .B2(n2897), 
        .ZN(n15354) );
  MOAI22 U24268 ( .A1(n28724), .A2(n2896), .B1(ram[11114]), .B2(n2897), 
        .ZN(n15355) );
  MOAI22 U24269 ( .A1(n28489), .A2(n2896), .B1(ram[11115]), .B2(n2897), 
        .ZN(n15356) );
  MOAI22 U24270 ( .A1(n28254), .A2(n2896), .B1(ram[11116]), .B2(n2897), 
        .ZN(n15357) );
  MOAI22 U24271 ( .A1(n28019), .A2(n2896), .B1(ram[11117]), .B2(n2897), 
        .ZN(n15358) );
  MOAI22 U24272 ( .A1(n27784), .A2(n2896), .B1(ram[11118]), .B2(n2897), 
        .ZN(n15359) );
  MOAI22 U24273 ( .A1(n27549), .A2(n2896), .B1(ram[11119]), .B2(n2897), 
        .ZN(n15360) );
  MOAI22 U24274 ( .A1(n29194), .A2(n2898), .B1(ram[11120]), .B2(n2899), 
        .ZN(n15361) );
  MOAI22 U24275 ( .A1(n28959), .A2(n2898), .B1(ram[11121]), .B2(n2899), 
        .ZN(n15362) );
  MOAI22 U24276 ( .A1(n28724), .A2(n2898), .B1(ram[11122]), .B2(n2899), 
        .ZN(n15363) );
  MOAI22 U24277 ( .A1(n28489), .A2(n2898), .B1(ram[11123]), .B2(n2899), 
        .ZN(n15364) );
  MOAI22 U24278 ( .A1(n28254), .A2(n2898), .B1(ram[11124]), .B2(n2899), 
        .ZN(n15365) );
  MOAI22 U24279 ( .A1(n28019), .A2(n2898), .B1(ram[11125]), .B2(n2899), 
        .ZN(n15366) );
  MOAI22 U24280 ( .A1(n27784), .A2(n2898), .B1(ram[11126]), .B2(n2899), 
        .ZN(n15367) );
  MOAI22 U24281 ( .A1(n27549), .A2(n2898), .B1(ram[11127]), .B2(n2899), 
        .ZN(n15368) );
  MOAI22 U24282 ( .A1(n29195), .A2(n2900), .B1(ram[11128]), .B2(n2901), 
        .ZN(n15369) );
  MOAI22 U24283 ( .A1(n28960), .A2(n2900), .B1(ram[11129]), .B2(n2901), 
        .ZN(n15370) );
  MOAI22 U24284 ( .A1(n28725), .A2(n2900), .B1(ram[11130]), .B2(n2901), 
        .ZN(n15371) );
  MOAI22 U24285 ( .A1(n28490), .A2(n2900), .B1(ram[11131]), .B2(n2901), 
        .ZN(n15372) );
  MOAI22 U24286 ( .A1(n28255), .A2(n2900), .B1(ram[11132]), .B2(n2901), 
        .ZN(n15373) );
  MOAI22 U24287 ( .A1(n28020), .A2(n2900), .B1(ram[11133]), .B2(n2901), 
        .ZN(n15374) );
  MOAI22 U24288 ( .A1(n27785), .A2(n2900), .B1(ram[11134]), .B2(n2901), 
        .ZN(n15375) );
  MOAI22 U24289 ( .A1(n27550), .A2(n2900), .B1(ram[11135]), .B2(n2901), 
        .ZN(n15376) );
  MOAI22 U24290 ( .A1(n29195), .A2(n2902), .B1(ram[11136]), .B2(n2903), 
        .ZN(n15377) );
  MOAI22 U24291 ( .A1(n28960), .A2(n2902), .B1(ram[11137]), .B2(n2903), 
        .ZN(n15378) );
  MOAI22 U24292 ( .A1(n28725), .A2(n2902), .B1(ram[11138]), .B2(n2903), 
        .ZN(n15379) );
  MOAI22 U24293 ( .A1(n28490), .A2(n2902), .B1(ram[11139]), .B2(n2903), 
        .ZN(n15380) );
  MOAI22 U24294 ( .A1(n28255), .A2(n2902), .B1(ram[11140]), .B2(n2903), 
        .ZN(n15381) );
  MOAI22 U24295 ( .A1(n28020), .A2(n2902), .B1(ram[11141]), .B2(n2903), 
        .ZN(n15382) );
  MOAI22 U24296 ( .A1(n27785), .A2(n2902), .B1(ram[11142]), .B2(n2903), 
        .ZN(n15383) );
  MOAI22 U24297 ( .A1(n27550), .A2(n2902), .B1(ram[11143]), .B2(n2903), 
        .ZN(n15384) );
  MOAI22 U24298 ( .A1(n29195), .A2(n2904), .B1(ram[11144]), .B2(n2905), 
        .ZN(n15385) );
  MOAI22 U24299 ( .A1(n28960), .A2(n2904), .B1(ram[11145]), .B2(n2905), 
        .ZN(n15386) );
  MOAI22 U24300 ( .A1(n28725), .A2(n2904), .B1(ram[11146]), .B2(n2905), 
        .ZN(n15387) );
  MOAI22 U24301 ( .A1(n28490), .A2(n2904), .B1(ram[11147]), .B2(n2905), 
        .ZN(n15388) );
  MOAI22 U24302 ( .A1(n28255), .A2(n2904), .B1(ram[11148]), .B2(n2905), 
        .ZN(n15389) );
  MOAI22 U24303 ( .A1(n28020), .A2(n2904), .B1(ram[11149]), .B2(n2905), 
        .ZN(n15390) );
  MOAI22 U24304 ( .A1(n27785), .A2(n2904), .B1(ram[11150]), .B2(n2905), 
        .ZN(n15391) );
  MOAI22 U24305 ( .A1(n27550), .A2(n2904), .B1(ram[11151]), .B2(n2905), 
        .ZN(n15392) );
  MOAI22 U24306 ( .A1(n29195), .A2(n2906), .B1(ram[11152]), .B2(n2907), 
        .ZN(n15393) );
  MOAI22 U24307 ( .A1(n28960), .A2(n2906), .B1(ram[11153]), .B2(n2907), 
        .ZN(n15394) );
  MOAI22 U24308 ( .A1(n28725), .A2(n2906), .B1(ram[11154]), .B2(n2907), 
        .ZN(n15395) );
  MOAI22 U24309 ( .A1(n28490), .A2(n2906), .B1(ram[11155]), .B2(n2907), 
        .ZN(n15396) );
  MOAI22 U24310 ( .A1(n28255), .A2(n2906), .B1(ram[11156]), .B2(n2907), 
        .ZN(n15397) );
  MOAI22 U24311 ( .A1(n28020), .A2(n2906), .B1(ram[11157]), .B2(n2907), 
        .ZN(n15398) );
  MOAI22 U24312 ( .A1(n27785), .A2(n2906), .B1(ram[11158]), .B2(n2907), 
        .ZN(n15399) );
  MOAI22 U24313 ( .A1(n27550), .A2(n2906), .B1(ram[11159]), .B2(n2907), 
        .ZN(n15400) );
  MOAI22 U24314 ( .A1(n29195), .A2(n2908), .B1(ram[11160]), .B2(n2909), 
        .ZN(n15401) );
  MOAI22 U24315 ( .A1(n28960), .A2(n2908), .B1(ram[11161]), .B2(n2909), 
        .ZN(n15402) );
  MOAI22 U24316 ( .A1(n28725), .A2(n2908), .B1(ram[11162]), .B2(n2909), 
        .ZN(n15403) );
  MOAI22 U24317 ( .A1(n28490), .A2(n2908), .B1(ram[11163]), .B2(n2909), 
        .ZN(n15404) );
  MOAI22 U24318 ( .A1(n28255), .A2(n2908), .B1(ram[11164]), .B2(n2909), 
        .ZN(n15405) );
  MOAI22 U24319 ( .A1(n28020), .A2(n2908), .B1(ram[11165]), .B2(n2909), 
        .ZN(n15406) );
  MOAI22 U24320 ( .A1(n27785), .A2(n2908), .B1(ram[11166]), .B2(n2909), 
        .ZN(n15407) );
  MOAI22 U24321 ( .A1(n27550), .A2(n2908), .B1(ram[11167]), .B2(n2909), 
        .ZN(n15408) );
  MOAI22 U24322 ( .A1(n29195), .A2(n2910), .B1(ram[11168]), .B2(n2911), 
        .ZN(n15409) );
  MOAI22 U24323 ( .A1(n28960), .A2(n2910), .B1(ram[11169]), .B2(n2911), 
        .ZN(n15410) );
  MOAI22 U24324 ( .A1(n28725), .A2(n2910), .B1(ram[11170]), .B2(n2911), 
        .ZN(n15411) );
  MOAI22 U24325 ( .A1(n28490), .A2(n2910), .B1(ram[11171]), .B2(n2911), 
        .ZN(n15412) );
  MOAI22 U24326 ( .A1(n28255), .A2(n2910), .B1(ram[11172]), .B2(n2911), 
        .ZN(n15413) );
  MOAI22 U24327 ( .A1(n28020), .A2(n2910), .B1(ram[11173]), .B2(n2911), 
        .ZN(n15414) );
  MOAI22 U24328 ( .A1(n27785), .A2(n2910), .B1(ram[11174]), .B2(n2911), 
        .ZN(n15415) );
  MOAI22 U24329 ( .A1(n27550), .A2(n2910), .B1(ram[11175]), .B2(n2911), 
        .ZN(n15416) );
  MOAI22 U24330 ( .A1(n29195), .A2(n2912), .B1(ram[11176]), .B2(n2913), 
        .ZN(n15417) );
  MOAI22 U24331 ( .A1(n28960), .A2(n2912), .B1(ram[11177]), .B2(n2913), 
        .ZN(n15418) );
  MOAI22 U24332 ( .A1(n28725), .A2(n2912), .B1(ram[11178]), .B2(n2913), 
        .ZN(n15419) );
  MOAI22 U24333 ( .A1(n28490), .A2(n2912), .B1(ram[11179]), .B2(n2913), 
        .ZN(n15420) );
  MOAI22 U24334 ( .A1(n28255), .A2(n2912), .B1(ram[11180]), .B2(n2913), 
        .ZN(n15421) );
  MOAI22 U24335 ( .A1(n28020), .A2(n2912), .B1(ram[11181]), .B2(n2913), 
        .ZN(n15422) );
  MOAI22 U24336 ( .A1(n27785), .A2(n2912), .B1(ram[11182]), .B2(n2913), 
        .ZN(n15423) );
  MOAI22 U24337 ( .A1(n27550), .A2(n2912), .B1(ram[11183]), .B2(n2913), 
        .ZN(n15424) );
  MOAI22 U24338 ( .A1(n29195), .A2(n2914), .B1(ram[11184]), .B2(n2915), 
        .ZN(n15425) );
  MOAI22 U24339 ( .A1(n28960), .A2(n2914), .B1(ram[11185]), .B2(n2915), 
        .ZN(n15426) );
  MOAI22 U24340 ( .A1(n28725), .A2(n2914), .B1(ram[11186]), .B2(n2915), 
        .ZN(n15427) );
  MOAI22 U24341 ( .A1(n28490), .A2(n2914), .B1(ram[11187]), .B2(n2915), 
        .ZN(n15428) );
  MOAI22 U24342 ( .A1(n28255), .A2(n2914), .B1(ram[11188]), .B2(n2915), 
        .ZN(n15429) );
  MOAI22 U24343 ( .A1(n28020), .A2(n2914), .B1(ram[11189]), .B2(n2915), 
        .ZN(n15430) );
  MOAI22 U24344 ( .A1(n27785), .A2(n2914), .B1(ram[11190]), .B2(n2915), 
        .ZN(n15431) );
  MOAI22 U24345 ( .A1(n27550), .A2(n2914), .B1(ram[11191]), .B2(n2915), 
        .ZN(n15432) );
  MOAI22 U24346 ( .A1(n29195), .A2(n2916), .B1(ram[11192]), .B2(n2917), 
        .ZN(n15433) );
  MOAI22 U24347 ( .A1(n28960), .A2(n2916), .B1(ram[11193]), .B2(n2917), 
        .ZN(n15434) );
  MOAI22 U24348 ( .A1(n28725), .A2(n2916), .B1(ram[11194]), .B2(n2917), 
        .ZN(n15435) );
  MOAI22 U24349 ( .A1(n28490), .A2(n2916), .B1(ram[11195]), .B2(n2917), 
        .ZN(n15436) );
  MOAI22 U24350 ( .A1(n28255), .A2(n2916), .B1(ram[11196]), .B2(n2917), 
        .ZN(n15437) );
  MOAI22 U24351 ( .A1(n28020), .A2(n2916), .B1(ram[11197]), .B2(n2917), 
        .ZN(n15438) );
  MOAI22 U24352 ( .A1(n27785), .A2(n2916), .B1(ram[11198]), .B2(n2917), 
        .ZN(n15439) );
  MOAI22 U24353 ( .A1(n27550), .A2(n2916), .B1(ram[11199]), .B2(n2917), 
        .ZN(n15440) );
  MOAI22 U24354 ( .A1(n29195), .A2(n2918), .B1(ram[11200]), .B2(n2919), 
        .ZN(n15441) );
  MOAI22 U24355 ( .A1(n28960), .A2(n2918), .B1(ram[11201]), .B2(n2919), 
        .ZN(n15442) );
  MOAI22 U24356 ( .A1(n28725), .A2(n2918), .B1(ram[11202]), .B2(n2919), 
        .ZN(n15443) );
  MOAI22 U24357 ( .A1(n28490), .A2(n2918), .B1(ram[11203]), .B2(n2919), 
        .ZN(n15444) );
  MOAI22 U24358 ( .A1(n28255), .A2(n2918), .B1(ram[11204]), .B2(n2919), 
        .ZN(n15445) );
  MOAI22 U24359 ( .A1(n28020), .A2(n2918), .B1(ram[11205]), .B2(n2919), 
        .ZN(n15446) );
  MOAI22 U24360 ( .A1(n27785), .A2(n2918), .B1(ram[11206]), .B2(n2919), 
        .ZN(n15447) );
  MOAI22 U24361 ( .A1(n27550), .A2(n2918), .B1(ram[11207]), .B2(n2919), 
        .ZN(n15448) );
  MOAI22 U24362 ( .A1(n29195), .A2(n2920), .B1(ram[11208]), .B2(n2921), 
        .ZN(n15449) );
  MOAI22 U24363 ( .A1(n28960), .A2(n2920), .B1(ram[11209]), .B2(n2921), 
        .ZN(n15450) );
  MOAI22 U24364 ( .A1(n28725), .A2(n2920), .B1(ram[11210]), .B2(n2921), 
        .ZN(n15451) );
  MOAI22 U24365 ( .A1(n28490), .A2(n2920), .B1(ram[11211]), .B2(n2921), 
        .ZN(n15452) );
  MOAI22 U24366 ( .A1(n28255), .A2(n2920), .B1(ram[11212]), .B2(n2921), 
        .ZN(n15453) );
  MOAI22 U24367 ( .A1(n28020), .A2(n2920), .B1(ram[11213]), .B2(n2921), 
        .ZN(n15454) );
  MOAI22 U24368 ( .A1(n27785), .A2(n2920), .B1(ram[11214]), .B2(n2921), 
        .ZN(n15455) );
  MOAI22 U24369 ( .A1(n27550), .A2(n2920), .B1(ram[11215]), .B2(n2921), 
        .ZN(n15456) );
  MOAI22 U24370 ( .A1(n29195), .A2(n2922), .B1(ram[11216]), .B2(n2923), 
        .ZN(n15457) );
  MOAI22 U24371 ( .A1(n28960), .A2(n2922), .B1(ram[11217]), .B2(n2923), 
        .ZN(n15458) );
  MOAI22 U24372 ( .A1(n28725), .A2(n2922), .B1(ram[11218]), .B2(n2923), 
        .ZN(n15459) );
  MOAI22 U24373 ( .A1(n28490), .A2(n2922), .B1(ram[11219]), .B2(n2923), 
        .ZN(n15460) );
  MOAI22 U24374 ( .A1(n28255), .A2(n2922), .B1(ram[11220]), .B2(n2923), 
        .ZN(n15461) );
  MOAI22 U24375 ( .A1(n28020), .A2(n2922), .B1(ram[11221]), .B2(n2923), 
        .ZN(n15462) );
  MOAI22 U24376 ( .A1(n27785), .A2(n2922), .B1(ram[11222]), .B2(n2923), 
        .ZN(n15463) );
  MOAI22 U24377 ( .A1(n27550), .A2(n2922), .B1(ram[11223]), .B2(n2923), 
        .ZN(n15464) );
  MOAI22 U24378 ( .A1(n29195), .A2(n2924), .B1(ram[11224]), .B2(n2925), 
        .ZN(n15465) );
  MOAI22 U24379 ( .A1(n28960), .A2(n2924), .B1(ram[11225]), .B2(n2925), 
        .ZN(n15466) );
  MOAI22 U24380 ( .A1(n28725), .A2(n2924), .B1(ram[11226]), .B2(n2925), 
        .ZN(n15467) );
  MOAI22 U24381 ( .A1(n28490), .A2(n2924), .B1(ram[11227]), .B2(n2925), 
        .ZN(n15468) );
  MOAI22 U24382 ( .A1(n28255), .A2(n2924), .B1(ram[11228]), .B2(n2925), 
        .ZN(n15469) );
  MOAI22 U24383 ( .A1(n28020), .A2(n2924), .B1(ram[11229]), .B2(n2925), 
        .ZN(n15470) );
  MOAI22 U24384 ( .A1(n27785), .A2(n2924), .B1(ram[11230]), .B2(n2925), 
        .ZN(n15471) );
  MOAI22 U24385 ( .A1(n27550), .A2(n2924), .B1(ram[11231]), .B2(n2925), 
        .ZN(n15472) );
  MOAI22 U24386 ( .A1(n29196), .A2(n2926), .B1(ram[11232]), .B2(n2927), 
        .ZN(n15473) );
  MOAI22 U24387 ( .A1(n28961), .A2(n2926), .B1(ram[11233]), .B2(n2927), 
        .ZN(n15474) );
  MOAI22 U24388 ( .A1(n28726), .A2(n2926), .B1(ram[11234]), .B2(n2927), 
        .ZN(n15475) );
  MOAI22 U24389 ( .A1(n28491), .A2(n2926), .B1(ram[11235]), .B2(n2927), 
        .ZN(n15476) );
  MOAI22 U24390 ( .A1(n28256), .A2(n2926), .B1(ram[11236]), .B2(n2927), 
        .ZN(n15477) );
  MOAI22 U24391 ( .A1(n28021), .A2(n2926), .B1(ram[11237]), .B2(n2927), 
        .ZN(n15478) );
  MOAI22 U24392 ( .A1(n27786), .A2(n2926), .B1(ram[11238]), .B2(n2927), 
        .ZN(n15479) );
  MOAI22 U24393 ( .A1(n27551), .A2(n2926), .B1(ram[11239]), .B2(n2927), 
        .ZN(n15480) );
  MOAI22 U24394 ( .A1(n29196), .A2(n2928), .B1(ram[11240]), .B2(n2929), 
        .ZN(n15481) );
  MOAI22 U24395 ( .A1(n28961), .A2(n2928), .B1(ram[11241]), .B2(n2929), 
        .ZN(n15482) );
  MOAI22 U24396 ( .A1(n28726), .A2(n2928), .B1(ram[11242]), .B2(n2929), 
        .ZN(n15483) );
  MOAI22 U24397 ( .A1(n28491), .A2(n2928), .B1(ram[11243]), .B2(n2929), 
        .ZN(n15484) );
  MOAI22 U24398 ( .A1(n28256), .A2(n2928), .B1(ram[11244]), .B2(n2929), 
        .ZN(n15485) );
  MOAI22 U24399 ( .A1(n28021), .A2(n2928), .B1(ram[11245]), .B2(n2929), 
        .ZN(n15486) );
  MOAI22 U24400 ( .A1(n27786), .A2(n2928), .B1(ram[11246]), .B2(n2929), 
        .ZN(n15487) );
  MOAI22 U24401 ( .A1(n27551), .A2(n2928), .B1(ram[11247]), .B2(n2929), 
        .ZN(n15488) );
  MOAI22 U24402 ( .A1(n29196), .A2(n2930), .B1(ram[11248]), .B2(n2931), 
        .ZN(n15489) );
  MOAI22 U24403 ( .A1(n28961), .A2(n2930), .B1(ram[11249]), .B2(n2931), 
        .ZN(n15490) );
  MOAI22 U24404 ( .A1(n28726), .A2(n2930), .B1(ram[11250]), .B2(n2931), 
        .ZN(n15491) );
  MOAI22 U24405 ( .A1(n28491), .A2(n2930), .B1(ram[11251]), .B2(n2931), 
        .ZN(n15492) );
  MOAI22 U24406 ( .A1(n28256), .A2(n2930), .B1(ram[11252]), .B2(n2931), 
        .ZN(n15493) );
  MOAI22 U24407 ( .A1(n28021), .A2(n2930), .B1(ram[11253]), .B2(n2931), 
        .ZN(n15494) );
  MOAI22 U24408 ( .A1(n27786), .A2(n2930), .B1(ram[11254]), .B2(n2931), 
        .ZN(n15495) );
  MOAI22 U24409 ( .A1(n27551), .A2(n2930), .B1(ram[11255]), .B2(n2931), 
        .ZN(n15496) );
  MOAI22 U24410 ( .A1(n29196), .A2(n2932), .B1(ram[11256]), .B2(n2933), 
        .ZN(n15497) );
  MOAI22 U24411 ( .A1(n28961), .A2(n2932), .B1(ram[11257]), .B2(n2933), 
        .ZN(n15498) );
  MOAI22 U24412 ( .A1(n28726), .A2(n2932), .B1(ram[11258]), .B2(n2933), 
        .ZN(n15499) );
  MOAI22 U24413 ( .A1(n28491), .A2(n2932), .B1(ram[11259]), .B2(n2933), 
        .ZN(n15500) );
  MOAI22 U24414 ( .A1(n28256), .A2(n2932), .B1(ram[11260]), .B2(n2933), 
        .ZN(n15501) );
  MOAI22 U24415 ( .A1(n28021), .A2(n2932), .B1(ram[11261]), .B2(n2933), 
        .ZN(n15502) );
  MOAI22 U24416 ( .A1(n27786), .A2(n2932), .B1(ram[11262]), .B2(n2933), 
        .ZN(n15503) );
  MOAI22 U24417 ( .A1(n27551), .A2(n2932), .B1(ram[11263]), .B2(n2933), 
        .ZN(n15504) );
  MOAI22 U24418 ( .A1(n29196), .A2(n2934), .B1(ram[11264]), .B2(n2935), 
        .ZN(n15505) );
  MOAI22 U24419 ( .A1(n28961), .A2(n2934), .B1(ram[11265]), .B2(n2935), 
        .ZN(n15506) );
  MOAI22 U24420 ( .A1(n28726), .A2(n2934), .B1(ram[11266]), .B2(n2935), 
        .ZN(n15507) );
  MOAI22 U24421 ( .A1(n28491), .A2(n2934), .B1(ram[11267]), .B2(n2935), 
        .ZN(n15508) );
  MOAI22 U24422 ( .A1(n28256), .A2(n2934), .B1(ram[11268]), .B2(n2935), 
        .ZN(n15509) );
  MOAI22 U24423 ( .A1(n28021), .A2(n2934), .B1(ram[11269]), .B2(n2935), 
        .ZN(n15510) );
  MOAI22 U24424 ( .A1(n27786), .A2(n2934), .B1(ram[11270]), .B2(n2935), 
        .ZN(n15511) );
  MOAI22 U24425 ( .A1(n27551), .A2(n2934), .B1(ram[11271]), .B2(n2935), 
        .ZN(n15512) );
  MOAI22 U24426 ( .A1(n29196), .A2(n2937), .B1(ram[11272]), .B2(n2938), 
        .ZN(n15513) );
  MOAI22 U24427 ( .A1(n28961), .A2(n2937), .B1(ram[11273]), .B2(n2938), 
        .ZN(n15514) );
  MOAI22 U24428 ( .A1(n28726), .A2(n2937), .B1(ram[11274]), .B2(n2938), 
        .ZN(n15515) );
  MOAI22 U24429 ( .A1(n28491), .A2(n2937), .B1(ram[11275]), .B2(n2938), 
        .ZN(n15516) );
  MOAI22 U24430 ( .A1(n28256), .A2(n2937), .B1(ram[11276]), .B2(n2938), 
        .ZN(n15517) );
  MOAI22 U24431 ( .A1(n28021), .A2(n2937), .B1(ram[11277]), .B2(n2938), 
        .ZN(n15518) );
  MOAI22 U24432 ( .A1(n27786), .A2(n2937), .B1(ram[11278]), .B2(n2938), 
        .ZN(n15519) );
  MOAI22 U24433 ( .A1(n27551), .A2(n2937), .B1(ram[11279]), .B2(n2938), 
        .ZN(n15520) );
  MOAI22 U24434 ( .A1(n29196), .A2(n2939), .B1(ram[11280]), .B2(n2940), 
        .ZN(n15521) );
  MOAI22 U24435 ( .A1(n28961), .A2(n2939), .B1(ram[11281]), .B2(n2940), 
        .ZN(n15522) );
  MOAI22 U24436 ( .A1(n28726), .A2(n2939), .B1(ram[11282]), .B2(n2940), 
        .ZN(n15523) );
  MOAI22 U24437 ( .A1(n28491), .A2(n2939), .B1(ram[11283]), .B2(n2940), 
        .ZN(n15524) );
  MOAI22 U24438 ( .A1(n28256), .A2(n2939), .B1(ram[11284]), .B2(n2940), 
        .ZN(n15525) );
  MOAI22 U24439 ( .A1(n28021), .A2(n2939), .B1(ram[11285]), .B2(n2940), 
        .ZN(n15526) );
  MOAI22 U24440 ( .A1(n27786), .A2(n2939), .B1(ram[11286]), .B2(n2940), 
        .ZN(n15527) );
  MOAI22 U24441 ( .A1(n27551), .A2(n2939), .B1(ram[11287]), .B2(n2940), 
        .ZN(n15528) );
  MOAI22 U24442 ( .A1(n29196), .A2(n2941), .B1(ram[11288]), .B2(n2942), 
        .ZN(n15529) );
  MOAI22 U24443 ( .A1(n28961), .A2(n2941), .B1(ram[11289]), .B2(n2942), 
        .ZN(n15530) );
  MOAI22 U24444 ( .A1(n28726), .A2(n2941), .B1(ram[11290]), .B2(n2942), 
        .ZN(n15531) );
  MOAI22 U24445 ( .A1(n28491), .A2(n2941), .B1(ram[11291]), .B2(n2942), 
        .ZN(n15532) );
  MOAI22 U24446 ( .A1(n28256), .A2(n2941), .B1(ram[11292]), .B2(n2942), 
        .ZN(n15533) );
  MOAI22 U24447 ( .A1(n28021), .A2(n2941), .B1(ram[11293]), .B2(n2942), 
        .ZN(n15534) );
  MOAI22 U24448 ( .A1(n27786), .A2(n2941), .B1(ram[11294]), .B2(n2942), 
        .ZN(n15535) );
  MOAI22 U24449 ( .A1(n27551), .A2(n2941), .B1(ram[11295]), .B2(n2942), 
        .ZN(n15536) );
  MOAI22 U24450 ( .A1(n29196), .A2(n2943), .B1(ram[11296]), .B2(n2944), 
        .ZN(n15537) );
  MOAI22 U24451 ( .A1(n28961), .A2(n2943), .B1(ram[11297]), .B2(n2944), 
        .ZN(n15538) );
  MOAI22 U24452 ( .A1(n28726), .A2(n2943), .B1(ram[11298]), .B2(n2944), 
        .ZN(n15539) );
  MOAI22 U24453 ( .A1(n28491), .A2(n2943), .B1(ram[11299]), .B2(n2944), 
        .ZN(n15540) );
  MOAI22 U24454 ( .A1(n28256), .A2(n2943), .B1(ram[11300]), .B2(n2944), 
        .ZN(n15541) );
  MOAI22 U24455 ( .A1(n28021), .A2(n2943), .B1(ram[11301]), .B2(n2944), 
        .ZN(n15542) );
  MOAI22 U24456 ( .A1(n27786), .A2(n2943), .B1(ram[11302]), .B2(n2944), 
        .ZN(n15543) );
  MOAI22 U24457 ( .A1(n27551), .A2(n2943), .B1(ram[11303]), .B2(n2944), 
        .ZN(n15544) );
  MOAI22 U24458 ( .A1(n29196), .A2(n2945), .B1(ram[11304]), .B2(n2946), 
        .ZN(n15545) );
  MOAI22 U24459 ( .A1(n28961), .A2(n2945), .B1(ram[11305]), .B2(n2946), 
        .ZN(n15546) );
  MOAI22 U24460 ( .A1(n28726), .A2(n2945), .B1(ram[11306]), .B2(n2946), 
        .ZN(n15547) );
  MOAI22 U24461 ( .A1(n28491), .A2(n2945), .B1(ram[11307]), .B2(n2946), 
        .ZN(n15548) );
  MOAI22 U24462 ( .A1(n28256), .A2(n2945), .B1(ram[11308]), .B2(n2946), 
        .ZN(n15549) );
  MOAI22 U24463 ( .A1(n28021), .A2(n2945), .B1(ram[11309]), .B2(n2946), 
        .ZN(n15550) );
  MOAI22 U24464 ( .A1(n27786), .A2(n2945), .B1(ram[11310]), .B2(n2946), 
        .ZN(n15551) );
  MOAI22 U24465 ( .A1(n27551), .A2(n2945), .B1(ram[11311]), .B2(n2946), 
        .ZN(n15552) );
  MOAI22 U24466 ( .A1(n29196), .A2(n2947), .B1(ram[11312]), .B2(n2948), 
        .ZN(n15553) );
  MOAI22 U24467 ( .A1(n28961), .A2(n2947), .B1(ram[11313]), .B2(n2948), 
        .ZN(n15554) );
  MOAI22 U24468 ( .A1(n28726), .A2(n2947), .B1(ram[11314]), .B2(n2948), 
        .ZN(n15555) );
  MOAI22 U24469 ( .A1(n28491), .A2(n2947), .B1(ram[11315]), .B2(n2948), 
        .ZN(n15556) );
  MOAI22 U24470 ( .A1(n28256), .A2(n2947), .B1(ram[11316]), .B2(n2948), 
        .ZN(n15557) );
  MOAI22 U24471 ( .A1(n28021), .A2(n2947), .B1(ram[11317]), .B2(n2948), 
        .ZN(n15558) );
  MOAI22 U24472 ( .A1(n27786), .A2(n2947), .B1(ram[11318]), .B2(n2948), 
        .ZN(n15559) );
  MOAI22 U24473 ( .A1(n27551), .A2(n2947), .B1(ram[11319]), .B2(n2948), 
        .ZN(n15560) );
  MOAI22 U24474 ( .A1(n29196), .A2(n2949), .B1(ram[11320]), .B2(n2950), 
        .ZN(n15561) );
  MOAI22 U24475 ( .A1(n28961), .A2(n2949), .B1(ram[11321]), .B2(n2950), 
        .ZN(n15562) );
  MOAI22 U24476 ( .A1(n28726), .A2(n2949), .B1(ram[11322]), .B2(n2950), 
        .ZN(n15563) );
  MOAI22 U24477 ( .A1(n28491), .A2(n2949), .B1(ram[11323]), .B2(n2950), 
        .ZN(n15564) );
  MOAI22 U24478 ( .A1(n28256), .A2(n2949), .B1(ram[11324]), .B2(n2950), 
        .ZN(n15565) );
  MOAI22 U24479 ( .A1(n28021), .A2(n2949), .B1(ram[11325]), .B2(n2950), 
        .ZN(n15566) );
  MOAI22 U24480 ( .A1(n27786), .A2(n2949), .B1(ram[11326]), .B2(n2950), 
        .ZN(n15567) );
  MOAI22 U24481 ( .A1(n27551), .A2(n2949), .B1(ram[11327]), .B2(n2950), 
        .ZN(n15568) );
  MOAI22 U24482 ( .A1(n29196), .A2(n2951), .B1(ram[11328]), .B2(n2952), 
        .ZN(n15569) );
  MOAI22 U24483 ( .A1(n28961), .A2(n2951), .B1(ram[11329]), .B2(n2952), 
        .ZN(n15570) );
  MOAI22 U24484 ( .A1(n28726), .A2(n2951), .B1(ram[11330]), .B2(n2952), 
        .ZN(n15571) );
  MOAI22 U24485 ( .A1(n28491), .A2(n2951), .B1(ram[11331]), .B2(n2952), 
        .ZN(n15572) );
  MOAI22 U24486 ( .A1(n28256), .A2(n2951), .B1(ram[11332]), .B2(n2952), 
        .ZN(n15573) );
  MOAI22 U24487 ( .A1(n28021), .A2(n2951), .B1(ram[11333]), .B2(n2952), 
        .ZN(n15574) );
  MOAI22 U24488 ( .A1(n27786), .A2(n2951), .B1(ram[11334]), .B2(n2952), 
        .ZN(n15575) );
  MOAI22 U24489 ( .A1(n27551), .A2(n2951), .B1(ram[11335]), .B2(n2952), 
        .ZN(n15576) );
  MOAI22 U24490 ( .A1(n29197), .A2(n2953), .B1(ram[11336]), .B2(n2954), 
        .ZN(n15577) );
  MOAI22 U24491 ( .A1(n28962), .A2(n2953), .B1(ram[11337]), .B2(n2954), 
        .ZN(n15578) );
  MOAI22 U24492 ( .A1(n28727), .A2(n2953), .B1(ram[11338]), .B2(n2954), 
        .ZN(n15579) );
  MOAI22 U24493 ( .A1(n28492), .A2(n2953), .B1(ram[11339]), .B2(n2954), 
        .ZN(n15580) );
  MOAI22 U24494 ( .A1(n28257), .A2(n2953), .B1(ram[11340]), .B2(n2954), 
        .ZN(n15581) );
  MOAI22 U24495 ( .A1(n28022), .A2(n2953), .B1(ram[11341]), .B2(n2954), 
        .ZN(n15582) );
  MOAI22 U24496 ( .A1(n27787), .A2(n2953), .B1(ram[11342]), .B2(n2954), 
        .ZN(n15583) );
  MOAI22 U24497 ( .A1(n27552), .A2(n2953), .B1(ram[11343]), .B2(n2954), 
        .ZN(n15584) );
  MOAI22 U24498 ( .A1(n29197), .A2(n2955), .B1(ram[11344]), .B2(n2956), 
        .ZN(n15585) );
  MOAI22 U24499 ( .A1(n28962), .A2(n2955), .B1(ram[11345]), .B2(n2956), 
        .ZN(n15586) );
  MOAI22 U24500 ( .A1(n28727), .A2(n2955), .B1(ram[11346]), .B2(n2956), 
        .ZN(n15587) );
  MOAI22 U24501 ( .A1(n28492), .A2(n2955), .B1(ram[11347]), .B2(n2956), 
        .ZN(n15588) );
  MOAI22 U24502 ( .A1(n28257), .A2(n2955), .B1(ram[11348]), .B2(n2956), 
        .ZN(n15589) );
  MOAI22 U24503 ( .A1(n28022), .A2(n2955), .B1(ram[11349]), .B2(n2956), 
        .ZN(n15590) );
  MOAI22 U24504 ( .A1(n27787), .A2(n2955), .B1(ram[11350]), .B2(n2956), 
        .ZN(n15591) );
  MOAI22 U24505 ( .A1(n27552), .A2(n2955), .B1(ram[11351]), .B2(n2956), 
        .ZN(n15592) );
  MOAI22 U24506 ( .A1(n29197), .A2(n2957), .B1(ram[11352]), .B2(n2958), 
        .ZN(n15593) );
  MOAI22 U24507 ( .A1(n28962), .A2(n2957), .B1(ram[11353]), .B2(n2958), 
        .ZN(n15594) );
  MOAI22 U24508 ( .A1(n28727), .A2(n2957), .B1(ram[11354]), .B2(n2958), 
        .ZN(n15595) );
  MOAI22 U24509 ( .A1(n28492), .A2(n2957), .B1(ram[11355]), .B2(n2958), 
        .ZN(n15596) );
  MOAI22 U24510 ( .A1(n28257), .A2(n2957), .B1(ram[11356]), .B2(n2958), 
        .ZN(n15597) );
  MOAI22 U24511 ( .A1(n28022), .A2(n2957), .B1(ram[11357]), .B2(n2958), 
        .ZN(n15598) );
  MOAI22 U24512 ( .A1(n27787), .A2(n2957), .B1(ram[11358]), .B2(n2958), 
        .ZN(n15599) );
  MOAI22 U24513 ( .A1(n27552), .A2(n2957), .B1(ram[11359]), .B2(n2958), 
        .ZN(n15600) );
  MOAI22 U24514 ( .A1(n29197), .A2(n2959), .B1(ram[11360]), .B2(n2960), 
        .ZN(n15601) );
  MOAI22 U24515 ( .A1(n28962), .A2(n2959), .B1(ram[11361]), .B2(n2960), 
        .ZN(n15602) );
  MOAI22 U24516 ( .A1(n28727), .A2(n2959), .B1(ram[11362]), .B2(n2960), 
        .ZN(n15603) );
  MOAI22 U24517 ( .A1(n28492), .A2(n2959), .B1(ram[11363]), .B2(n2960), 
        .ZN(n15604) );
  MOAI22 U24518 ( .A1(n28257), .A2(n2959), .B1(ram[11364]), .B2(n2960), 
        .ZN(n15605) );
  MOAI22 U24519 ( .A1(n28022), .A2(n2959), .B1(ram[11365]), .B2(n2960), 
        .ZN(n15606) );
  MOAI22 U24520 ( .A1(n27787), .A2(n2959), .B1(ram[11366]), .B2(n2960), 
        .ZN(n15607) );
  MOAI22 U24521 ( .A1(n27552), .A2(n2959), .B1(ram[11367]), .B2(n2960), 
        .ZN(n15608) );
  MOAI22 U24522 ( .A1(n29197), .A2(n2961), .B1(ram[11368]), .B2(n2962), 
        .ZN(n15609) );
  MOAI22 U24523 ( .A1(n28962), .A2(n2961), .B1(ram[11369]), .B2(n2962), 
        .ZN(n15610) );
  MOAI22 U24524 ( .A1(n28727), .A2(n2961), .B1(ram[11370]), .B2(n2962), 
        .ZN(n15611) );
  MOAI22 U24525 ( .A1(n28492), .A2(n2961), .B1(ram[11371]), .B2(n2962), 
        .ZN(n15612) );
  MOAI22 U24526 ( .A1(n28257), .A2(n2961), .B1(ram[11372]), .B2(n2962), 
        .ZN(n15613) );
  MOAI22 U24527 ( .A1(n28022), .A2(n2961), .B1(ram[11373]), .B2(n2962), 
        .ZN(n15614) );
  MOAI22 U24528 ( .A1(n27787), .A2(n2961), .B1(ram[11374]), .B2(n2962), 
        .ZN(n15615) );
  MOAI22 U24529 ( .A1(n27552), .A2(n2961), .B1(ram[11375]), .B2(n2962), 
        .ZN(n15616) );
  MOAI22 U24530 ( .A1(n29197), .A2(n2963), .B1(ram[11376]), .B2(n2964), 
        .ZN(n15617) );
  MOAI22 U24531 ( .A1(n28962), .A2(n2963), .B1(ram[11377]), .B2(n2964), 
        .ZN(n15618) );
  MOAI22 U24532 ( .A1(n28727), .A2(n2963), .B1(ram[11378]), .B2(n2964), 
        .ZN(n15619) );
  MOAI22 U24533 ( .A1(n28492), .A2(n2963), .B1(ram[11379]), .B2(n2964), 
        .ZN(n15620) );
  MOAI22 U24534 ( .A1(n28257), .A2(n2963), .B1(ram[11380]), .B2(n2964), 
        .ZN(n15621) );
  MOAI22 U24535 ( .A1(n28022), .A2(n2963), .B1(ram[11381]), .B2(n2964), 
        .ZN(n15622) );
  MOAI22 U24536 ( .A1(n27787), .A2(n2963), .B1(ram[11382]), .B2(n2964), 
        .ZN(n15623) );
  MOAI22 U24537 ( .A1(n27552), .A2(n2963), .B1(ram[11383]), .B2(n2964), 
        .ZN(n15624) );
  MOAI22 U24538 ( .A1(n29197), .A2(n2965), .B1(ram[11384]), .B2(n2966), 
        .ZN(n15625) );
  MOAI22 U24539 ( .A1(n28962), .A2(n2965), .B1(ram[11385]), .B2(n2966), 
        .ZN(n15626) );
  MOAI22 U24540 ( .A1(n28727), .A2(n2965), .B1(ram[11386]), .B2(n2966), 
        .ZN(n15627) );
  MOAI22 U24541 ( .A1(n28492), .A2(n2965), .B1(ram[11387]), .B2(n2966), 
        .ZN(n15628) );
  MOAI22 U24542 ( .A1(n28257), .A2(n2965), .B1(ram[11388]), .B2(n2966), 
        .ZN(n15629) );
  MOAI22 U24543 ( .A1(n28022), .A2(n2965), .B1(ram[11389]), .B2(n2966), 
        .ZN(n15630) );
  MOAI22 U24544 ( .A1(n27787), .A2(n2965), .B1(ram[11390]), .B2(n2966), 
        .ZN(n15631) );
  MOAI22 U24545 ( .A1(n27552), .A2(n2965), .B1(ram[11391]), .B2(n2966), 
        .ZN(n15632) );
  MOAI22 U24546 ( .A1(n29197), .A2(n2967), .B1(ram[11392]), .B2(n2968), 
        .ZN(n15633) );
  MOAI22 U24547 ( .A1(n28962), .A2(n2967), .B1(ram[11393]), .B2(n2968), 
        .ZN(n15634) );
  MOAI22 U24548 ( .A1(n28727), .A2(n2967), .B1(ram[11394]), .B2(n2968), 
        .ZN(n15635) );
  MOAI22 U24549 ( .A1(n28492), .A2(n2967), .B1(ram[11395]), .B2(n2968), 
        .ZN(n15636) );
  MOAI22 U24550 ( .A1(n28257), .A2(n2967), .B1(ram[11396]), .B2(n2968), 
        .ZN(n15637) );
  MOAI22 U24551 ( .A1(n28022), .A2(n2967), .B1(ram[11397]), .B2(n2968), 
        .ZN(n15638) );
  MOAI22 U24552 ( .A1(n27787), .A2(n2967), .B1(ram[11398]), .B2(n2968), 
        .ZN(n15639) );
  MOAI22 U24553 ( .A1(n27552), .A2(n2967), .B1(ram[11399]), .B2(n2968), 
        .ZN(n15640) );
  MOAI22 U24554 ( .A1(n29197), .A2(n2969), .B1(ram[11400]), .B2(n2970), 
        .ZN(n15641) );
  MOAI22 U24555 ( .A1(n28962), .A2(n2969), .B1(ram[11401]), .B2(n2970), 
        .ZN(n15642) );
  MOAI22 U24556 ( .A1(n28727), .A2(n2969), .B1(ram[11402]), .B2(n2970), 
        .ZN(n15643) );
  MOAI22 U24557 ( .A1(n28492), .A2(n2969), .B1(ram[11403]), .B2(n2970), 
        .ZN(n15644) );
  MOAI22 U24558 ( .A1(n28257), .A2(n2969), .B1(ram[11404]), .B2(n2970), 
        .ZN(n15645) );
  MOAI22 U24559 ( .A1(n28022), .A2(n2969), .B1(ram[11405]), .B2(n2970), 
        .ZN(n15646) );
  MOAI22 U24560 ( .A1(n27787), .A2(n2969), .B1(ram[11406]), .B2(n2970), 
        .ZN(n15647) );
  MOAI22 U24561 ( .A1(n27552), .A2(n2969), .B1(ram[11407]), .B2(n2970), 
        .ZN(n15648) );
  MOAI22 U24562 ( .A1(n29197), .A2(n2971), .B1(ram[11408]), .B2(n2972), 
        .ZN(n15649) );
  MOAI22 U24563 ( .A1(n28962), .A2(n2971), .B1(ram[11409]), .B2(n2972), 
        .ZN(n15650) );
  MOAI22 U24564 ( .A1(n28727), .A2(n2971), .B1(ram[11410]), .B2(n2972), 
        .ZN(n15651) );
  MOAI22 U24565 ( .A1(n28492), .A2(n2971), .B1(ram[11411]), .B2(n2972), 
        .ZN(n15652) );
  MOAI22 U24566 ( .A1(n28257), .A2(n2971), .B1(ram[11412]), .B2(n2972), 
        .ZN(n15653) );
  MOAI22 U24567 ( .A1(n28022), .A2(n2971), .B1(ram[11413]), .B2(n2972), 
        .ZN(n15654) );
  MOAI22 U24568 ( .A1(n27787), .A2(n2971), .B1(ram[11414]), .B2(n2972), 
        .ZN(n15655) );
  MOAI22 U24569 ( .A1(n27552), .A2(n2971), .B1(ram[11415]), .B2(n2972), 
        .ZN(n15656) );
  MOAI22 U24570 ( .A1(n29197), .A2(n2973), .B1(ram[11416]), .B2(n2974), 
        .ZN(n15657) );
  MOAI22 U24571 ( .A1(n28962), .A2(n2973), .B1(ram[11417]), .B2(n2974), 
        .ZN(n15658) );
  MOAI22 U24572 ( .A1(n28727), .A2(n2973), .B1(ram[11418]), .B2(n2974), 
        .ZN(n15659) );
  MOAI22 U24573 ( .A1(n28492), .A2(n2973), .B1(ram[11419]), .B2(n2974), 
        .ZN(n15660) );
  MOAI22 U24574 ( .A1(n28257), .A2(n2973), .B1(ram[11420]), .B2(n2974), 
        .ZN(n15661) );
  MOAI22 U24575 ( .A1(n28022), .A2(n2973), .B1(ram[11421]), .B2(n2974), 
        .ZN(n15662) );
  MOAI22 U24576 ( .A1(n27787), .A2(n2973), .B1(ram[11422]), .B2(n2974), 
        .ZN(n15663) );
  MOAI22 U24577 ( .A1(n27552), .A2(n2973), .B1(ram[11423]), .B2(n2974), 
        .ZN(n15664) );
  MOAI22 U24578 ( .A1(n29197), .A2(n2975), .B1(ram[11424]), .B2(n2976), 
        .ZN(n15665) );
  MOAI22 U24579 ( .A1(n28962), .A2(n2975), .B1(ram[11425]), .B2(n2976), 
        .ZN(n15666) );
  MOAI22 U24580 ( .A1(n28727), .A2(n2975), .B1(ram[11426]), .B2(n2976), 
        .ZN(n15667) );
  MOAI22 U24581 ( .A1(n28492), .A2(n2975), .B1(ram[11427]), .B2(n2976), 
        .ZN(n15668) );
  MOAI22 U24582 ( .A1(n28257), .A2(n2975), .B1(ram[11428]), .B2(n2976), 
        .ZN(n15669) );
  MOAI22 U24583 ( .A1(n28022), .A2(n2975), .B1(ram[11429]), .B2(n2976), 
        .ZN(n15670) );
  MOAI22 U24584 ( .A1(n27787), .A2(n2975), .B1(ram[11430]), .B2(n2976), 
        .ZN(n15671) );
  MOAI22 U24585 ( .A1(n27552), .A2(n2975), .B1(ram[11431]), .B2(n2976), 
        .ZN(n15672) );
  MOAI22 U24586 ( .A1(n29197), .A2(n2977), .B1(ram[11432]), .B2(n2978), 
        .ZN(n15673) );
  MOAI22 U24587 ( .A1(n28962), .A2(n2977), .B1(ram[11433]), .B2(n2978), 
        .ZN(n15674) );
  MOAI22 U24588 ( .A1(n28727), .A2(n2977), .B1(ram[11434]), .B2(n2978), 
        .ZN(n15675) );
  MOAI22 U24589 ( .A1(n28492), .A2(n2977), .B1(ram[11435]), .B2(n2978), 
        .ZN(n15676) );
  MOAI22 U24590 ( .A1(n28257), .A2(n2977), .B1(ram[11436]), .B2(n2978), 
        .ZN(n15677) );
  MOAI22 U24591 ( .A1(n28022), .A2(n2977), .B1(ram[11437]), .B2(n2978), 
        .ZN(n15678) );
  MOAI22 U24592 ( .A1(n27787), .A2(n2977), .B1(ram[11438]), .B2(n2978), 
        .ZN(n15679) );
  MOAI22 U24593 ( .A1(n27552), .A2(n2977), .B1(ram[11439]), .B2(n2978), 
        .ZN(n15680) );
  MOAI22 U24594 ( .A1(n29198), .A2(n2979), .B1(ram[11440]), .B2(n2980), 
        .ZN(n15681) );
  MOAI22 U24595 ( .A1(n28963), .A2(n2979), .B1(ram[11441]), .B2(n2980), 
        .ZN(n15682) );
  MOAI22 U24596 ( .A1(n28728), .A2(n2979), .B1(ram[11442]), .B2(n2980), 
        .ZN(n15683) );
  MOAI22 U24597 ( .A1(n28493), .A2(n2979), .B1(ram[11443]), .B2(n2980), 
        .ZN(n15684) );
  MOAI22 U24598 ( .A1(n28258), .A2(n2979), .B1(ram[11444]), .B2(n2980), 
        .ZN(n15685) );
  MOAI22 U24599 ( .A1(n28023), .A2(n2979), .B1(ram[11445]), .B2(n2980), 
        .ZN(n15686) );
  MOAI22 U24600 ( .A1(n27788), .A2(n2979), .B1(ram[11446]), .B2(n2980), 
        .ZN(n15687) );
  MOAI22 U24601 ( .A1(n27553), .A2(n2979), .B1(ram[11447]), .B2(n2980), 
        .ZN(n15688) );
  MOAI22 U24602 ( .A1(n29198), .A2(n2981), .B1(ram[11448]), .B2(n2982), 
        .ZN(n15689) );
  MOAI22 U24603 ( .A1(n28963), .A2(n2981), .B1(ram[11449]), .B2(n2982), 
        .ZN(n15690) );
  MOAI22 U24604 ( .A1(n28728), .A2(n2981), .B1(ram[11450]), .B2(n2982), 
        .ZN(n15691) );
  MOAI22 U24605 ( .A1(n28493), .A2(n2981), .B1(ram[11451]), .B2(n2982), 
        .ZN(n15692) );
  MOAI22 U24606 ( .A1(n28258), .A2(n2981), .B1(ram[11452]), .B2(n2982), 
        .ZN(n15693) );
  MOAI22 U24607 ( .A1(n28023), .A2(n2981), .B1(ram[11453]), .B2(n2982), 
        .ZN(n15694) );
  MOAI22 U24608 ( .A1(n27788), .A2(n2981), .B1(ram[11454]), .B2(n2982), 
        .ZN(n15695) );
  MOAI22 U24609 ( .A1(n27553), .A2(n2981), .B1(ram[11455]), .B2(n2982), 
        .ZN(n15696) );
  MOAI22 U24610 ( .A1(n29198), .A2(n2983), .B1(ram[11456]), .B2(n2984), 
        .ZN(n15697) );
  MOAI22 U24611 ( .A1(n28963), .A2(n2983), .B1(ram[11457]), .B2(n2984), 
        .ZN(n15698) );
  MOAI22 U24612 ( .A1(n28728), .A2(n2983), .B1(ram[11458]), .B2(n2984), 
        .ZN(n15699) );
  MOAI22 U24613 ( .A1(n28493), .A2(n2983), .B1(ram[11459]), .B2(n2984), 
        .ZN(n15700) );
  MOAI22 U24614 ( .A1(n28258), .A2(n2983), .B1(ram[11460]), .B2(n2984), 
        .ZN(n15701) );
  MOAI22 U24615 ( .A1(n28023), .A2(n2983), .B1(ram[11461]), .B2(n2984), 
        .ZN(n15702) );
  MOAI22 U24616 ( .A1(n27788), .A2(n2983), .B1(ram[11462]), .B2(n2984), 
        .ZN(n15703) );
  MOAI22 U24617 ( .A1(n27553), .A2(n2983), .B1(ram[11463]), .B2(n2984), 
        .ZN(n15704) );
  MOAI22 U24618 ( .A1(n29198), .A2(n2985), .B1(ram[11464]), .B2(n2986), 
        .ZN(n15705) );
  MOAI22 U24619 ( .A1(n28963), .A2(n2985), .B1(ram[11465]), .B2(n2986), 
        .ZN(n15706) );
  MOAI22 U24620 ( .A1(n28728), .A2(n2985), .B1(ram[11466]), .B2(n2986), 
        .ZN(n15707) );
  MOAI22 U24621 ( .A1(n28493), .A2(n2985), .B1(ram[11467]), .B2(n2986), 
        .ZN(n15708) );
  MOAI22 U24622 ( .A1(n28258), .A2(n2985), .B1(ram[11468]), .B2(n2986), 
        .ZN(n15709) );
  MOAI22 U24623 ( .A1(n28023), .A2(n2985), .B1(ram[11469]), .B2(n2986), 
        .ZN(n15710) );
  MOAI22 U24624 ( .A1(n27788), .A2(n2985), .B1(ram[11470]), .B2(n2986), 
        .ZN(n15711) );
  MOAI22 U24625 ( .A1(n27553), .A2(n2985), .B1(ram[11471]), .B2(n2986), 
        .ZN(n15712) );
  MOAI22 U24626 ( .A1(n29198), .A2(n2987), .B1(ram[11472]), .B2(n2988), 
        .ZN(n15713) );
  MOAI22 U24627 ( .A1(n28963), .A2(n2987), .B1(ram[11473]), .B2(n2988), 
        .ZN(n15714) );
  MOAI22 U24628 ( .A1(n28728), .A2(n2987), .B1(ram[11474]), .B2(n2988), 
        .ZN(n15715) );
  MOAI22 U24629 ( .A1(n28493), .A2(n2987), .B1(ram[11475]), .B2(n2988), 
        .ZN(n15716) );
  MOAI22 U24630 ( .A1(n28258), .A2(n2987), .B1(ram[11476]), .B2(n2988), 
        .ZN(n15717) );
  MOAI22 U24631 ( .A1(n28023), .A2(n2987), .B1(ram[11477]), .B2(n2988), 
        .ZN(n15718) );
  MOAI22 U24632 ( .A1(n27788), .A2(n2987), .B1(ram[11478]), .B2(n2988), 
        .ZN(n15719) );
  MOAI22 U24633 ( .A1(n27553), .A2(n2987), .B1(ram[11479]), .B2(n2988), 
        .ZN(n15720) );
  MOAI22 U24634 ( .A1(n29198), .A2(n2989), .B1(ram[11480]), .B2(n2990), 
        .ZN(n15721) );
  MOAI22 U24635 ( .A1(n28963), .A2(n2989), .B1(ram[11481]), .B2(n2990), 
        .ZN(n15722) );
  MOAI22 U24636 ( .A1(n28728), .A2(n2989), .B1(ram[11482]), .B2(n2990), 
        .ZN(n15723) );
  MOAI22 U24637 ( .A1(n28493), .A2(n2989), .B1(ram[11483]), .B2(n2990), 
        .ZN(n15724) );
  MOAI22 U24638 ( .A1(n28258), .A2(n2989), .B1(ram[11484]), .B2(n2990), 
        .ZN(n15725) );
  MOAI22 U24639 ( .A1(n28023), .A2(n2989), .B1(ram[11485]), .B2(n2990), 
        .ZN(n15726) );
  MOAI22 U24640 ( .A1(n27788), .A2(n2989), .B1(ram[11486]), .B2(n2990), 
        .ZN(n15727) );
  MOAI22 U24641 ( .A1(n27553), .A2(n2989), .B1(ram[11487]), .B2(n2990), 
        .ZN(n15728) );
  MOAI22 U24642 ( .A1(n29198), .A2(n2991), .B1(ram[11488]), .B2(n2992), 
        .ZN(n15729) );
  MOAI22 U24643 ( .A1(n28963), .A2(n2991), .B1(ram[11489]), .B2(n2992), 
        .ZN(n15730) );
  MOAI22 U24644 ( .A1(n28728), .A2(n2991), .B1(ram[11490]), .B2(n2992), 
        .ZN(n15731) );
  MOAI22 U24645 ( .A1(n28493), .A2(n2991), .B1(ram[11491]), .B2(n2992), 
        .ZN(n15732) );
  MOAI22 U24646 ( .A1(n28258), .A2(n2991), .B1(ram[11492]), .B2(n2992), 
        .ZN(n15733) );
  MOAI22 U24647 ( .A1(n28023), .A2(n2991), .B1(ram[11493]), .B2(n2992), 
        .ZN(n15734) );
  MOAI22 U24648 ( .A1(n27788), .A2(n2991), .B1(ram[11494]), .B2(n2992), 
        .ZN(n15735) );
  MOAI22 U24649 ( .A1(n27553), .A2(n2991), .B1(ram[11495]), .B2(n2992), 
        .ZN(n15736) );
  MOAI22 U24650 ( .A1(n29198), .A2(n2993), .B1(ram[11496]), .B2(n2994), 
        .ZN(n15737) );
  MOAI22 U24651 ( .A1(n28963), .A2(n2993), .B1(ram[11497]), .B2(n2994), 
        .ZN(n15738) );
  MOAI22 U24652 ( .A1(n28728), .A2(n2993), .B1(ram[11498]), .B2(n2994), 
        .ZN(n15739) );
  MOAI22 U24653 ( .A1(n28493), .A2(n2993), .B1(ram[11499]), .B2(n2994), 
        .ZN(n15740) );
  MOAI22 U24654 ( .A1(n28258), .A2(n2993), .B1(ram[11500]), .B2(n2994), 
        .ZN(n15741) );
  MOAI22 U24655 ( .A1(n28023), .A2(n2993), .B1(ram[11501]), .B2(n2994), 
        .ZN(n15742) );
  MOAI22 U24656 ( .A1(n27788), .A2(n2993), .B1(ram[11502]), .B2(n2994), 
        .ZN(n15743) );
  MOAI22 U24657 ( .A1(n27553), .A2(n2993), .B1(ram[11503]), .B2(n2994), 
        .ZN(n15744) );
  MOAI22 U24658 ( .A1(n29198), .A2(n2995), .B1(ram[11504]), .B2(n2996), 
        .ZN(n15745) );
  MOAI22 U24659 ( .A1(n28963), .A2(n2995), .B1(ram[11505]), .B2(n2996), 
        .ZN(n15746) );
  MOAI22 U24660 ( .A1(n28728), .A2(n2995), .B1(ram[11506]), .B2(n2996), 
        .ZN(n15747) );
  MOAI22 U24661 ( .A1(n28493), .A2(n2995), .B1(ram[11507]), .B2(n2996), 
        .ZN(n15748) );
  MOAI22 U24662 ( .A1(n28258), .A2(n2995), .B1(ram[11508]), .B2(n2996), 
        .ZN(n15749) );
  MOAI22 U24663 ( .A1(n28023), .A2(n2995), .B1(ram[11509]), .B2(n2996), 
        .ZN(n15750) );
  MOAI22 U24664 ( .A1(n27788), .A2(n2995), .B1(ram[11510]), .B2(n2996), 
        .ZN(n15751) );
  MOAI22 U24665 ( .A1(n27553), .A2(n2995), .B1(ram[11511]), .B2(n2996), 
        .ZN(n15752) );
  MOAI22 U24666 ( .A1(n29198), .A2(n2997), .B1(ram[11512]), .B2(n2998), 
        .ZN(n15753) );
  MOAI22 U24667 ( .A1(n28963), .A2(n2997), .B1(ram[11513]), .B2(n2998), 
        .ZN(n15754) );
  MOAI22 U24668 ( .A1(n28728), .A2(n2997), .B1(ram[11514]), .B2(n2998), 
        .ZN(n15755) );
  MOAI22 U24669 ( .A1(n28493), .A2(n2997), .B1(ram[11515]), .B2(n2998), 
        .ZN(n15756) );
  MOAI22 U24670 ( .A1(n28258), .A2(n2997), .B1(ram[11516]), .B2(n2998), 
        .ZN(n15757) );
  MOAI22 U24671 ( .A1(n28023), .A2(n2997), .B1(ram[11517]), .B2(n2998), 
        .ZN(n15758) );
  MOAI22 U24672 ( .A1(n27788), .A2(n2997), .B1(ram[11518]), .B2(n2998), 
        .ZN(n15759) );
  MOAI22 U24673 ( .A1(n27553), .A2(n2997), .B1(ram[11519]), .B2(n2998), 
        .ZN(n15760) );
  MOAI22 U24674 ( .A1(n29198), .A2(n2999), .B1(ram[11520]), .B2(n3000), 
        .ZN(n15761) );
  MOAI22 U24675 ( .A1(n28963), .A2(n2999), .B1(ram[11521]), .B2(n3000), 
        .ZN(n15762) );
  MOAI22 U24676 ( .A1(n28728), .A2(n2999), .B1(ram[11522]), .B2(n3000), 
        .ZN(n15763) );
  MOAI22 U24677 ( .A1(n28493), .A2(n2999), .B1(ram[11523]), .B2(n3000), 
        .ZN(n15764) );
  MOAI22 U24678 ( .A1(n28258), .A2(n2999), .B1(ram[11524]), .B2(n3000), 
        .ZN(n15765) );
  MOAI22 U24679 ( .A1(n28023), .A2(n2999), .B1(ram[11525]), .B2(n3000), 
        .ZN(n15766) );
  MOAI22 U24680 ( .A1(n27788), .A2(n2999), .B1(ram[11526]), .B2(n3000), 
        .ZN(n15767) );
  MOAI22 U24681 ( .A1(n27553), .A2(n2999), .B1(ram[11527]), .B2(n3000), 
        .ZN(n15768) );
  MOAI22 U24682 ( .A1(n29198), .A2(n3001), .B1(ram[11528]), .B2(n3002), 
        .ZN(n15769) );
  MOAI22 U24683 ( .A1(n28963), .A2(n3001), .B1(ram[11529]), .B2(n3002), 
        .ZN(n15770) );
  MOAI22 U24684 ( .A1(n28728), .A2(n3001), .B1(ram[11530]), .B2(n3002), 
        .ZN(n15771) );
  MOAI22 U24685 ( .A1(n28493), .A2(n3001), .B1(ram[11531]), .B2(n3002), 
        .ZN(n15772) );
  MOAI22 U24686 ( .A1(n28258), .A2(n3001), .B1(ram[11532]), .B2(n3002), 
        .ZN(n15773) );
  MOAI22 U24687 ( .A1(n28023), .A2(n3001), .B1(ram[11533]), .B2(n3002), 
        .ZN(n15774) );
  MOAI22 U24688 ( .A1(n27788), .A2(n3001), .B1(ram[11534]), .B2(n3002), 
        .ZN(n15775) );
  MOAI22 U24689 ( .A1(n27553), .A2(n3001), .B1(ram[11535]), .B2(n3002), 
        .ZN(n15776) );
  MOAI22 U24690 ( .A1(n29198), .A2(n3003), .B1(ram[11536]), .B2(n3004), 
        .ZN(n15777) );
  MOAI22 U24691 ( .A1(n28963), .A2(n3003), .B1(ram[11537]), .B2(n3004), 
        .ZN(n15778) );
  MOAI22 U24692 ( .A1(n28728), .A2(n3003), .B1(ram[11538]), .B2(n3004), 
        .ZN(n15779) );
  MOAI22 U24693 ( .A1(n28493), .A2(n3003), .B1(ram[11539]), .B2(n3004), 
        .ZN(n15780) );
  MOAI22 U24694 ( .A1(n28258), .A2(n3003), .B1(ram[11540]), .B2(n3004), 
        .ZN(n15781) );
  MOAI22 U24695 ( .A1(n28023), .A2(n3003), .B1(ram[11541]), .B2(n3004), 
        .ZN(n15782) );
  MOAI22 U24696 ( .A1(n27788), .A2(n3003), .B1(ram[11542]), .B2(n3004), 
        .ZN(n15783) );
  MOAI22 U24697 ( .A1(n27553), .A2(n3003), .B1(ram[11543]), .B2(n3004), 
        .ZN(n15784) );
  MOAI22 U24698 ( .A1(n29199), .A2(n3005), .B1(ram[11544]), .B2(n3006), 
        .ZN(n15785) );
  MOAI22 U24699 ( .A1(n28964), .A2(n3005), .B1(ram[11545]), .B2(n3006), 
        .ZN(n15786) );
  MOAI22 U24700 ( .A1(n28729), .A2(n3005), .B1(ram[11546]), .B2(n3006), 
        .ZN(n15787) );
  MOAI22 U24701 ( .A1(n28494), .A2(n3005), .B1(ram[11547]), .B2(n3006), 
        .ZN(n15788) );
  MOAI22 U24702 ( .A1(n28259), .A2(n3005), .B1(ram[11548]), .B2(n3006), 
        .ZN(n15789) );
  MOAI22 U24703 ( .A1(n28024), .A2(n3005), .B1(ram[11549]), .B2(n3006), 
        .ZN(n15790) );
  MOAI22 U24704 ( .A1(n27789), .A2(n3005), .B1(ram[11550]), .B2(n3006), 
        .ZN(n15791) );
  MOAI22 U24705 ( .A1(n27554), .A2(n3005), .B1(ram[11551]), .B2(n3006), 
        .ZN(n15792) );
  MOAI22 U24706 ( .A1(n29199), .A2(n3007), .B1(ram[11552]), .B2(n3008), 
        .ZN(n15793) );
  MOAI22 U24707 ( .A1(n28964), .A2(n3007), .B1(ram[11553]), .B2(n3008), 
        .ZN(n15794) );
  MOAI22 U24708 ( .A1(n28729), .A2(n3007), .B1(ram[11554]), .B2(n3008), 
        .ZN(n15795) );
  MOAI22 U24709 ( .A1(n28494), .A2(n3007), .B1(ram[11555]), .B2(n3008), 
        .ZN(n15796) );
  MOAI22 U24710 ( .A1(n28259), .A2(n3007), .B1(ram[11556]), .B2(n3008), 
        .ZN(n15797) );
  MOAI22 U24711 ( .A1(n28024), .A2(n3007), .B1(ram[11557]), .B2(n3008), 
        .ZN(n15798) );
  MOAI22 U24712 ( .A1(n27789), .A2(n3007), .B1(ram[11558]), .B2(n3008), 
        .ZN(n15799) );
  MOAI22 U24713 ( .A1(n27554), .A2(n3007), .B1(ram[11559]), .B2(n3008), 
        .ZN(n15800) );
  MOAI22 U24714 ( .A1(n29199), .A2(n3009), .B1(ram[11560]), .B2(n3010), 
        .ZN(n15801) );
  MOAI22 U24715 ( .A1(n28964), .A2(n3009), .B1(ram[11561]), .B2(n3010), 
        .ZN(n15802) );
  MOAI22 U24716 ( .A1(n28729), .A2(n3009), .B1(ram[11562]), .B2(n3010), 
        .ZN(n15803) );
  MOAI22 U24717 ( .A1(n28494), .A2(n3009), .B1(ram[11563]), .B2(n3010), 
        .ZN(n15804) );
  MOAI22 U24718 ( .A1(n28259), .A2(n3009), .B1(ram[11564]), .B2(n3010), 
        .ZN(n15805) );
  MOAI22 U24719 ( .A1(n28024), .A2(n3009), .B1(ram[11565]), .B2(n3010), 
        .ZN(n15806) );
  MOAI22 U24720 ( .A1(n27789), .A2(n3009), .B1(ram[11566]), .B2(n3010), 
        .ZN(n15807) );
  MOAI22 U24721 ( .A1(n27554), .A2(n3009), .B1(ram[11567]), .B2(n3010), 
        .ZN(n15808) );
  MOAI22 U24722 ( .A1(n29199), .A2(n3011), .B1(ram[11568]), .B2(n3012), 
        .ZN(n15809) );
  MOAI22 U24723 ( .A1(n28964), .A2(n3011), .B1(ram[11569]), .B2(n3012), 
        .ZN(n15810) );
  MOAI22 U24724 ( .A1(n28729), .A2(n3011), .B1(ram[11570]), .B2(n3012), 
        .ZN(n15811) );
  MOAI22 U24725 ( .A1(n28494), .A2(n3011), .B1(ram[11571]), .B2(n3012), 
        .ZN(n15812) );
  MOAI22 U24726 ( .A1(n28259), .A2(n3011), .B1(ram[11572]), .B2(n3012), 
        .ZN(n15813) );
  MOAI22 U24727 ( .A1(n28024), .A2(n3011), .B1(ram[11573]), .B2(n3012), 
        .ZN(n15814) );
  MOAI22 U24728 ( .A1(n27789), .A2(n3011), .B1(ram[11574]), .B2(n3012), 
        .ZN(n15815) );
  MOAI22 U24729 ( .A1(n27554), .A2(n3011), .B1(ram[11575]), .B2(n3012), 
        .ZN(n15816) );
  MOAI22 U24730 ( .A1(n29199), .A2(n3013), .B1(ram[11576]), .B2(n3014), 
        .ZN(n15817) );
  MOAI22 U24731 ( .A1(n28964), .A2(n3013), .B1(ram[11577]), .B2(n3014), 
        .ZN(n15818) );
  MOAI22 U24732 ( .A1(n28729), .A2(n3013), .B1(ram[11578]), .B2(n3014), 
        .ZN(n15819) );
  MOAI22 U24733 ( .A1(n28494), .A2(n3013), .B1(ram[11579]), .B2(n3014), 
        .ZN(n15820) );
  MOAI22 U24734 ( .A1(n28259), .A2(n3013), .B1(ram[11580]), .B2(n3014), 
        .ZN(n15821) );
  MOAI22 U24735 ( .A1(n28024), .A2(n3013), .B1(ram[11581]), .B2(n3014), 
        .ZN(n15822) );
  MOAI22 U24736 ( .A1(n27789), .A2(n3013), .B1(ram[11582]), .B2(n3014), 
        .ZN(n15823) );
  MOAI22 U24737 ( .A1(n27554), .A2(n3013), .B1(ram[11583]), .B2(n3014), 
        .ZN(n15824) );
  MOAI22 U24738 ( .A1(n29199), .A2(n3015), .B1(ram[11584]), .B2(n3016), 
        .ZN(n15825) );
  MOAI22 U24739 ( .A1(n28964), .A2(n3015), .B1(ram[11585]), .B2(n3016), 
        .ZN(n15826) );
  MOAI22 U24740 ( .A1(n28729), .A2(n3015), .B1(ram[11586]), .B2(n3016), 
        .ZN(n15827) );
  MOAI22 U24741 ( .A1(n28494), .A2(n3015), .B1(ram[11587]), .B2(n3016), 
        .ZN(n15828) );
  MOAI22 U24742 ( .A1(n28259), .A2(n3015), .B1(ram[11588]), .B2(n3016), 
        .ZN(n15829) );
  MOAI22 U24743 ( .A1(n28024), .A2(n3015), .B1(ram[11589]), .B2(n3016), 
        .ZN(n15830) );
  MOAI22 U24744 ( .A1(n27789), .A2(n3015), .B1(ram[11590]), .B2(n3016), 
        .ZN(n15831) );
  MOAI22 U24745 ( .A1(n27554), .A2(n3015), .B1(ram[11591]), .B2(n3016), 
        .ZN(n15832) );
  MOAI22 U24746 ( .A1(n29199), .A2(n3017), .B1(ram[11592]), .B2(n3018), 
        .ZN(n15833) );
  MOAI22 U24747 ( .A1(n28964), .A2(n3017), .B1(ram[11593]), .B2(n3018), 
        .ZN(n15834) );
  MOAI22 U24748 ( .A1(n28729), .A2(n3017), .B1(ram[11594]), .B2(n3018), 
        .ZN(n15835) );
  MOAI22 U24749 ( .A1(n28494), .A2(n3017), .B1(ram[11595]), .B2(n3018), 
        .ZN(n15836) );
  MOAI22 U24750 ( .A1(n28259), .A2(n3017), .B1(ram[11596]), .B2(n3018), 
        .ZN(n15837) );
  MOAI22 U24751 ( .A1(n28024), .A2(n3017), .B1(ram[11597]), .B2(n3018), 
        .ZN(n15838) );
  MOAI22 U24752 ( .A1(n27789), .A2(n3017), .B1(ram[11598]), .B2(n3018), 
        .ZN(n15839) );
  MOAI22 U24753 ( .A1(n27554), .A2(n3017), .B1(ram[11599]), .B2(n3018), 
        .ZN(n15840) );
  MOAI22 U24754 ( .A1(n29199), .A2(n3019), .B1(ram[11600]), .B2(n3020), 
        .ZN(n15841) );
  MOAI22 U24755 ( .A1(n28964), .A2(n3019), .B1(ram[11601]), .B2(n3020), 
        .ZN(n15842) );
  MOAI22 U24756 ( .A1(n28729), .A2(n3019), .B1(ram[11602]), .B2(n3020), 
        .ZN(n15843) );
  MOAI22 U24757 ( .A1(n28494), .A2(n3019), .B1(ram[11603]), .B2(n3020), 
        .ZN(n15844) );
  MOAI22 U24758 ( .A1(n28259), .A2(n3019), .B1(ram[11604]), .B2(n3020), 
        .ZN(n15845) );
  MOAI22 U24759 ( .A1(n28024), .A2(n3019), .B1(ram[11605]), .B2(n3020), 
        .ZN(n15846) );
  MOAI22 U24760 ( .A1(n27789), .A2(n3019), .B1(ram[11606]), .B2(n3020), 
        .ZN(n15847) );
  MOAI22 U24761 ( .A1(n27554), .A2(n3019), .B1(ram[11607]), .B2(n3020), 
        .ZN(n15848) );
  MOAI22 U24762 ( .A1(n29199), .A2(n3021), .B1(ram[11608]), .B2(n3022), 
        .ZN(n15849) );
  MOAI22 U24763 ( .A1(n28964), .A2(n3021), .B1(ram[11609]), .B2(n3022), 
        .ZN(n15850) );
  MOAI22 U24764 ( .A1(n28729), .A2(n3021), .B1(ram[11610]), .B2(n3022), 
        .ZN(n15851) );
  MOAI22 U24765 ( .A1(n28494), .A2(n3021), .B1(ram[11611]), .B2(n3022), 
        .ZN(n15852) );
  MOAI22 U24766 ( .A1(n28259), .A2(n3021), .B1(ram[11612]), .B2(n3022), 
        .ZN(n15853) );
  MOAI22 U24767 ( .A1(n28024), .A2(n3021), .B1(ram[11613]), .B2(n3022), 
        .ZN(n15854) );
  MOAI22 U24768 ( .A1(n27789), .A2(n3021), .B1(ram[11614]), .B2(n3022), 
        .ZN(n15855) );
  MOAI22 U24769 ( .A1(n27554), .A2(n3021), .B1(ram[11615]), .B2(n3022), 
        .ZN(n15856) );
  MOAI22 U24770 ( .A1(n29199), .A2(n3023), .B1(ram[11616]), .B2(n3024), 
        .ZN(n15857) );
  MOAI22 U24771 ( .A1(n28964), .A2(n3023), .B1(ram[11617]), .B2(n3024), 
        .ZN(n15858) );
  MOAI22 U24772 ( .A1(n28729), .A2(n3023), .B1(ram[11618]), .B2(n3024), 
        .ZN(n15859) );
  MOAI22 U24773 ( .A1(n28494), .A2(n3023), .B1(ram[11619]), .B2(n3024), 
        .ZN(n15860) );
  MOAI22 U24774 ( .A1(n28259), .A2(n3023), .B1(ram[11620]), .B2(n3024), 
        .ZN(n15861) );
  MOAI22 U24775 ( .A1(n28024), .A2(n3023), .B1(ram[11621]), .B2(n3024), 
        .ZN(n15862) );
  MOAI22 U24776 ( .A1(n27789), .A2(n3023), .B1(ram[11622]), .B2(n3024), 
        .ZN(n15863) );
  MOAI22 U24777 ( .A1(n27554), .A2(n3023), .B1(ram[11623]), .B2(n3024), 
        .ZN(n15864) );
  MOAI22 U24778 ( .A1(n29199), .A2(n3025), .B1(ram[11624]), .B2(n3026), 
        .ZN(n15865) );
  MOAI22 U24779 ( .A1(n28964), .A2(n3025), .B1(ram[11625]), .B2(n3026), 
        .ZN(n15866) );
  MOAI22 U24780 ( .A1(n28729), .A2(n3025), .B1(ram[11626]), .B2(n3026), 
        .ZN(n15867) );
  MOAI22 U24781 ( .A1(n28494), .A2(n3025), .B1(ram[11627]), .B2(n3026), 
        .ZN(n15868) );
  MOAI22 U24782 ( .A1(n28259), .A2(n3025), .B1(ram[11628]), .B2(n3026), 
        .ZN(n15869) );
  MOAI22 U24783 ( .A1(n28024), .A2(n3025), .B1(ram[11629]), .B2(n3026), 
        .ZN(n15870) );
  MOAI22 U24784 ( .A1(n27789), .A2(n3025), .B1(ram[11630]), .B2(n3026), 
        .ZN(n15871) );
  MOAI22 U24785 ( .A1(n27554), .A2(n3025), .B1(ram[11631]), .B2(n3026), 
        .ZN(n15872) );
  MOAI22 U24786 ( .A1(n29199), .A2(n3027), .B1(ram[11632]), .B2(n3028), 
        .ZN(n15873) );
  MOAI22 U24787 ( .A1(n28964), .A2(n3027), .B1(ram[11633]), .B2(n3028), 
        .ZN(n15874) );
  MOAI22 U24788 ( .A1(n28729), .A2(n3027), .B1(ram[11634]), .B2(n3028), 
        .ZN(n15875) );
  MOAI22 U24789 ( .A1(n28494), .A2(n3027), .B1(ram[11635]), .B2(n3028), 
        .ZN(n15876) );
  MOAI22 U24790 ( .A1(n28259), .A2(n3027), .B1(ram[11636]), .B2(n3028), 
        .ZN(n15877) );
  MOAI22 U24791 ( .A1(n28024), .A2(n3027), .B1(ram[11637]), .B2(n3028), 
        .ZN(n15878) );
  MOAI22 U24792 ( .A1(n27789), .A2(n3027), .B1(ram[11638]), .B2(n3028), 
        .ZN(n15879) );
  MOAI22 U24793 ( .A1(n27554), .A2(n3027), .B1(ram[11639]), .B2(n3028), 
        .ZN(n15880) );
  MOAI22 U24794 ( .A1(n29199), .A2(n3029), .B1(ram[11640]), .B2(n3030), 
        .ZN(n15881) );
  MOAI22 U24795 ( .A1(n28964), .A2(n3029), .B1(ram[11641]), .B2(n3030), 
        .ZN(n15882) );
  MOAI22 U24796 ( .A1(n28729), .A2(n3029), .B1(ram[11642]), .B2(n3030), 
        .ZN(n15883) );
  MOAI22 U24797 ( .A1(n28494), .A2(n3029), .B1(ram[11643]), .B2(n3030), 
        .ZN(n15884) );
  MOAI22 U24798 ( .A1(n28259), .A2(n3029), .B1(ram[11644]), .B2(n3030), 
        .ZN(n15885) );
  MOAI22 U24799 ( .A1(n28024), .A2(n3029), .B1(ram[11645]), .B2(n3030), 
        .ZN(n15886) );
  MOAI22 U24800 ( .A1(n27789), .A2(n3029), .B1(ram[11646]), .B2(n3030), 
        .ZN(n15887) );
  MOAI22 U24801 ( .A1(n27554), .A2(n3029), .B1(ram[11647]), .B2(n3030), 
        .ZN(n15888) );
  MOAI22 U24802 ( .A1(n29200), .A2(n3031), .B1(ram[11648]), .B2(n3032), 
        .ZN(n15889) );
  MOAI22 U24803 ( .A1(n28965), .A2(n3031), .B1(ram[11649]), .B2(n3032), 
        .ZN(n15890) );
  MOAI22 U24804 ( .A1(n28730), .A2(n3031), .B1(ram[11650]), .B2(n3032), 
        .ZN(n15891) );
  MOAI22 U24805 ( .A1(n28495), .A2(n3031), .B1(ram[11651]), .B2(n3032), 
        .ZN(n15892) );
  MOAI22 U24806 ( .A1(n28260), .A2(n3031), .B1(ram[11652]), .B2(n3032), 
        .ZN(n15893) );
  MOAI22 U24807 ( .A1(n28025), .A2(n3031), .B1(ram[11653]), .B2(n3032), 
        .ZN(n15894) );
  MOAI22 U24808 ( .A1(n27790), .A2(n3031), .B1(ram[11654]), .B2(n3032), 
        .ZN(n15895) );
  MOAI22 U24809 ( .A1(n27555), .A2(n3031), .B1(ram[11655]), .B2(n3032), 
        .ZN(n15896) );
  MOAI22 U24810 ( .A1(n29200), .A2(n3033), .B1(ram[11656]), .B2(n3034), 
        .ZN(n15897) );
  MOAI22 U24811 ( .A1(n28965), .A2(n3033), .B1(ram[11657]), .B2(n3034), 
        .ZN(n15898) );
  MOAI22 U24812 ( .A1(n28730), .A2(n3033), .B1(ram[11658]), .B2(n3034), 
        .ZN(n15899) );
  MOAI22 U24813 ( .A1(n28495), .A2(n3033), .B1(ram[11659]), .B2(n3034), 
        .ZN(n15900) );
  MOAI22 U24814 ( .A1(n28260), .A2(n3033), .B1(ram[11660]), .B2(n3034), 
        .ZN(n15901) );
  MOAI22 U24815 ( .A1(n28025), .A2(n3033), .B1(ram[11661]), .B2(n3034), 
        .ZN(n15902) );
  MOAI22 U24816 ( .A1(n27790), .A2(n3033), .B1(ram[11662]), .B2(n3034), 
        .ZN(n15903) );
  MOAI22 U24817 ( .A1(n27555), .A2(n3033), .B1(ram[11663]), .B2(n3034), 
        .ZN(n15904) );
  MOAI22 U24818 ( .A1(n29200), .A2(n3035), .B1(ram[11664]), .B2(n3036), 
        .ZN(n15905) );
  MOAI22 U24819 ( .A1(n28965), .A2(n3035), .B1(ram[11665]), .B2(n3036), 
        .ZN(n15906) );
  MOAI22 U24820 ( .A1(n28730), .A2(n3035), .B1(ram[11666]), .B2(n3036), 
        .ZN(n15907) );
  MOAI22 U24821 ( .A1(n28495), .A2(n3035), .B1(ram[11667]), .B2(n3036), 
        .ZN(n15908) );
  MOAI22 U24822 ( .A1(n28260), .A2(n3035), .B1(ram[11668]), .B2(n3036), 
        .ZN(n15909) );
  MOAI22 U24823 ( .A1(n28025), .A2(n3035), .B1(ram[11669]), .B2(n3036), 
        .ZN(n15910) );
  MOAI22 U24824 ( .A1(n27790), .A2(n3035), .B1(ram[11670]), .B2(n3036), 
        .ZN(n15911) );
  MOAI22 U24825 ( .A1(n27555), .A2(n3035), .B1(ram[11671]), .B2(n3036), 
        .ZN(n15912) );
  MOAI22 U24826 ( .A1(n29200), .A2(n3037), .B1(ram[11672]), .B2(n3038), 
        .ZN(n15913) );
  MOAI22 U24827 ( .A1(n28965), .A2(n3037), .B1(ram[11673]), .B2(n3038), 
        .ZN(n15914) );
  MOAI22 U24828 ( .A1(n28730), .A2(n3037), .B1(ram[11674]), .B2(n3038), 
        .ZN(n15915) );
  MOAI22 U24829 ( .A1(n28495), .A2(n3037), .B1(ram[11675]), .B2(n3038), 
        .ZN(n15916) );
  MOAI22 U24830 ( .A1(n28260), .A2(n3037), .B1(ram[11676]), .B2(n3038), 
        .ZN(n15917) );
  MOAI22 U24831 ( .A1(n28025), .A2(n3037), .B1(ram[11677]), .B2(n3038), 
        .ZN(n15918) );
  MOAI22 U24832 ( .A1(n27790), .A2(n3037), .B1(ram[11678]), .B2(n3038), 
        .ZN(n15919) );
  MOAI22 U24833 ( .A1(n27555), .A2(n3037), .B1(ram[11679]), .B2(n3038), 
        .ZN(n15920) );
  MOAI22 U24834 ( .A1(n29200), .A2(n3039), .B1(ram[11680]), .B2(n3040), 
        .ZN(n15921) );
  MOAI22 U24835 ( .A1(n28965), .A2(n3039), .B1(ram[11681]), .B2(n3040), 
        .ZN(n15922) );
  MOAI22 U24836 ( .A1(n28730), .A2(n3039), .B1(ram[11682]), .B2(n3040), 
        .ZN(n15923) );
  MOAI22 U24837 ( .A1(n28495), .A2(n3039), .B1(ram[11683]), .B2(n3040), 
        .ZN(n15924) );
  MOAI22 U24838 ( .A1(n28260), .A2(n3039), .B1(ram[11684]), .B2(n3040), 
        .ZN(n15925) );
  MOAI22 U24839 ( .A1(n28025), .A2(n3039), .B1(ram[11685]), .B2(n3040), 
        .ZN(n15926) );
  MOAI22 U24840 ( .A1(n27790), .A2(n3039), .B1(ram[11686]), .B2(n3040), 
        .ZN(n15927) );
  MOAI22 U24841 ( .A1(n27555), .A2(n3039), .B1(ram[11687]), .B2(n3040), 
        .ZN(n15928) );
  MOAI22 U24842 ( .A1(n29200), .A2(n3041), .B1(ram[11688]), .B2(n3042), 
        .ZN(n15929) );
  MOAI22 U24843 ( .A1(n28965), .A2(n3041), .B1(ram[11689]), .B2(n3042), 
        .ZN(n15930) );
  MOAI22 U24844 ( .A1(n28730), .A2(n3041), .B1(ram[11690]), .B2(n3042), 
        .ZN(n15931) );
  MOAI22 U24845 ( .A1(n28495), .A2(n3041), .B1(ram[11691]), .B2(n3042), 
        .ZN(n15932) );
  MOAI22 U24846 ( .A1(n28260), .A2(n3041), .B1(ram[11692]), .B2(n3042), 
        .ZN(n15933) );
  MOAI22 U24847 ( .A1(n28025), .A2(n3041), .B1(ram[11693]), .B2(n3042), 
        .ZN(n15934) );
  MOAI22 U24848 ( .A1(n27790), .A2(n3041), .B1(ram[11694]), .B2(n3042), 
        .ZN(n15935) );
  MOAI22 U24849 ( .A1(n27555), .A2(n3041), .B1(ram[11695]), .B2(n3042), 
        .ZN(n15936) );
  MOAI22 U24850 ( .A1(n29200), .A2(n3043), .B1(ram[11696]), .B2(n3044), 
        .ZN(n15937) );
  MOAI22 U24851 ( .A1(n28965), .A2(n3043), .B1(ram[11697]), .B2(n3044), 
        .ZN(n15938) );
  MOAI22 U24852 ( .A1(n28730), .A2(n3043), .B1(ram[11698]), .B2(n3044), 
        .ZN(n15939) );
  MOAI22 U24853 ( .A1(n28495), .A2(n3043), .B1(ram[11699]), .B2(n3044), 
        .ZN(n15940) );
  MOAI22 U24854 ( .A1(n28260), .A2(n3043), .B1(ram[11700]), .B2(n3044), 
        .ZN(n15941) );
  MOAI22 U24855 ( .A1(n28025), .A2(n3043), .B1(ram[11701]), .B2(n3044), 
        .ZN(n15942) );
  MOAI22 U24856 ( .A1(n27790), .A2(n3043), .B1(ram[11702]), .B2(n3044), 
        .ZN(n15943) );
  MOAI22 U24857 ( .A1(n27555), .A2(n3043), .B1(ram[11703]), .B2(n3044), 
        .ZN(n15944) );
  MOAI22 U24858 ( .A1(n29200), .A2(n3045), .B1(ram[11704]), .B2(n3046), 
        .ZN(n15945) );
  MOAI22 U24859 ( .A1(n28965), .A2(n3045), .B1(ram[11705]), .B2(n3046), 
        .ZN(n15946) );
  MOAI22 U24860 ( .A1(n28730), .A2(n3045), .B1(ram[11706]), .B2(n3046), 
        .ZN(n15947) );
  MOAI22 U24861 ( .A1(n28495), .A2(n3045), .B1(ram[11707]), .B2(n3046), 
        .ZN(n15948) );
  MOAI22 U24862 ( .A1(n28260), .A2(n3045), .B1(ram[11708]), .B2(n3046), 
        .ZN(n15949) );
  MOAI22 U24863 ( .A1(n28025), .A2(n3045), .B1(ram[11709]), .B2(n3046), 
        .ZN(n15950) );
  MOAI22 U24864 ( .A1(n27790), .A2(n3045), .B1(ram[11710]), .B2(n3046), 
        .ZN(n15951) );
  MOAI22 U24865 ( .A1(n27555), .A2(n3045), .B1(ram[11711]), .B2(n3046), 
        .ZN(n15952) );
  MOAI22 U24866 ( .A1(n29200), .A2(n3047), .B1(ram[11712]), .B2(n3048), 
        .ZN(n15953) );
  MOAI22 U24867 ( .A1(n28965), .A2(n3047), .B1(ram[11713]), .B2(n3048), 
        .ZN(n15954) );
  MOAI22 U24868 ( .A1(n28730), .A2(n3047), .B1(ram[11714]), .B2(n3048), 
        .ZN(n15955) );
  MOAI22 U24869 ( .A1(n28495), .A2(n3047), .B1(ram[11715]), .B2(n3048), 
        .ZN(n15956) );
  MOAI22 U24870 ( .A1(n28260), .A2(n3047), .B1(ram[11716]), .B2(n3048), 
        .ZN(n15957) );
  MOAI22 U24871 ( .A1(n28025), .A2(n3047), .B1(ram[11717]), .B2(n3048), 
        .ZN(n15958) );
  MOAI22 U24872 ( .A1(n27790), .A2(n3047), .B1(ram[11718]), .B2(n3048), 
        .ZN(n15959) );
  MOAI22 U24873 ( .A1(n27555), .A2(n3047), .B1(ram[11719]), .B2(n3048), 
        .ZN(n15960) );
  MOAI22 U24874 ( .A1(n29200), .A2(n3049), .B1(ram[11720]), .B2(n3050), 
        .ZN(n15961) );
  MOAI22 U24875 ( .A1(n28965), .A2(n3049), .B1(ram[11721]), .B2(n3050), 
        .ZN(n15962) );
  MOAI22 U24876 ( .A1(n28730), .A2(n3049), .B1(ram[11722]), .B2(n3050), 
        .ZN(n15963) );
  MOAI22 U24877 ( .A1(n28495), .A2(n3049), .B1(ram[11723]), .B2(n3050), 
        .ZN(n15964) );
  MOAI22 U24878 ( .A1(n28260), .A2(n3049), .B1(ram[11724]), .B2(n3050), 
        .ZN(n15965) );
  MOAI22 U24879 ( .A1(n28025), .A2(n3049), .B1(ram[11725]), .B2(n3050), 
        .ZN(n15966) );
  MOAI22 U24880 ( .A1(n27790), .A2(n3049), .B1(ram[11726]), .B2(n3050), 
        .ZN(n15967) );
  MOAI22 U24881 ( .A1(n27555), .A2(n3049), .B1(ram[11727]), .B2(n3050), 
        .ZN(n15968) );
  MOAI22 U24882 ( .A1(n29200), .A2(n3051), .B1(ram[11728]), .B2(n3052), 
        .ZN(n15969) );
  MOAI22 U24883 ( .A1(n28965), .A2(n3051), .B1(ram[11729]), .B2(n3052), 
        .ZN(n15970) );
  MOAI22 U24884 ( .A1(n28730), .A2(n3051), .B1(ram[11730]), .B2(n3052), 
        .ZN(n15971) );
  MOAI22 U24885 ( .A1(n28495), .A2(n3051), .B1(ram[11731]), .B2(n3052), 
        .ZN(n15972) );
  MOAI22 U24886 ( .A1(n28260), .A2(n3051), .B1(ram[11732]), .B2(n3052), 
        .ZN(n15973) );
  MOAI22 U24887 ( .A1(n28025), .A2(n3051), .B1(ram[11733]), .B2(n3052), 
        .ZN(n15974) );
  MOAI22 U24888 ( .A1(n27790), .A2(n3051), .B1(ram[11734]), .B2(n3052), 
        .ZN(n15975) );
  MOAI22 U24889 ( .A1(n27555), .A2(n3051), .B1(ram[11735]), .B2(n3052), 
        .ZN(n15976) );
  MOAI22 U24890 ( .A1(n29200), .A2(n3053), .B1(ram[11736]), .B2(n3054), 
        .ZN(n15977) );
  MOAI22 U24891 ( .A1(n28965), .A2(n3053), .B1(ram[11737]), .B2(n3054), 
        .ZN(n15978) );
  MOAI22 U24892 ( .A1(n28730), .A2(n3053), .B1(ram[11738]), .B2(n3054), 
        .ZN(n15979) );
  MOAI22 U24893 ( .A1(n28495), .A2(n3053), .B1(ram[11739]), .B2(n3054), 
        .ZN(n15980) );
  MOAI22 U24894 ( .A1(n28260), .A2(n3053), .B1(ram[11740]), .B2(n3054), 
        .ZN(n15981) );
  MOAI22 U24895 ( .A1(n28025), .A2(n3053), .B1(ram[11741]), .B2(n3054), 
        .ZN(n15982) );
  MOAI22 U24896 ( .A1(n27790), .A2(n3053), .B1(ram[11742]), .B2(n3054), 
        .ZN(n15983) );
  MOAI22 U24897 ( .A1(n27555), .A2(n3053), .B1(ram[11743]), .B2(n3054), 
        .ZN(n15984) );
  MOAI22 U24898 ( .A1(n29200), .A2(n3055), .B1(ram[11744]), .B2(n3056), 
        .ZN(n15985) );
  MOAI22 U24899 ( .A1(n28965), .A2(n3055), .B1(ram[11745]), .B2(n3056), 
        .ZN(n15986) );
  MOAI22 U24900 ( .A1(n28730), .A2(n3055), .B1(ram[11746]), .B2(n3056), 
        .ZN(n15987) );
  MOAI22 U24901 ( .A1(n28495), .A2(n3055), .B1(ram[11747]), .B2(n3056), 
        .ZN(n15988) );
  MOAI22 U24902 ( .A1(n28260), .A2(n3055), .B1(ram[11748]), .B2(n3056), 
        .ZN(n15989) );
  MOAI22 U24903 ( .A1(n28025), .A2(n3055), .B1(ram[11749]), .B2(n3056), 
        .ZN(n15990) );
  MOAI22 U24904 ( .A1(n27790), .A2(n3055), .B1(ram[11750]), .B2(n3056), 
        .ZN(n15991) );
  MOAI22 U24905 ( .A1(n27555), .A2(n3055), .B1(ram[11751]), .B2(n3056), 
        .ZN(n15992) );
  MOAI22 U24906 ( .A1(n29201), .A2(n3057), .B1(ram[11752]), .B2(n3058), 
        .ZN(n15993) );
  MOAI22 U24907 ( .A1(n28966), .A2(n3057), .B1(ram[11753]), .B2(n3058), 
        .ZN(n15994) );
  MOAI22 U24908 ( .A1(n28731), .A2(n3057), .B1(ram[11754]), .B2(n3058), 
        .ZN(n15995) );
  MOAI22 U24909 ( .A1(n28496), .A2(n3057), .B1(ram[11755]), .B2(n3058), 
        .ZN(n15996) );
  MOAI22 U24910 ( .A1(n28261), .A2(n3057), .B1(ram[11756]), .B2(n3058), 
        .ZN(n15997) );
  MOAI22 U24911 ( .A1(n28026), .A2(n3057), .B1(ram[11757]), .B2(n3058), 
        .ZN(n15998) );
  MOAI22 U24912 ( .A1(n27791), .A2(n3057), .B1(ram[11758]), .B2(n3058), 
        .ZN(n15999) );
  MOAI22 U24913 ( .A1(n27556), .A2(n3057), .B1(ram[11759]), .B2(n3058), 
        .ZN(n16000) );
  MOAI22 U24914 ( .A1(n29201), .A2(n3059), .B1(ram[11760]), .B2(n3060), 
        .ZN(n16001) );
  MOAI22 U24915 ( .A1(n28966), .A2(n3059), .B1(ram[11761]), .B2(n3060), 
        .ZN(n16002) );
  MOAI22 U24916 ( .A1(n28731), .A2(n3059), .B1(ram[11762]), .B2(n3060), 
        .ZN(n16003) );
  MOAI22 U24917 ( .A1(n28496), .A2(n3059), .B1(ram[11763]), .B2(n3060), 
        .ZN(n16004) );
  MOAI22 U24918 ( .A1(n28261), .A2(n3059), .B1(ram[11764]), .B2(n3060), 
        .ZN(n16005) );
  MOAI22 U24919 ( .A1(n28026), .A2(n3059), .B1(ram[11765]), .B2(n3060), 
        .ZN(n16006) );
  MOAI22 U24920 ( .A1(n27791), .A2(n3059), .B1(ram[11766]), .B2(n3060), 
        .ZN(n16007) );
  MOAI22 U24921 ( .A1(n27556), .A2(n3059), .B1(ram[11767]), .B2(n3060), 
        .ZN(n16008) );
  MOAI22 U24922 ( .A1(n29201), .A2(n3061), .B1(ram[11768]), .B2(n3062), 
        .ZN(n16009) );
  MOAI22 U24923 ( .A1(n28966), .A2(n3061), .B1(ram[11769]), .B2(n3062), 
        .ZN(n16010) );
  MOAI22 U24924 ( .A1(n28731), .A2(n3061), .B1(ram[11770]), .B2(n3062), 
        .ZN(n16011) );
  MOAI22 U24925 ( .A1(n28496), .A2(n3061), .B1(ram[11771]), .B2(n3062), 
        .ZN(n16012) );
  MOAI22 U24926 ( .A1(n28261), .A2(n3061), .B1(ram[11772]), .B2(n3062), 
        .ZN(n16013) );
  MOAI22 U24927 ( .A1(n28026), .A2(n3061), .B1(ram[11773]), .B2(n3062), 
        .ZN(n16014) );
  MOAI22 U24928 ( .A1(n27791), .A2(n3061), .B1(ram[11774]), .B2(n3062), 
        .ZN(n16015) );
  MOAI22 U24929 ( .A1(n27556), .A2(n3061), .B1(ram[11775]), .B2(n3062), 
        .ZN(n16016) );
  MOAI22 U24930 ( .A1(n29201), .A2(n3063), .B1(ram[11776]), .B2(n3064), 
        .ZN(n16017) );
  MOAI22 U24931 ( .A1(n28966), .A2(n3063), .B1(ram[11777]), .B2(n3064), 
        .ZN(n16018) );
  MOAI22 U24932 ( .A1(n28731), .A2(n3063), .B1(ram[11778]), .B2(n3064), 
        .ZN(n16019) );
  MOAI22 U24933 ( .A1(n28496), .A2(n3063), .B1(ram[11779]), .B2(n3064), 
        .ZN(n16020) );
  MOAI22 U24934 ( .A1(n28261), .A2(n3063), .B1(ram[11780]), .B2(n3064), 
        .ZN(n16021) );
  MOAI22 U24935 ( .A1(n28026), .A2(n3063), .B1(ram[11781]), .B2(n3064), 
        .ZN(n16022) );
  MOAI22 U24936 ( .A1(n27791), .A2(n3063), .B1(ram[11782]), .B2(n3064), 
        .ZN(n16023) );
  MOAI22 U24937 ( .A1(n27556), .A2(n3063), .B1(ram[11783]), .B2(n3064), 
        .ZN(n16024) );
  MOAI22 U24938 ( .A1(n29201), .A2(n3066), .B1(ram[11784]), .B2(n3067), 
        .ZN(n16025) );
  MOAI22 U24939 ( .A1(n28966), .A2(n3066), .B1(ram[11785]), .B2(n3067), 
        .ZN(n16026) );
  MOAI22 U24940 ( .A1(n28731), .A2(n3066), .B1(ram[11786]), .B2(n3067), 
        .ZN(n16027) );
  MOAI22 U24941 ( .A1(n28496), .A2(n3066), .B1(ram[11787]), .B2(n3067), 
        .ZN(n16028) );
  MOAI22 U24942 ( .A1(n28261), .A2(n3066), .B1(ram[11788]), .B2(n3067), 
        .ZN(n16029) );
  MOAI22 U24943 ( .A1(n28026), .A2(n3066), .B1(ram[11789]), .B2(n3067), 
        .ZN(n16030) );
  MOAI22 U24944 ( .A1(n27791), .A2(n3066), .B1(ram[11790]), .B2(n3067), 
        .ZN(n16031) );
  MOAI22 U24945 ( .A1(n27556), .A2(n3066), .B1(ram[11791]), .B2(n3067), 
        .ZN(n16032) );
  MOAI22 U24946 ( .A1(n29201), .A2(n3068), .B1(ram[11792]), .B2(n3069), 
        .ZN(n16033) );
  MOAI22 U24947 ( .A1(n28966), .A2(n3068), .B1(ram[11793]), .B2(n3069), 
        .ZN(n16034) );
  MOAI22 U24948 ( .A1(n28731), .A2(n3068), .B1(ram[11794]), .B2(n3069), 
        .ZN(n16035) );
  MOAI22 U24949 ( .A1(n28496), .A2(n3068), .B1(ram[11795]), .B2(n3069), 
        .ZN(n16036) );
  MOAI22 U24950 ( .A1(n28261), .A2(n3068), .B1(ram[11796]), .B2(n3069), 
        .ZN(n16037) );
  MOAI22 U24951 ( .A1(n28026), .A2(n3068), .B1(ram[11797]), .B2(n3069), 
        .ZN(n16038) );
  MOAI22 U24952 ( .A1(n27791), .A2(n3068), .B1(ram[11798]), .B2(n3069), 
        .ZN(n16039) );
  MOAI22 U24953 ( .A1(n27556), .A2(n3068), .B1(ram[11799]), .B2(n3069), 
        .ZN(n16040) );
  MOAI22 U24954 ( .A1(n29201), .A2(n3070), .B1(ram[11800]), .B2(n3071), 
        .ZN(n16041) );
  MOAI22 U24955 ( .A1(n28966), .A2(n3070), .B1(ram[11801]), .B2(n3071), 
        .ZN(n16042) );
  MOAI22 U24956 ( .A1(n28731), .A2(n3070), .B1(ram[11802]), .B2(n3071), 
        .ZN(n16043) );
  MOAI22 U24957 ( .A1(n28496), .A2(n3070), .B1(ram[11803]), .B2(n3071), 
        .ZN(n16044) );
  MOAI22 U24958 ( .A1(n28261), .A2(n3070), .B1(ram[11804]), .B2(n3071), 
        .ZN(n16045) );
  MOAI22 U24959 ( .A1(n28026), .A2(n3070), .B1(ram[11805]), .B2(n3071), 
        .ZN(n16046) );
  MOAI22 U24960 ( .A1(n27791), .A2(n3070), .B1(ram[11806]), .B2(n3071), 
        .ZN(n16047) );
  MOAI22 U24961 ( .A1(n27556), .A2(n3070), .B1(ram[11807]), .B2(n3071), 
        .ZN(n16048) );
  MOAI22 U24962 ( .A1(n29201), .A2(n3072), .B1(ram[11808]), .B2(n3073), 
        .ZN(n16049) );
  MOAI22 U24963 ( .A1(n28966), .A2(n3072), .B1(ram[11809]), .B2(n3073), 
        .ZN(n16050) );
  MOAI22 U24964 ( .A1(n28731), .A2(n3072), .B1(ram[11810]), .B2(n3073), 
        .ZN(n16051) );
  MOAI22 U24965 ( .A1(n28496), .A2(n3072), .B1(ram[11811]), .B2(n3073), 
        .ZN(n16052) );
  MOAI22 U24966 ( .A1(n28261), .A2(n3072), .B1(ram[11812]), .B2(n3073), 
        .ZN(n16053) );
  MOAI22 U24967 ( .A1(n28026), .A2(n3072), .B1(ram[11813]), .B2(n3073), 
        .ZN(n16054) );
  MOAI22 U24968 ( .A1(n27791), .A2(n3072), .B1(ram[11814]), .B2(n3073), 
        .ZN(n16055) );
  MOAI22 U24969 ( .A1(n27556), .A2(n3072), .B1(ram[11815]), .B2(n3073), 
        .ZN(n16056) );
  MOAI22 U24970 ( .A1(n29201), .A2(n3074), .B1(ram[11816]), .B2(n3075), 
        .ZN(n16057) );
  MOAI22 U24971 ( .A1(n28966), .A2(n3074), .B1(ram[11817]), .B2(n3075), 
        .ZN(n16058) );
  MOAI22 U24972 ( .A1(n28731), .A2(n3074), .B1(ram[11818]), .B2(n3075), 
        .ZN(n16059) );
  MOAI22 U24973 ( .A1(n28496), .A2(n3074), .B1(ram[11819]), .B2(n3075), 
        .ZN(n16060) );
  MOAI22 U24974 ( .A1(n28261), .A2(n3074), .B1(ram[11820]), .B2(n3075), 
        .ZN(n16061) );
  MOAI22 U24975 ( .A1(n28026), .A2(n3074), .B1(ram[11821]), .B2(n3075), 
        .ZN(n16062) );
  MOAI22 U24976 ( .A1(n27791), .A2(n3074), .B1(ram[11822]), .B2(n3075), 
        .ZN(n16063) );
  MOAI22 U24977 ( .A1(n27556), .A2(n3074), .B1(ram[11823]), .B2(n3075), 
        .ZN(n16064) );
  MOAI22 U24978 ( .A1(n29201), .A2(n3076), .B1(ram[11824]), .B2(n3077), 
        .ZN(n16065) );
  MOAI22 U24979 ( .A1(n28966), .A2(n3076), .B1(ram[11825]), .B2(n3077), 
        .ZN(n16066) );
  MOAI22 U24980 ( .A1(n28731), .A2(n3076), .B1(ram[11826]), .B2(n3077), 
        .ZN(n16067) );
  MOAI22 U24981 ( .A1(n28496), .A2(n3076), .B1(ram[11827]), .B2(n3077), 
        .ZN(n16068) );
  MOAI22 U24982 ( .A1(n28261), .A2(n3076), .B1(ram[11828]), .B2(n3077), 
        .ZN(n16069) );
  MOAI22 U24983 ( .A1(n28026), .A2(n3076), .B1(ram[11829]), .B2(n3077), 
        .ZN(n16070) );
  MOAI22 U24984 ( .A1(n27791), .A2(n3076), .B1(ram[11830]), .B2(n3077), 
        .ZN(n16071) );
  MOAI22 U24985 ( .A1(n27556), .A2(n3076), .B1(ram[11831]), .B2(n3077), 
        .ZN(n16072) );
  MOAI22 U24986 ( .A1(n29201), .A2(n3078), .B1(ram[11832]), .B2(n3079), 
        .ZN(n16073) );
  MOAI22 U24987 ( .A1(n28966), .A2(n3078), .B1(ram[11833]), .B2(n3079), 
        .ZN(n16074) );
  MOAI22 U24988 ( .A1(n28731), .A2(n3078), .B1(ram[11834]), .B2(n3079), 
        .ZN(n16075) );
  MOAI22 U24989 ( .A1(n28496), .A2(n3078), .B1(ram[11835]), .B2(n3079), 
        .ZN(n16076) );
  MOAI22 U24990 ( .A1(n28261), .A2(n3078), .B1(ram[11836]), .B2(n3079), 
        .ZN(n16077) );
  MOAI22 U24991 ( .A1(n28026), .A2(n3078), .B1(ram[11837]), .B2(n3079), 
        .ZN(n16078) );
  MOAI22 U24992 ( .A1(n27791), .A2(n3078), .B1(ram[11838]), .B2(n3079), 
        .ZN(n16079) );
  MOAI22 U24993 ( .A1(n27556), .A2(n3078), .B1(ram[11839]), .B2(n3079), 
        .ZN(n16080) );
  MOAI22 U24994 ( .A1(n29201), .A2(n3080), .B1(ram[11840]), .B2(n3081), 
        .ZN(n16081) );
  MOAI22 U24995 ( .A1(n28966), .A2(n3080), .B1(ram[11841]), .B2(n3081), 
        .ZN(n16082) );
  MOAI22 U24996 ( .A1(n28731), .A2(n3080), .B1(ram[11842]), .B2(n3081), 
        .ZN(n16083) );
  MOAI22 U24997 ( .A1(n28496), .A2(n3080), .B1(ram[11843]), .B2(n3081), 
        .ZN(n16084) );
  MOAI22 U24998 ( .A1(n28261), .A2(n3080), .B1(ram[11844]), .B2(n3081), 
        .ZN(n16085) );
  MOAI22 U24999 ( .A1(n28026), .A2(n3080), .B1(ram[11845]), .B2(n3081), 
        .ZN(n16086) );
  MOAI22 U25000 ( .A1(n27791), .A2(n3080), .B1(ram[11846]), .B2(n3081), 
        .ZN(n16087) );
  MOAI22 U25001 ( .A1(n27556), .A2(n3080), .B1(ram[11847]), .B2(n3081), 
        .ZN(n16088) );
  MOAI22 U25002 ( .A1(n29201), .A2(n3082), .B1(ram[11848]), .B2(n3083), 
        .ZN(n16089) );
  MOAI22 U25003 ( .A1(n28966), .A2(n3082), .B1(ram[11849]), .B2(n3083), 
        .ZN(n16090) );
  MOAI22 U25004 ( .A1(n28731), .A2(n3082), .B1(ram[11850]), .B2(n3083), 
        .ZN(n16091) );
  MOAI22 U25005 ( .A1(n28496), .A2(n3082), .B1(ram[11851]), .B2(n3083), 
        .ZN(n16092) );
  MOAI22 U25006 ( .A1(n28261), .A2(n3082), .B1(ram[11852]), .B2(n3083), 
        .ZN(n16093) );
  MOAI22 U25007 ( .A1(n28026), .A2(n3082), .B1(ram[11853]), .B2(n3083), 
        .ZN(n16094) );
  MOAI22 U25008 ( .A1(n27791), .A2(n3082), .B1(ram[11854]), .B2(n3083), 
        .ZN(n16095) );
  MOAI22 U25009 ( .A1(n27556), .A2(n3082), .B1(ram[11855]), .B2(n3083), 
        .ZN(n16096) );
  MOAI22 U25010 ( .A1(n29202), .A2(n3084), .B1(ram[11856]), .B2(n3085), 
        .ZN(n16097) );
  MOAI22 U25011 ( .A1(n28967), .A2(n3084), .B1(ram[11857]), .B2(n3085), 
        .ZN(n16098) );
  MOAI22 U25012 ( .A1(n28732), .A2(n3084), .B1(ram[11858]), .B2(n3085), 
        .ZN(n16099) );
  MOAI22 U25013 ( .A1(n28497), .A2(n3084), .B1(ram[11859]), .B2(n3085), 
        .ZN(n16100) );
  MOAI22 U25014 ( .A1(n28262), .A2(n3084), .B1(ram[11860]), .B2(n3085), 
        .ZN(n16101) );
  MOAI22 U25015 ( .A1(n28027), .A2(n3084), .B1(ram[11861]), .B2(n3085), 
        .ZN(n16102) );
  MOAI22 U25016 ( .A1(n27792), .A2(n3084), .B1(ram[11862]), .B2(n3085), 
        .ZN(n16103) );
  MOAI22 U25017 ( .A1(n27557), .A2(n3084), .B1(ram[11863]), .B2(n3085), 
        .ZN(n16104) );
  MOAI22 U25018 ( .A1(n29202), .A2(n3086), .B1(ram[11864]), .B2(n3087), 
        .ZN(n16105) );
  MOAI22 U25019 ( .A1(n28967), .A2(n3086), .B1(ram[11865]), .B2(n3087), 
        .ZN(n16106) );
  MOAI22 U25020 ( .A1(n28732), .A2(n3086), .B1(ram[11866]), .B2(n3087), 
        .ZN(n16107) );
  MOAI22 U25021 ( .A1(n28497), .A2(n3086), .B1(ram[11867]), .B2(n3087), 
        .ZN(n16108) );
  MOAI22 U25022 ( .A1(n28262), .A2(n3086), .B1(ram[11868]), .B2(n3087), 
        .ZN(n16109) );
  MOAI22 U25023 ( .A1(n28027), .A2(n3086), .B1(ram[11869]), .B2(n3087), 
        .ZN(n16110) );
  MOAI22 U25024 ( .A1(n27792), .A2(n3086), .B1(ram[11870]), .B2(n3087), 
        .ZN(n16111) );
  MOAI22 U25025 ( .A1(n27557), .A2(n3086), .B1(ram[11871]), .B2(n3087), 
        .ZN(n16112) );
  MOAI22 U25026 ( .A1(n29202), .A2(n3088), .B1(ram[11872]), .B2(n3089), 
        .ZN(n16113) );
  MOAI22 U25027 ( .A1(n28967), .A2(n3088), .B1(ram[11873]), .B2(n3089), 
        .ZN(n16114) );
  MOAI22 U25028 ( .A1(n28732), .A2(n3088), .B1(ram[11874]), .B2(n3089), 
        .ZN(n16115) );
  MOAI22 U25029 ( .A1(n28497), .A2(n3088), .B1(ram[11875]), .B2(n3089), 
        .ZN(n16116) );
  MOAI22 U25030 ( .A1(n28262), .A2(n3088), .B1(ram[11876]), .B2(n3089), 
        .ZN(n16117) );
  MOAI22 U25031 ( .A1(n28027), .A2(n3088), .B1(ram[11877]), .B2(n3089), 
        .ZN(n16118) );
  MOAI22 U25032 ( .A1(n27792), .A2(n3088), .B1(ram[11878]), .B2(n3089), 
        .ZN(n16119) );
  MOAI22 U25033 ( .A1(n27557), .A2(n3088), .B1(ram[11879]), .B2(n3089), 
        .ZN(n16120) );
  MOAI22 U25034 ( .A1(n29202), .A2(n3090), .B1(ram[11880]), .B2(n3091), 
        .ZN(n16121) );
  MOAI22 U25035 ( .A1(n28967), .A2(n3090), .B1(ram[11881]), .B2(n3091), 
        .ZN(n16122) );
  MOAI22 U25036 ( .A1(n28732), .A2(n3090), .B1(ram[11882]), .B2(n3091), 
        .ZN(n16123) );
  MOAI22 U25037 ( .A1(n28497), .A2(n3090), .B1(ram[11883]), .B2(n3091), 
        .ZN(n16124) );
  MOAI22 U25038 ( .A1(n28262), .A2(n3090), .B1(ram[11884]), .B2(n3091), 
        .ZN(n16125) );
  MOAI22 U25039 ( .A1(n28027), .A2(n3090), .B1(ram[11885]), .B2(n3091), 
        .ZN(n16126) );
  MOAI22 U25040 ( .A1(n27792), .A2(n3090), .B1(ram[11886]), .B2(n3091), 
        .ZN(n16127) );
  MOAI22 U25041 ( .A1(n27557), .A2(n3090), .B1(ram[11887]), .B2(n3091), 
        .ZN(n16128) );
  MOAI22 U25042 ( .A1(n29202), .A2(n3092), .B1(ram[11888]), .B2(n3093), 
        .ZN(n16129) );
  MOAI22 U25043 ( .A1(n28967), .A2(n3092), .B1(ram[11889]), .B2(n3093), 
        .ZN(n16130) );
  MOAI22 U25044 ( .A1(n28732), .A2(n3092), .B1(ram[11890]), .B2(n3093), 
        .ZN(n16131) );
  MOAI22 U25045 ( .A1(n28497), .A2(n3092), .B1(ram[11891]), .B2(n3093), 
        .ZN(n16132) );
  MOAI22 U25046 ( .A1(n28262), .A2(n3092), .B1(ram[11892]), .B2(n3093), 
        .ZN(n16133) );
  MOAI22 U25047 ( .A1(n28027), .A2(n3092), .B1(ram[11893]), .B2(n3093), 
        .ZN(n16134) );
  MOAI22 U25048 ( .A1(n27792), .A2(n3092), .B1(ram[11894]), .B2(n3093), 
        .ZN(n16135) );
  MOAI22 U25049 ( .A1(n27557), .A2(n3092), .B1(ram[11895]), .B2(n3093), 
        .ZN(n16136) );
  MOAI22 U25050 ( .A1(n29202), .A2(n3094), .B1(ram[11896]), .B2(n3095), 
        .ZN(n16137) );
  MOAI22 U25051 ( .A1(n28967), .A2(n3094), .B1(ram[11897]), .B2(n3095), 
        .ZN(n16138) );
  MOAI22 U25052 ( .A1(n28732), .A2(n3094), .B1(ram[11898]), .B2(n3095), 
        .ZN(n16139) );
  MOAI22 U25053 ( .A1(n28497), .A2(n3094), .B1(ram[11899]), .B2(n3095), 
        .ZN(n16140) );
  MOAI22 U25054 ( .A1(n28262), .A2(n3094), .B1(ram[11900]), .B2(n3095), 
        .ZN(n16141) );
  MOAI22 U25055 ( .A1(n28027), .A2(n3094), .B1(ram[11901]), .B2(n3095), 
        .ZN(n16142) );
  MOAI22 U25056 ( .A1(n27792), .A2(n3094), .B1(ram[11902]), .B2(n3095), 
        .ZN(n16143) );
  MOAI22 U25057 ( .A1(n27557), .A2(n3094), .B1(ram[11903]), .B2(n3095), 
        .ZN(n16144) );
  MOAI22 U25058 ( .A1(n29202), .A2(n3096), .B1(ram[11904]), .B2(n3097), 
        .ZN(n16145) );
  MOAI22 U25059 ( .A1(n28967), .A2(n3096), .B1(ram[11905]), .B2(n3097), 
        .ZN(n16146) );
  MOAI22 U25060 ( .A1(n28732), .A2(n3096), .B1(ram[11906]), .B2(n3097), 
        .ZN(n16147) );
  MOAI22 U25061 ( .A1(n28497), .A2(n3096), .B1(ram[11907]), .B2(n3097), 
        .ZN(n16148) );
  MOAI22 U25062 ( .A1(n28262), .A2(n3096), .B1(ram[11908]), .B2(n3097), 
        .ZN(n16149) );
  MOAI22 U25063 ( .A1(n28027), .A2(n3096), .B1(ram[11909]), .B2(n3097), 
        .ZN(n16150) );
  MOAI22 U25064 ( .A1(n27792), .A2(n3096), .B1(ram[11910]), .B2(n3097), 
        .ZN(n16151) );
  MOAI22 U25065 ( .A1(n27557), .A2(n3096), .B1(ram[11911]), .B2(n3097), 
        .ZN(n16152) );
  MOAI22 U25066 ( .A1(n29202), .A2(n3098), .B1(ram[11912]), .B2(n3099), 
        .ZN(n16153) );
  MOAI22 U25067 ( .A1(n28967), .A2(n3098), .B1(ram[11913]), .B2(n3099), 
        .ZN(n16154) );
  MOAI22 U25068 ( .A1(n28732), .A2(n3098), .B1(ram[11914]), .B2(n3099), 
        .ZN(n16155) );
  MOAI22 U25069 ( .A1(n28497), .A2(n3098), .B1(ram[11915]), .B2(n3099), 
        .ZN(n16156) );
  MOAI22 U25070 ( .A1(n28262), .A2(n3098), .B1(ram[11916]), .B2(n3099), 
        .ZN(n16157) );
  MOAI22 U25071 ( .A1(n28027), .A2(n3098), .B1(ram[11917]), .B2(n3099), 
        .ZN(n16158) );
  MOAI22 U25072 ( .A1(n27792), .A2(n3098), .B1(ram[11918]), .B2(n3099), 
        .ZN(n16159) );
  MOAI22 U25073 ( .A1(n27557), .A2(n3098), .B1(ram[11919]), .B2(n3099), 
        .ZN(n16160) );
  MOAI22 U25074 ( .A1(n29202), .A2(n3100), .B1(ram[11920]), .B2(n3101), 
        .ZN(n16161) );
  MOAI22 U25075 ( .A1(n28967), .A2(n3100), .B1(ram[11921]), .B2(n3101), 
        .ZN(n16162) );
  MOAI22 U25076 ( .A1(n28732), .A2(n3100), .B1(ram[11922]), .B2(n3101), 
        .ZN(n16163) );
  MOAI22 U25077 ( .A1(n28497), .A2(n3100), .B1(ram[11923]), .B2(n3101), 
        .ZN(n16164) );
  MOAI22 U25078 ( .A1(n28262), .A2(n3100), .B1(ram[11924]), .B2(n3101), 
        .ZN(n16165) );
  MOAI22 U25079 ( .A1(n28027), .A2(n3100), .B1(ram[11925]), .B2(n3101), 
        .ZN(n16166) );
  MOAI22 U25080 ( .A1(n27792), .A2(n3100), .B1(ram[11926]), .B2(n3101), 
        .ZN(n16167) );
  MOAI22 U25081 ( .A1(n27557), .A2(n3100), .B1(ram[11927]), .B2(n3101), 
        .ZN(n16168) );
  MOAI22 U25082 ( .A1(n29202), .A2(n3102), .B1(ram[11928]), .B2(n3103), 
        .ZN(n16169) );
  MOAI22 U25083 ( .A1(n28967), .A2(n3102), .B1(ram[11929]), .B2(n3103), 
        .ZN(n16170) );
  MOAI22 U25084 ( .A1(n28732), .A2(n3102), .B1(ram[11930]), .B2(n3103), 
        .ZN(n16171) );
  MOAI22 U25085 ( .A1(n28497), .A2(n3102), .B1(ram[11931]), .B2(n3103), 
        .ZN(n16172) );
  MOAI22 U25086 ( .A1(n28262), .A2(n3102), .B1(ram[11932]), .B2(n3103), 
        .ZN(n16173) );
  MOAI22 U25087 ( .A1(n28027), .A2(n3102), .B1(ram[11933]), .B2(n3103), 
        .ZN(n16174) );
  MOAI22 U25088 ( .A1(n27792), .A2(n3102), .B1(ram[11934]), .B2(n3103), 
        .ZN(n16175) );
  MOAI22 U25089 ( .A1(n27557), .A2(n3102), .B1(ram[11935]), .B2(n3103), 
        .ZN(n16176) );
  MOAI22 U25090 ( .A1(n29202), .A2(n3104), .B1(ram[11936]), .B2(n3105), 
        .ZN(n16177) );
  MOAI22 U25091 ( .A1(n28967), .A2(n3104), .B1(ram[11937]), .B2(n3105), 
        .ZN(n16178) );
  MOAI22 U25092 ( .A1(n28732), .A2(n3104), .B1(ram[11938]), .B2(n3105), 
        .ZN(n16179) );
  MOAI22 U25093 ( .A1(n28497), .A2(n3104), .B1(ram[11939]), .B2(n3105), 
        .ZN(n16180) );
  MOAI22 U25094 ( .A1(n28262), .A2(n3104), .B1(ram[11940]), .B2(n3105), 
        .ZN(n16181) );
  MOAI22 U25095 ( .A1(n28027), .A2(n3104), .B1(ram[11941]), .B2(n3105), 
        .ZN(n16182) );
  MOAI22 U25096 ( .A1(n27792), .A2(n3104), .B1(ram[11942]), .B2(n3105), 
        .ZN(n16183) );
  MOAI22 U25097 ( .A1(n27557), .A2(n3104), .B1(ram[11943]), .B2(n3105), 
        .ZN(n16184) );
  MOAI22 U25098 ( .A1(n29202), .A2(n3106), .B1(ram[11944]), .B2(n3107), 
        .ZN(n16185) );
  MOAI22 U25099 ( .A1(n28967), .A2(n3106), .B1(ram[11945]), .B2(n3107), 
        .ZN(n16186) );
  MOAI22 U25100 ( .A1(n28732), .A2(n3106), .B1(ram[11946]), .B2(n3107), 
        .ZN(n16187) );
  MOAI22 U25101 ( .A1(n28497), .A2(n3106), .B1(ram[11947]), .B2(n3107), 
        .ZN(n16188) );
  MOAI22 U25102 ( .A1(n28262), .A2(n3106), .B1(ram[11948]), .B2(n3107), 
        .ZN(n16189) );
  MOAI22 U25103 ( .A1(n28027), .A2(n3106), .B1(ram[11949]), .B2(n3107), 
        .ZN(n16190) );
  MOAI22 U25104 ( .A1(n27792), .A2(n3106), .B1(ram[11950]), .B2(n3107), 
        .ZN(n16191) );
  MOAI22 U25105 ( .A1(n27557), .A2(n3106), .B1(ram[11951]), .B2(n3107), 
        .ZN(n16192) );
  MOAI22 U25106 ( .A1(n29202), .A2(n3108), .B1(ram[11952]), .B2(n3109), 
        .ZN(n16193) );
  MOAI22 U25107 ( .A1(n28967), .A2(n3108), .B1(ram[11953]), .B2(n3109), 
        .ZN(n16194) );
  MOAI22 U25108 ( .A1(n28732), .A2(n3108), .B1(ram[11954]), .B2(n3109), 
        .ZN(n16195) );
  MOAI22 U25109 ( .A1(n28497), .A2(n3108), .B1(ram[11955]), .B2(n3109), 
        .ZN(n16196) );
  MOAI22 U25110 ( .A1(n28262), .A2(n3108), .B1(ram[11956]), .B2(n3109), 
        .ZN(n16197) );
  MOAI22 U25111 ( .A1(n28027), .A2(n3108), .B1(ram[11957]), .B2(n3109), 
        .ZN(n16198) );
  MOAI22 U25112 ( .A1(n27792), .A2(n3108), .B1(ram[11958]), .B2(n3109), 
        .ZN(n16199) );
  MOAI22 U25113 ( .A1(n27557), .A2(n3108), .B1(ram[11959]), .B2(n3109), 
        .ZN(n16200) );
  MOAI22 U25114 ( .A1(n29203), .A2(n3110), .B1(ram[11960]), .B2(n3111), 
        .ZN(n16201) );
  MOAI22 U25115 ( .A1(n28968), .A2(n3110), .B1(ram[11961]), .B2(n3111), 
        .ZN(n16202) );
  MOAI22 U25116 ( .A1(n28733), .A2(n3110), .B1(ram[11962]), .B2(n3111), 
        .ZN(n16203) );
  MOAI22 U25117 ( .A1(n28498), .A2(n3110), .B1(ram[11963]), .B2(n3111), 
        .ZN(n16204) );
  MOAI22 U25118 ( .A1(n28263), .A2(n3110), .B1(ram[11964]), .B2(n3111), 
        .ZN(n16205) );
  MOAI22 U25119 ( .A1(n28028), .A2(n3110), .B1(ram[11965]), .B2(n3111), 
        .ZN(n16206) );
  MOAI22 U25120 ( .A1(n27793), .A2(n3110), .B1(ram[11966]), .B2(n3111), 
        .ZN(n16207) );
  MOAI22 U25121 ( .A1(n27558), .A2(n3110), .B1(ram[11967]), .B2(n3111), 
        .ZN(n16208) );
  MOAI22 U25122 ( .A1(n29203), .A2(n3112), .B1(ram[11968]), .B2(n3113), 
        .ZN(n16209) );
  MOAI22 U25123 ( .A1(n28968), .A2(n3112), .B1(ram[11969]), .B2(n3113), 
        .ZN(n16210) );
  MOAI22 U25124 ( .A1(n28733), .A2(n3112), .B1(ram[11970]), .B2(n3113), 
        .ZN(n16211) );
  MOAI22 U25125 ( .A1(n28498), .A2(n3112), .B1(ram[11971]), .B2(n3113), 
        .ZN(n16212) );
  MOAI22 U25126 ( .A1(n28263), .A2(n3112), .B1(ram[11972]), .B2(n3113), 
        .ZN(n16213) );
  MOAI22 U25127 ( .A1(n28028), .A2(n3112), .B1(ram[11973]), .B2(n3113), 
        .ZN(n16214) );
  MOAI22 U25128 ( .A1(n27793), .A2(n3112), .B1(ram[11974]), .B2(n3113), 
        .ZN(n16215) );
  MOAI22 U25129 ( .A1(n27558), .A2(n3112), .B1(ram[11975]), .B2(n3113), 
        .ZN(n16216) );
  MOAI22 U25130 ( .A1(n29203), .A2(n3114), .B1(ram[11976]), .B2(n3115), 
        .ZN(n16217) );
  MOAI22 U25131 ( .A1(n28968), .A2(n3114), .B1(ram[11977]), .B2(n3115), 
        .ZN(n16218) );
  MOAI22 U25132 ( .A1(n28733), .A2(n3114), .B1(ram[11978]), .B2(n3115), 
        .ZN(n16219) );
  MOAI22 U25133 ( .A1(n28498), .A2(n3114), .B1(ram[11979]), .B2(n3115), 
        .ZN(n16220) );
  MOAI22 U25134 ( .A1(n28263), .A2(n3114), .B1(ram[11980]), .B2(n3115), 
        .ZN(n16221) );
  MOAI22 U25135 ( .A1(n28028), .A2(n3114), .B1(ram[11981]), .B2(n3115), 
        .ZN(n16222) );
  MOAI22 U25136 ( .A1(n27793), .A2(n3114), .B1(ram[11982]), .B2(n3115), 
        .ZN(n16223) );
  MOAI22 U25137 ( .A1(n27558), .A2(n3114), .B1(ram[11983]), .B2(n3115), 
        .ZN(n16224) );
  MOAI22 U25138 ( .A1(n29203), .A2(n3116), .B1(ram[11984]), .B2(n3117), 
        .ZN(n16225) );
  MOAI22 U25139 ( .A1(n28968), .A2(n3116), .B1(ram[11985]), .B2(n3117), 
        .ZN(n16226) );
  MOAI22 U25140 ( .A1(n28733), .A2(n3116), .B1(ram[11986]), .B2(n3117), 
        .ZN(n16227) );
  MOAI22 U25141 ( .A1(n28498), .A2(n3116), .B1(ram[11987]), .B2(n3117), 
        .ZN(n16228) );
  MOAI22 U25142 ( .A1(n28263), .A2(n3116), .B1(ram[11988]), .B2(n3117), 
        .ZN(n16229) );
  MOAI22 U25143 ( .A1(n28028), .A2(n3116), .B1(ram[11989]), .B2(n3117), 
        .ZN(n16230) );
  MOAI22 U25144 ( .A1(n27793), .A2(n3116), .B1(ram[11990]), .B2(n3117), 
        .ZN(n16231) );
  MOAI22 U25145 ( .A1(n27558), .A2(n3116), .B1(ram[11991]), .B2(n3117), 
        .ZN(n16232) );
  MOAI22 U25146 ( .A1(n29203), .A2(n3118), .B1(ram[11992]), .B2(n3119), 
        .ZN(n16233) );
  MOAI22 U25147 ( .A1(n28968), .A2(n3118), .B1(ram[11993]), .B2(n3119), 
        .ZN(n16234) );
  MOAI22 U25148 ( .A1(n28733), .A2(n3118), .B1(ram[11994]), .B2(n3119), 
        .ZN(n16235) );
  MOAI22 U25149 ( .A1(n28498), .A2(n3118), .B1(ram[11995]), .B2(n3119), 
        .ZN(n16236) );
  MOAI22 U25150 ( .A1(n28263), .A2(n3118), .B1(ram[11996]), .B2(n3119), 
        .ZN(n16237) );
  MOAI22 U25151 ( .A1(n28028), .A2(n3118), .B1(ram[11997]), .B2(n3119), 
        .ZN(n16238) );
  MOAI22 U25152 ( .A1(n27793), .A2(n3118), .B1(ram[11998]), .B2(n3119), 
        .ZN(n16239) );
  MOAI22 U25153 ( .A1(n27558), .A2(n3118), .B1(ram[11999]), .B2(n3119), 
        .ZN(n16240) );
  MOAI22 U25154 ( .A1(n29203), .A2(n3120), .B1(ram[12000]), .B2(n3121), 
        .ZN(n16241) );
  MOAI22 U25155 ( .A1(n28968), .A2(n3120), .B1(ram[12001]), .B2(n3121), 
        .ZN(n16242) );
  MOAI22 U25156 ( .A1(n28733), .A2(n3120), .B1(ram[12002]), .B2(n3121), 
        .ZN(n16243) );
  MOAI22 U25157 ( .A1(n28498), .A2(n3120), .B1(ram[12003]), .B2(n3121), 
        .ZN(n16244) );
  MOAI22 U25158 ( .A1(n28263), .A2(n3120), .B1(ram[12004]), .B2(n3121), 
        .ZN(n16245) );
  MOAI22 U25159 ( .A1(n28028), .A2(n3120), .B1(ram[12005]), .B2(n3121), 
        .ZN(n16246) );
  MOAI22 U25160 ( .A1(n27793), .A2(n3120), .B1(ram[12006]), .B2(n3121), 
        .ZN(n16247) );
  MOAI22 U25161 ( .A1(n27558), .A2(n3120), .B1(ram[12007]), .B2(n3121), 
        .ZN(n16248) );
  MOAI22 U25162 ( .A1(n29203), .A2(n3122), .B1(ram[12008]), .B2(n3123), 
        .ZN(n16249) );
  MOAI22 U25163 ( .A1(n28968), .A2(n3122), .B1(ram[12009]), .B2(n3123), 
        .ZN(n16250) );
  MOAI22 U25164 ( .A1(n28733), .A2(n3122), .B1(ram[12010]), .B2(n3123), 
        .ZN(n16251) );
  MOAI22 U25165 ( .A1(n28498), .A2(n3122), .B1(ram[12011]), .B2(n3123), 
        .ZN(n16252) );
  MOAI22 U25166 ( .A1(n28263), .A2(n3122), .B1(ram[12012]), .B2(n3123), 
        .ZN(n16253) );
  MOAI22 U25167 ( .A1(n28028), .A2(n3122), .B1(ram[12013]), .B2(n3123), 
        .ZN(n16254) );
  MOAI22 U25168 ( .A1(n27793), .A2(n3122), .B1(ram[12014]), .B2(n3123), 
        .ZN(n16255) );
  MOAI22 U25169 ( .A1(n27558), .A2(n3122), .B1(ram[12015]), .B2(n3123), 
        .ZN(n16256) );
  MOAI22 U25170 ( .A1(n29203), .A2(n3124), .B1(ram[12016]), .B2(n3125), 
        .ZN(n16257) );
  MOAI22 U25171 ( .A1(n28968), .A2(n3124), .B1(ram[12017]), .B2(n3125), 
        .ZN(n16258) );
  MOAI22 U25172 ( .A1(n28733), .A2(n3124), .B1(ram[12018]), .B2(n3125), 
        .ZN(n16259) );
  MOAI22 U25173 ( .A1(n28498), .A2(n3124), .B1(ram[12019]), .B2(n3125), 
        .ZN(n16260) );
  MOAI22 U25174 ( .A1(n28263), .A2(n3124), .B1(ram[12020]), .B2(n3125), 
        .ZN(n16261) );
  MOAI22 U25175 ( .A1(n28028), .A2(n3124), .B1(ram[12021]), .B2(n3125), 
        .ZN(n16262) );
  MOAI22 U25176 ( .A1(n27793), .A2(n3124), .B1(ram[12022]), .B2(n3125), 
        .ZN(n16263) );
  MOAI22 U25177 ( .A1(n27558), .A2(n3124), .B1(ram[12023]), .B2(n3125), 
        .ZN(n16264) );
  MOAI22 U25178 ( .A1(n29203), .A2(n3126), .B1(ram[12024]), .B2(n3127), 
        .ZN(n16265) );
  MOAI22 U25179 ( .A1(n28968), .A2(n3126), .B1(ram[12025]), .B2(n3127), 
        .ZN(n16266) );
  MOAI22 U25180 ( .A1(n28733), .A2(n3126), .B1(ram[12026]), .B2(n3127), 
        .ZN(n16267) );
  MOAI22 U25181 ( .A1(n28498), .A2(n3126), .B1(ram[12027]), .B2(n3127), 
        .ZN(n16268) );
  MOAI22 U25182 ( .A1(n28263), .A2(n3126), .B1(ram[12028]), .B2(n3127), 
        .ZN(n16269) );
  MOAI22 U25183 ( .A1(n28028), .A2(n3126), .B1(ram[12029]), .B2(n3127), 
        .ZN(n16270) );
  MOAI22 U25184 ( .A1(n27793), .A2(n3126), .B1(ram[12030]), .B2(n3127), 
        .ZN(n16271) );
  MOAI22 U25185 ( .A1(n27558), .A2(n3126), .B1(ram[12031]), .B2(n3127), 
        .ZN(n16272) );
  MOAI22 U25186 ( .A1(n29203), .A2(n3128), .B1(ram[12032]), .B2(n3129), 
        .ZN(n16273) );
  MOAI22 U25187 ( .A1(n28968), .A2(n3128), .B1(ram[12033]), .B2(n3129), 
        .ZN(n16274) );
  MOAI22 U25188 ( .A1(n28733), .A2(n3128), .B1(ram[12034]), .B2(n3129), 
        .ZN(n16275) );
  MOAI22 U25189 ( .A1(n28498), .A2(n3128), .B1(ram[12035]), .B2(n3129), 
        .ZN(n16276) );
  MOAI22 U25190 ( .A1(n28263), .A2(n3128), .B1(ram[12036]), .B2(n3129), 
        .ZN(n16277) );
  MOAI22 U25191 ( .A1(n28028), .A2(n3128), .B1(ram[12037]), .B2(n3129), 
        .ZN(n16278) );
  MOAI22 U25192 ( .A1(n27793), .A2(n3128), .B1(ram[12038]), .B2(n3129), 
        .ZN(n16279) );
  MOAI22 U25193 ( .A1(n27558), .A2(n3128), .B1(ram[12039]), .B2(n3129), 
        .ZN(n16280) );
  MOAI22 U25194 ( .A1(n29203), .A2(n3130), .B1(ram[12040]), .B2(n3131), 
        .ZN(n16281) );
  MOAI22 U25195 ( .A1(n28968), .A2(n3130), .B1(ram[12041]), .B2(n3131), 
        .ZN(n16282) );
  MOAI22 U25196 ( .A1(n28733), .A2(n3130), .B1(ram[12042]), .B2(n3131), 
        .ZN(n16283) );
  MOAI22 U25197 ( .A1(n28498), .A2(n3130), .B1(ram[12043]), .B2(n3131), 
        .ZN(n16284) );
  MOAI22 U25198 ( .A1(n28263), .A2(n3130), .B1(ram[12044]), .B2(n3131), 
        .ZN(n16285) );
  MOAI22 U25199 ( .A1(n28028), .A2(n3130), .B1(ram[12045]), .B2(n3131), 
        .ZN(n16286) );
  MOAI22 U25200 ( .A1(n27793), .A2(n3130), .B1(ram[12046]), .B2(n3131), 
        .ZN(n16287) );
  MOAI22 U25201 ( .A1(n27558), .A2(n3130), .B1(ram[12047]), .B2(n3131), 
        .ZN(n16288) );
  MOAI22 U25202 ( .A1(n29203), .A2(n3132), .B1(ram[12048]), .B2(n3133), 
        .ZN(n16289) );
  MOAI22 U25203 ( .A1(n28968), .A2(n3132), .B1(ram[12049]), .B2(n3133), 
        .ZN(n16290) );
  MOAI22 U25204 ( .A1(n28733), .A2(n3132), .B1(ram[12050]), .B2(n3133), 
        .ZN(n16291) );
  MOAI22 U25205 ( .A1(n28498), .A2(n3132), .B1(ram[12051]), .B2(n3133), 
        .ZN(n16292) );
  MOAI22 U25206 ( .A1(n28263), .A2(n3132), .B1(ram[12052]), .B2(n3133), 
        .ZN(n16293) );
  MOAI22 U25207 ( .A1(n28028), .A2(n3132), .B1(ram[12053]), .B2(n3133), 
        .ZN(n16294) );
  MOAI22 U25208 ( .A1(n27793), .A2(n3132), .B1(ram[12054]), .B2(n3133), 
        .ZN(n16295) );
  MOAI22 U25209 ( .A1(n27558), .A2(n3132), .B1(ram[12055]), .B2(n3133), 
        .ZN(n16296) );
  MOAI22 U25210 ( .A1(n29203), .A2(n3134), .B1(ram[12056]), .B2(n3135), 
        .ZN(n16297) );
  MOAI22 U25211 ( .A1(n28968), .A2(n3134), .B1(ram[12057]), .B2(n3135), 
        .ZN(n16298) );
  MOAI22 U25212 ( .A1(n28733), .A2(n3134), .B1(ram[12058]), .B2(n3135), 
        .ZN(n16299) );
  MOAI22 U25213 ( .A1(n28498), .A2(n3134), .B1(ram[12059]), .B2(n3135), 
        .ZN(n16300) );
  MOAI22 U25214 ( .A1(n28263), .A2(n3134), .B1(ram[12060]), .B2(n3135), 
        .ZN(n16301) );
  MOAI22 U25215 ( .A1(n28028), .A2(n3134), .B1(ram[12061]), .B2(n3135), 
        .ZN(n16302) );
  MOAI22 U25216 ( .A1(n27793), .A2(n3134), .B1(ram[12062]), .B2(n3135), 
        .ZN(n16303) );
  MOAI22 U25217 ( .A1(n27558), .A2(n3134), .B1(ram[12063]), .B2(n3135), 
        .ZN(n16304) );
  MOAI22 U25218 ( .A1(n29204), .A2(n3136), .B1(ram[12064]), .B2(n3137), 
        .ZN(n16305) );
  MOAI22 U25219 ( .A1(n28969), .A2(n3136), .B1(ram[12065]), .B2(n3137), 
        .ZN(n16306) );
  MOAI22 U25220 ( .A1(n28734), .A2(n3136), .B1(ram[12066]), .B2(n3137), 
        .ZN(n16307) );
  MOAI22 U25221 ( .A1(n28499), .A2(n3136), .B1(ram[12067]), .B2(n3137), 
        .ZN(n16308) );
  MOAI22 U25222 ( .A1(n28264), .A2(n3136), .B1(ram[12068]), .B2(n3137), 
        .ZN(n16309) );
  MOAI22 U25223 ( .A1(n28029), .A2(n3136), .B1(ram[12069]), .B2(n3137), 
        .ZN(n16310) );
  MOAI22 U25224 ( .A1(n27794), .A2(n3136), .B1(ram[12070]), .B2(n3137), 
        .ZN(n16311) );
  MOAI22 U25225 ( .A1(n27559), .A2(n3136), .B1(ram[12071]), .B2(n3137), 
        .ZN(n16312) );
  MOAI22 U25226 ( .A1(n29204), .A2(n3138), .B1(ram[12072]), .B2(n3139), 
        .ZN(n16313) );
  MOAI22 U25227 ( .A1(n28969), .A2(n3138), .B1(ram[12073]), .B2(n3139), 
        .ZN(n16314) );
  MOAI22 U25228 ( .A1(n28734), .A2(n3138), .B1(ram[12074]), .B2(n3139), 
        .ZN(n16315) );
  MOAI22 U25229 ( .A1(n28499), .A2(n3138), .B1(ram[12075]), .B2(n3139), 
        .ZN(n16316) );
  MOAI22 U25230 ( .A1(n28264), .A2(n3138), .B1(ram[12076]), .B2(n3139), 
        .ZN(n16317) );
  MOAI22 U25231 ( .A1(n28029), .A2(n3138), .B1(ram[12077]), .B2(n3139), 
        .ZN(n16318) );
  MOAI22 U25232 ( .A1(n27794), .A2(n3138), .B1(ram[12078]), .B2(n3139), 
        .ZN(n16319) );
  MOAI22 U25233 ( .A1(n27559), .A2(n3138), .B1(ram[12079]), .B2(n3139), 
        .ZN(n16320) );
  MOAI22 U25234 ( .A1(n29204), .A2(n3140), .B1(ram[12080]), .B2(n3141), 
        .ZN(n16321) );
  MOAI22 U25235 ( .A1(n28969), .A2(n3140), .B1(ram[12081]), .B2(n3141), 
        .ZN(n16322) );
  MOAI22 U25236 ( .A1(n28734), .A2(n3140), .B1(ram[12082]), .B2(n3141), 
        .ZN(n16323) );
  MOAI22 U25237 ( .A1(n28499), .A2(n3140), .B1(ram[12083]), .B2(n3141), 
        .ZN(n16324) );
  MOAI22 U25238 ( .A1(n28264), .A2(n3140), .B1(ram[12084]), .B2(n3141), 
        .ZN(n16325) );
  MOAI22 U25239 ( .A1(n28029), .A2(n3140), .B1(ram[12085]), .B2(n3141), 
        .ZN(n16326) );
  MOAI22 U25240 ( .A1(n27794), .A2(n3140), .B1(ram[12086]), .B2(n3141), 
        .ZN(n16327) );
  MOAI22 U25241 ( .A1(n27559), .A2(n3140), .B1(ram[12087]), .B2(n3141), 
        .ZN(n16328) );
  MOAI22 U25242 ( .A1(n29204), .A2(n3142), .B1(ram[12088]), .B2(n3143), 
        .ZN(n16329) );
  MOAI22 U25243 ( .A1(n28969), .A2(n3142), .B1(ram[12089]), .B2(n3143), 
        .ZN(n16330) );
  MOAI22 U25244 ( .A1(n28734), .A2(n3142), .B1(ram[12090]), .B2(n3143), 
        .ZN(n16331) );
  MOAI22 U25245 ( .A1(n28499), .A2(n3142), .B1(ram[12091]), .B2(n3143), 
        .ZN(n16332) );
  MOAI22 U25246 ( .A1(n28264), .A2(n3142), .B1(ram[12092]), .B2(n3143), 
        .ZN(n16333) );
  MOAI22 U25247 ( .A1(n28029), .A2(n3142), .B1(ram[12093]), .B2(n3143), 
        .ZN(n16334) );
  MOAI22 U25248 ( .A1(n27794), .A2(n3142), .B1(ram[12094]), .B2(n3143), 
        .ZN(n16335) );
  MOAI22 U25249 ( .A1(n27559), .A2(n3142), .B1(ram[12095]), .B2(n3143), 
        .ZN(n16336) );
  MOAI22 U25250 ( .A1(n29204), .A2(n3144), .B1(ram[12096]), .B2(n3145), 
        .ZN(n16337) );
  MOAI22 U25251 ( .A1(n28969), .A2(n3144), .B1(ram[12097]), .B2(n3145), 
        .ZN(n16338) );
  MOAI22 U25252 ( .A1(n28734), .A2(n3144), .B1(ram[12098]), .B2(n3145), 
        .ZN(n16339) );
  MOAI22 U25253 ( .A1(n28499), .A2(n3144), .B1(ram[12099]), .B2(n3145), 
        .ZN(n16340) );
  MOAI22 U25254 ( .A1(n28264), .A2(n3144), .B1(ram[12100]), .B2(n3145), 
        .ZN(n16341) );
  MOAI22 U25255 ( .A1(n28029), .A2(n3144), .B1(ram[12101]), .B2(n3145), 
        .ZN(n16342) );
  MOAI22 U25256 ( .A1(n27794), .A2(n3144), .B1(ram[12102]), .B2(n3145), 
        .ZN(n16343) );
  MOAI22 U25257 ( .A1(n27559), .A2(n3144), .B1(ram[12103]), .B2(n3145), 
        .ZN(n16344) );
  MOAI22 U25258 ( .A1(n29204), .A2(n3146), .B1(ram[12104]), .B2(n3147), 
        .ZN(n16345) );
  MOAI22 U25259 ( .A1(n28969), .A2(n3146), .B1(ram[12105]), .B2(n3147), 
        .ZN(n16346) );
  MOAI22 U25260 ( .A1(n28734), .A2(n3146), .B1(ram[12106]), .B2(n3147), 
        .ZN(n16347) );
  MOAI22 U25261 ( .A1(n28499), .A2(n3146), .B1(ram[12107]), .B2(n3147), 
        .ZN(n16348) );
  MOAI22 U25262 ( .A1(n28264), .A2(n3146), .B1(ram[12108]), .B2(n3147), 
        .ZN(n16349) );
  MOAI22 U25263 ( .A1(n28029), .A2(n3146), .B1(ram[12109]), .B2(n3147), 
        .ZN(n16350) );
  MOAI22 U25264 ( .A1(n27794), .A2(n3146), .B1(ram[12110]), .B2(n3147), 
        .ZN(n16351) );
  MOAI22 U25265 ( .A1(n27559), .A2(n3146), .B1(ram[12111]), .B2(n3147), 
        .ZN(n16352) );
  MOAI22 U25266 ( .A1(n29204), .A2(n3148), .B1(ram[12112]), .B2(n3149), 
        .ZN(n16353) );
  MOAI22 U25267 ( .A1(n28969), .A2(n3148), .B1(ram[12113]), .B2(n3149), 
        .ZN(n16354) );
  MOAI22 U25268 ( .A1(n28734), .A2(n3148), .B1(ram[12114]), .B2(n3149), 
        .ZN(n16355) );
  MOAI22 U25269 ( .A1(n28499), .A2(n3148), .B1(ram[12115]), .B2(n3149), 
        .ZN(n16356) );
  MOAI22 U25270 ( .A1(n28264), .A2(n3148), .B1(ram[12116]), .B2(n3149), 
        .ZN(n16357) );
  MOAI22 U25271 ( .A1(n28029), .A2(n3148), .B1(ram[12117]), .B2(n3149), 
        .ZN(n16358) );
  MOAI22 U25272 ( .A1(n27794), .A2(n3148), .B1(ram[12118]), .B2(n3149), 
        .ZN(n16359) );
  MOAI22 U25273 ( .A1(n27559), .A2(n3148), .B1(ram[12119]), .B2(n3149), 
        .ZN(n16360) );
  MOAI22 U25274 ( .A1(n29204), .A2(n3150), .B1(ram[12120]), .B2(n3151), 
        .ZN(n16361) );
  MOAI22 U25275 ( .A1(n28969), .A2(n3150), .B1(ram[12121]), .B2(n3151), 
        .ZN(n16362) );
  MOAI22 U25276 ( .A1(n28734), .A2(n3150), .B1(ram[12122]), .B2(n3151), 
        .ZN(n16363) );
  MOAI22 U25277 ( .A1(n28499), .A2(n3150), .B1(ram[12123]), .B2(n3151), 
        .ZN(n16364) );
  MOAI22 U25278 ( .A1(n28264), .A2(n3150), .B1(ram[12124]), .B2(n3151), 
        .ZN(n16365) );
  MOAI22 U25279 ( .A1(n28029), .A2(n3150), .B1(ram[12125]), .B2(n3151), 
        .ZN(n16366) );
  MOAI22 U25280 ( .A1(n27794), .A2(n3150), .B1(ram[12126]), .B2(n3151), 
        .ZN(n16367) );
  MOAI22 U25281 ( .A1(n27559), .A2(n3150), .B1(ram[12127]), .B2(n3151), 
        .ZN(n16368) );
  MOAI22 U25282 ( .A1(n29204), .A2(n3152), .B1(ram[12128]), .B2(n3153), 
        .ZN(n16369) );
  MOAI22 U25283 ( .A1(n28969), .A2(n3152), .B1(ram[12129]), .B2(n3153), 
        .ZN(n16370) );
  MOAI22 U25284 ( .A1(n28734), .A2(n3152), .B1(ram[12130]), .B2(n3153), 
        .ZN(n16371) );
  MOAI22 U25285 ( .A1(n28499), .A2(n3152), .B1(ram[12131]), .B2(n3153), 
        .ZN(n16372) );
  MOAI22 U25286 ( .A1(n28264), .A2(n3152), .B1(ram[12132]), .B2(n3153), 
        .ZN(n16373) );
  MOAI22 U25287 ( .A1(n28029), .A2(n3152), .B1(ram[12133]), .B2(n3153), 
        .ZN(n16374) );
  MOAI22 U25288 ( .A1(n27794), .A2(n3152), .B1(ram[12134]), .B2(n3153), 
        .ZN(n16375) );
  MOAI22 U25289 ( .A1(n27559), .A2(n3152), .B1(ram[12135]), .B2(n3153), 
        .ZN(n16376) );
  MOAI22 U25290 ( .A1(n29204), .A2(n3154), .B1(ram[12136]), .B2(n3155), 
        .ZN(n16377) );
  MOAI22 U25291 ( .A1(n28969), .A2(n3154), .B1(ram[12137]), .B2(n3155), 
        .ZN(n16378) );
  MOAI22 U25292 ( .A1(n28734), .A2(n3154), .B1(ram[12138]), .B2(n3155), 
        .ZN(n16379) );
  MOAI22 U25293 ( .A1(n28499), .A2(n3154), .B1(ram[12139]), .B2(n3155), 
        .ZN(n16380) );
  MOAI22 U25294 ( .A1(n28264), .A2(n3154), .B1(ram[12140]), .B2(n3155), 
        .ZN(n16381) );
  MOAI22 U25295 ( .A1(n28029), .A2(n3154), .B1(ram[12141]), .B2(n3155), 
        .ZN(n16382) );
  MOAI22 U25296 ( .A1(n27794), .A2(n3154), .B1(ram[12142]), .B2(n3155), 
        .ZN(n16383) );
  MOAI22 U25297 ( .A1(n27559), .A2(n3154), .B1(ram[12143]), .B2(n3155), 
        .ZN(n16384) );
  MOAI22 U25298 ( .A1(n29204), .A2(n3156), .B1(ram[12144]), .B2(n3157), 
        .ZN(n16385) );
  MOAI22 U25299 ( .A1(n28969), .A2(n3156), .B1(ram[12145]), .B2(n3157), 
        .ZN(n16386) );
  MOAI22 U25300 ( .A1(n28734), .A2(n3156), .B1(ram[12146]), .B2(n3157), 
        .ZN(n16387) );
  MOAI22 U25301 ( .A1(n28499), .A2(n3156), .B1(ram[12147]), .B2(n3157), 
        .ZN(n16388) );
  MOAI22 U25302 ( .A1(n28264), .A2(n3156), .B1(ram[12148]), .B2(n3157), 
        .ZN(n16389) );
  MOAI22 U25303 ( .A1(n28029), .A2(n3156), .B1(ram[12149]), .B2(n3157), 
        .ZN(n16390) );
  MOAI22 U25304 ( .A1(n27794), .A2(n3156), .B1(ram[12150]), .B2(n3157), 
        .ZN(n16391) );
  MOAI22 U25305 ( .A1(n27559), .A2(n3156), .B1(ram[12151]), .B2(n3157), 
        .ZN(n16392) );
  MOAI22 U25306 ( .A1(n29204), .A2(n3158), .B1(ram[12152]), .B2(n3159), 
        .ZN(n16393) );
  MOAI22 U25307 ( .A1(n28969), .A2(n3158), .B1(ram[12153]), .B2(n3159), 
        .ZN(n16394) );
  MOAI22 U25308 ( .A1(n28734), .A2(n3158), .B1(ram[12154]), .B2(n3159), 
        .ZN(n16395) );
  MOAI22 U25309 ( .A1(n28499), .A2(n3158), .B1(ram[12155]), .B2(n3159), 
        .ZN(n16396) );
  MOAI22 U25310 ( .A1(n28264), .A2(n3158), .B1(ram[12156]), .B2(n3159), 
        .ZN(n16397) );
  MOAI22 U25311 ( .A1(n28029), .A2(n3158), .B1(ram[12157]), .B2(n3159), 
        .ZN(n16398) );
  MOAI22 U25312 ( .A1(n27794), .A2(n3158), .B1(ram[12158]), .B2(n3159), 
        .ZN(n16399) );
  MOAI22 U25313 ( .A1(n27559), .A2(n3158), .B1(ram[12159]), .B2(n3159), 
        .ZN(n16400) );
  MOAI22 U25314 ( .A1(n29204), .A2(n3160), .B1(ram[12160]), .B2(n3161), 
        .ZN(n16401) );
  MOAI22 U25315 ( .A1(n28969), .A2(n3160), .B1(ram[12161]), .B2(n3161), 
        .ZN(n16402) );
  MOAI22 U25316 ( .A1(n28734), .A2(n3160), .B1(ram[12162]), .B2(n3161), 
        .ZN(n16403) );
  MOAI22 U25317 ( .A1(n28499), .A2(n3160), .B1(ram[12163]), .B2(n3161), 
        .ZN(n16404) );
  MOAI22 U25318 ( .A1(n28264), .A2(n3160), .B1(ram[12164]), .B2(n3161), 
        .ZN(n16405) );
  MOAI22 U25319 ( .A1(n28029), .A2(n3160), .B1(ram[12165]), .B2(n3161), 
        .ZN(n16406) );
  MOAI22 U25320 ( .A1(n27794), .A2(n3160), .B1(ram[12166]), .B2(n3161), 
        .ZN(n16407) );
  MOAI22 U25321 ( .A1(n27559), .A2(n3160), .B1(ram[12167]), .B2(n3161), 
        .ZN(n16408) );
  MOAI22 U25322 ( .A1(n29205), .A2(n3162), .B1(ram[12168]), .B2(n3163), 
        .ZN(n16409) );
  MOAI22 U25323 ( .A1(n28970), .A2(n3162), .B1(ram[12169]), .B2(n3163), 
        .ZN(n16410) );
  MOAI22 U25324 ( .A1(n28735), .A2(n3162), .B1(ram[12170]), .B2(n3163), 
        .ZN(n16411) );
  MOAI22 U25325 ( .A1(n28500), .A2(n3162), .B1(ram[12171]), .B2(n3163), 
        .ZN(n16412) );
  MOAI22 U25326 ( .A1(n28265), .A2(n3162), .B1(ram[12172]), .B2(n3163), 
        .ZN(n16413) );
  MOAI22 U25327 ( .A1(n28030), .A2(n3162), .B1(ram[12173]), .B2(n3163), 
        .ZN(n16414) );
  MOAI22 U25328 ( .A1(n27795), .A2(n3162), .B1(ram[12174]), .B2(n3163), 
        .ZN(n16415) );
  MOAI22 U25329 ( .A1(n27560), .A2(n3162), .B1(ram[12175]), .B2(n3163), 
        .ZN(n16416) );
  MOAI22 U25330 ( .A1(n29205), .A2(n3164), .B1(ram[12176]), .B2(n3165), 
        .ZN(n16417) );
  MOAI22 U25331 ( .A1(n28970), .A2(n3164), .B1(ram[12177]), .B2(n3165), 
        .ZN(n16418) );
  MOAI22 U25332 ( .A1(n28735), .A2(n3164), .B1(ram[12178]), .B2(n3165), 
        .ZN(n16419) );
  MOAI22 U25333 ( .A1(n28500), .A2(n3164), .B1(ram[12179]), .B2(n3165), 
        .ZN(n16420) );
  MOAI22 U25334 ( .A1(n28265), .A2(n3164), .B1(ram[12180]), .B2(n3165), 
        .ZN(n16421) );
  MOAI22 U25335 ( .A1(n28030), .A2(n3164), .B1(ram[12181]), .B2(n3165), 
        .ZN(n16422) );
  MOAI22 U25336 ( .A1(n27795), .A2(n3164), .B1(ram[12182]), .B2(n3165), 
        .ZN(n16423) );
  MOAI22 U25337 ( .A1(n27560), .A2(n3164), .B1(ram[12183]), .B2(n3165), 
        .ZN(n16424) );
  MOAI22 U25338 ( .A1(n29205), .A2(n3166), .B1(ram[12184]), .B2(n3167), 
        .ZN(n16425) );
  MOAI22 U25339 ( .A1(n28970), .A2(n3166), .B1(ram[12185]), .B2(n3167), 
        .ZN(n16426) );
  MOAI22 U25340 ( .A1(n28735), .A2(n3166), .B1(ram[12186]), .B2(n3167), 
        .ZN(n16427) );
  MOAI22 U25341 ( .A1(n28500), .A2(n3166), .B1(ram[12187]), .B2(n3167), 
        .ZN(n16428) );
  MOAI22 U25342 ( .A1(n28265), .A2(n3166), .B1(ram[12188]), .B2(n3167), 
        .ZN(n16429) );
  MOAI22 U25343 ( .A1(n28030), .A2(n3166), .B1(ram[12189]), .B2(n3167), 
        .ZN(n16430) );
  MOAI22 U25344 ( .A1(n27795), .A2(n3166), .B1(ram[12190]), .B2(n3167), 
        .ZN(n16431) );
  MOAI22 U25345 ( .A1(n27560), .A2(n3166), .B1(ram[12191]), .B2(n3167), 
        .ZN(n16432) );
  MOAI22 U25346 ( .A1(n29205), .A2(n3168), .B1(ram[12192]), .B2(n3169), 
        .ZN(n16433) );
  MOAI22 U25347 ( .A1(n28970), .A2(n3168), .B1(ram[12193]), .B2(n3169), 
        .ZN(n16434) );
  MOAI22 U25348 ( .A1(n28735), .A2(n3168), .B1(ram[12194]), .B2(n3169), 
        .ZN(n16435) );
  MOAI22 U25349 ( .A1(n28500), .A2(n3168), .B1(ram[12195]), .B2(n3169), 
        .ZN(n16436) );
  MOAI22 U25350 ( .A1(n28265), .A2(n3168), .B1(ram[12196]), .B2(n3169), 
        .ZN(n16437) );
  MOAI22 U25351 ( .A1(n28030), .A2(n3168), .B1(ram[12197]), .B2(n3169), 
        .ZN(n16438) );
  MOAI22 U25352 ( .A1(n27795), .A2(n3168), .B1(ram[12198]), .B2(n3169), 
        .ZN(n16439) );
  MOAI22 U25353 ( .A1(n27560), .A2(n3168), .B1(ram[12199]), .B2(n3169), 
        .ZN(n16440) );
  MOAI22 U25354 ( .A1(n29205), .A2(n3170), .B1(ram[12200]), .B2(n3171), 
        .ZN(n16441) );
  MOAI22 U25355 ( .A1(n28970), .A2(n3170), .B1(ram[12201]), .B2(n3171), 
        .ZN(n16442) );
  MOAI22 U25356 ( .A1(n28735), .A2(n3170), .B1(ram[12202]), .B2(n3171), 
        .ZN(n16443) );
  MOAI22 U25357 ( .A1(n28500), .A2(n3170), .B1(ram[12203]), .B2(n3171), 
        .ZN(n16444) );
  MOAI22 U25358 ( .A1(n28265), .A2(n3170), .B1(ram[12204]), .B2(n3171), 
        .ZN(n16445) );
  MOAI22 U25359 ( .A1(n28030), .A2(n3170), .B1(ram[12205]), .B2(n3171), 
        .ZN(n16446) );
  MOAI22 U25360 ( .A1(n27795), .A2(n3170), .B1(ram[12206]), .B2(n3171), 
        .ZN(n16447) );
  MOAI22 U25361 ( .A1(n27560), .A2(n3170), .B1(ram[12207]), .B2(n3171), 
        .ZN(n16448) );
  MOAI22 U25362 ( .A1(n29205), .A2(n3172), .B1(ram[12208]), .B2(n3173), 
        .ZN(n16449) );
  MOAI22 U25363 ( .A1(n28970), .A2(n3172), .B1(ram[12209]), .B2(n3173), 
        .ZN(n16450) );
  MOAI22 U25364 ( .A1(n28735), .A2(n3172), .B1(ram[12210]), .B2(n3173), 
        .ZN(n16451) );
  MOAI22 U25365 ( .A1(n28500), .A2(n3172), .B1(ram[12211]), .B2(n3173), 
        .ZN(n16452) );
  MOAI22 U25366 ( .A1(n28265), .A2(n3172), .B1(ram[12212]), .B2(n3173), 
        .ZN(n16453) );
  MOAI22 U25367 ( .A1(n28030), .A2(n3172), .B1(ram[12213]), .B2(n3173), 
        .ZN(n16454) );
  MOAI22 U25368 ( .A1(n27795), .A2(n3172), .B1(ram[12214]), .B2(n3173), 
        .ZN(n16455) );
  MOAI22 U25369 ( .A1(n27560), .A2(n3172), .B1(ram[12215]), .B2(n3173), 
        .ZN(n16456) );
  MOAI22 U25370 ( .A1(n29205), .A2(n3174), .B1(ram[12216]), .B2(n3175), 
        .ZN(n16457) );
  MOAI22 U25371 ( .A1(n28970), .A2(n3174), .B1(ram[12217]), .B2(n3175), 
        .ZN(n16458) );
  MOAI22 U25372 ( .A1(n28735), .A2(n3174), .B1(ram[12218]), .B2(n3175), 
        .ZN(n16459) );
  MOAI22 U25373 ( .A1(n28500), .A2(n3174), .B1(ram[12219]), .B2(n3175), 
        .ZN(n16460) );
  MOAI22 U25374 ( .A1(n28265), .A2(n3174), .B1(ram[12220]), .B2(n3175), 
        .ZN(n16461) );
  MOAI22 U25375 ( .A1(n28030), .A2(n3174), .B1(ram[12221]), .B2(n3175), 
        .ZN(n16462) );
  MOAI22 U25376 ( .A1(n27795), .A2(n3174), .B1(ram[12222]), .B2(n3175), 
        .ZN(n16463) );
  MOAI22 U25377 ( .A1(n27560), .A2(n3174), .B1(ram[12223]), .B2(n3175), 
        .ZN(n16464) );
  MOAI22 U25378 ( .A1(n29205), .A2(n3176), .B1(ram[12224]), .B2(n3177), 
        .ZN(n16465) );
  MOAI22 U25379 ( .A1(n28970), .A2(n3176), .B1(ram[12225]), .B2(n3177), 
        .ZN(n16466) );
  MOAI22 U25380 ( .A1(n28735), .A2(n3176), .B1(ram[12226]), .B2(n3177), 
        .ZN(n16467) );
  MOAI22 U25381 ( .A1(n28500), .A2(n3176), .B1(ram[12227]), .B2(n3177), 
        .ZN(n16468) );
  MOAI22 U25382 ( .A1(n28265), .A2(n3176), .B1(ram[12228]), .B2(n3177), 
        .ZN(n16469) );
  MOAI22 U25383 ( .A1(n28030), .A2(n3176), .B1(ram[12229]), .B2(n3177), 
        .ZN(n16470) );
  MOAI22 U25384 ( .A1(n27795), .A2(n3176), .B1(ram[12230]), .B2(n3177), 
        .ZN(n16471) );
  MOAI22 U25385 ( .A1(n27560), .A2(n3176), .B1(ram[12231]), .B2(n3177), 
        .ZN(n16472) );
  MOAI22 U25386 ( .A1(n29205), .A2(n3178), .B1(ram[12232]), .B2(n3179), 
        .ZN(n16473) );
  MOAI22 U25387 ( .A1(n28970), .A2(n3178), .B1(ram[12233]), .B2(n3179), 
        .ZN(n16474) );
  MOAI22 U25388 ( .A1(n28735), .A2(n3178), .B1(ram[12234]), .B2(n3179), 
        .ZN(n16475) );
  MOAI22 U25389 ( .A1(n28500), .A2(n3178), .B1(ram[12235]), .B2(n3179), 
        .ZN(n16476) );
  MOAI22 U25390 ( .A1(n28265), .A2(n3178), .B1(ram[12236]), .B2(n3179), 
        .ZN(n16477) );
  MOAI22 U25391 ( .A1(n28030), .A2(n3178), .B1(ram[12237]), .B2(n3179), 
        .ZN(n16478) );
  MOAI22 U25392 ( .A1(n27795), .A2(n3178), .B1(ram[12238]), .B2(n3179), 
        .ZN(n16479) );
  MOAI22 U25393 ( .A1(n27560), .A2(n3178), .B1(ram[12239]), .B2(n3179), 
        .ZN(n16480) );
  MOAI22 U25394 ( .A1(n29205), .A2(n3180), .B1(ram[12240]), .B2(n3181), 
        .ZN(n16481) );
  MOAI22 U25395 ( .A1(n28970), .A2(n3180), .B1(ram[12241]), .B2(n3181), 
        .ZN(n16482) );
  MOAI22 U25396 ( .A1(n28735), .A2(n3180), .B1(ram[12242]), .B2(n3181), 
        .ZN(n16483) );
  MOAI22 U25397 ( .A1(n28500), .A2(n3180), .B1(ram[12243]), .B2(n3181), 
        .ZN(n16484) );
  MOAI22 U25398 ( .A1(n28265), .A2(n3180), .B1(ram[12244]), .B2(n3181), 
        .ZN(n16485) );
  MOAI22 U25399 ( .A1(n28030), .A2(n3180), .B1(ram[12245]), .B2(n3181), 
        .ZN(n16486) );
  MOAI22 U25400 ( .A1(n27795), .A2(n3180), .B1(ram[12246]), .B2(n3181), 
        .ZN(n16487) );
  MOAI22 U25401 ( .A1(n27560), .A2(n3180), .B1(ram[12247]), .B2(n3181), 
        .ZN(n16488) );
  MOAI22 U25402 ( .A1(n29205), .A2(n3182), .B1(ram[12248]), .B2(n3183), 
        .ZN(n16489) );
  MOAI22 U25403 ( .A1(n28970), .A2(n3182), .B1(ram[12249]), .B2(n3183), 
        .ZN(n16490) );
  MOAI22 U25404 ( .A1(n28735), .A2(n3182), .B1(ram[12250]), .B2(n3183), 
        .ZN(n16491) );
  MOAI22 U25405 ( .A1(n28500), .A2(n3182), .B1(ram[12251]), .B2(n3183), 
        .ZN(n16492) );
  MOAI22 U25406 ( .A1(n28265), .A2(n3182), .B1(ram[12252]), .B2(n3183), 
        .ZN(n16493) );
  MOAI22 U25407 ( .A1(n28030), .A2(n3182), .B1(ram[12253]), .B2(n3183), 
        .ZN(n16494) );
  MOAI22 U25408 ( .A1(n27795), .A2(n3182), .B1(ram[12254]), .B2(n3183), 
        .ZN(n16495) );
  MOAI22 U25409 ( .A1(n27560), .A2(n3182), .B1(ram[12255]), .B2(n3183), 
        .ZN(n16496) );
  MOAI22 U25410 ( .A1(n29205), .A2(n3184), .B1(ram[12256]), .B2(n3185), 
        .ZN(n16497) );
  MOAI22 U25411 ( .A1(n28970), .A2(n3184), .B1(ram[12257]), .B2(n3185), 
        .ZN(n16498) );
  MOAI22 U25412 ( .A1(n28735), .A2(n3184), .B1(ram[12258]), .B2(n3185), 
        .ZN(n16499) );
  MOAI22 U25413 ( .A1(n28500), .A2(n3184), .B1(ram[12259]), .B2(n3185), 
        .ZN(n16500) );
  MOAI22 U25414 ( .A1(n28265), .A2(n3184), .B1(ram[12260]), .B2(n3185), 
        .ZN(n16501) );
  MOAI22 U25415 ( .A1(n28030), .A2(n3184), .B1(ram[12261]), .B2(n3185), 
        .ZN(n16502) );
  MOAI22 U25416 ( .A1(n27795), .A2(n3184), .B1(ram[12262]), .B2(n3185), 
        .ZN(n16503) );
  MOAI22 U25417 ( .A1(n27560), .A2(n3184), .B1(ram[12263]), .B2(n3185), 
        .ZN(n16504) );
  MOAI22 U25418 ( .A1(n29205), .A2(n3186), .B1(ram[12264]), .B2(n3187), 
        .ZN(n16505) );
  MOAI22 U25419 ( .A1(n28970), .A2(n3186), .B1(ram[12265]), .B2(n3187), 
        .ZN(n16506) );
  MOAI22 U25420 ( .A1(n28735), .A2(n3186), .B1(ram[12266]), .B2(n3187), 
        .ZN(n16507) );
  MOAI22 U25421 ( .A1(n28500), .A2(n3186), .B1(ram[12267]), .B2(n3187), 
        .ZN(n16508) );
  MOAI22 U25422 ( .A1(n28265), .A2(n3186), .B1(ram[12268]), .B2(n3187), 
        .ZN(n16509) );
  MOAI22 U25423 ( .A1(n28030), .A2(n3186), .B1(ram[12269]), .B2(n3187), 
        .ZN(n16510) );
  MOAI22 U25424 ( .A1(n27795), .A2(n3186), .B1(ram[12270]), .B2(n3187), 
        .ZN(n16511) );
  MOAI22 U25425 ( .A1(n27560), .A2(n3186), .B1(ram[12271]), .B2(n3187), 
        .ZN(n16512) );
  MOAI22 U25426 ( .A1(n29206), .A2(n3188), .B1(ram[12272]), .B2(n3189), 
        .ZN(n16513) );
  MOAI22 U25427 ( .A1(n28971), .A2(n3188), .B1(ram[12273]), .B2(n3189), 
        .ZN(n16514) );
  MOAI22 U25428 ( .A1(n28736), .A2(n3188), .B1(ram[12274]), .B2(n3189), 
        .ZN(n16515) );
  MOAI22 U25429 ( .A1(n28501), .A2(n3188), .B1(ram[12275]), .B2(n3189), 
        .ZN(n16516) );
  MOAI22 U25430 ( .A1(n28266), .A2(n3188), .B1(ram[12276]), .B2(n3189), 
        .ZN(n16517) );
  MOAI22 U25431 ( .A1(n28031), .A2(n3188), .B1(ram[12277]), .B2(n3189), 
        .ZN(n16518) );
  MOAI22 U25432 ( .A1(n27796), .A2(n3188), .B1(ram[12278]), .B2(n3189), 
        .ZN(n16519) );
  MOAI22 U25433 ( .A1(n27561), .A2(n3188), .B1(ram[12279]), .B2(n3189), 
        .ZN(n16520) );
  MOAI22 U25434 ( .A1(n29206), .A2(n3192), .B1(ram[12288]), .B2(n3193), 
        .ZN(n16529) );
  MOAI22 U25435 ( .A1(n28971), .A2(n3192), .B1(ram[12289]), .B2(n3193), 
        .ZN(n16530) );
  MOAI22 U25436 ( .A1(n28736), .A2(n3192), .B1(ram[12290]), .B2(n3193), 
        .ZN(n16531) );
  MOAI22 U25437 ( .A1(n28501), .A2(n3192), .B1(ram[12291]), .B2(n3193), 
        .ZN(n16532) );
  MOAI22 U25438 ( .A1(n28266), .A2(n3192), .B1(ram[12292]), .B2(n3193), 
        .ZN(n16533) );
  MOAI22 U25439 ( .A1(n28031), .A2(n3192), .B1(ram[12293]), .B2(n3193), 
        .ZN(n16534) );
  MOAI22 U25440 ( .A1(n27796), .A2(n3192), .B1(ram[12294]), .B2(n3193), 
        .ZN(n16535) );
  MOAI22 U25441 ( .A1(n27561), .A2(n3192), .B1(ram[12295]), .B2(n3193), 
        .ZN(n16536) );
  MOAI22 U25442 ( .A1(n29206), .A2(n3195), .B1(ram[12296]), .B2(n3196), 
        .ZN(n16537) );
  MOAI22 U25443 ( .A1(n28971), .A2(n3195), .B1(ram[12297]), .B2(n3196), 
        .ZN(n16538) );
  MOAI22 U25444 ( .A1(n28736), .A2(n3195), .B1(ram[12298]), .B2(n3196), 
        .ZN(n16539) );
  MOAI22 U25445 ( .A1(n28501), .A2(n3195), .B1(ram[12299]), .B2(n3196), 
        .ZN(n16540) );
  MOAI22 U25446 ( .A1(n28266), .A2(n3195), .B1(ram[12300]), .B2(n3196), 
        .ZN(n16541) );
  MOAI22 U25447 ( .A1(n28031), .A2(n3195), .B1(ram[12301]), .B2(n3196), 
        .ZN(n16542) );
  MOAI22 U25448 ( .A1(n27796), .A2(n3195), .B1(ram[12302]), .B2(n3196), 
        .ZN(n16543) );
  MOAI22 U25449 ( .A1(n27561), .A2(n3195), .B1(ram[12303]), .B2(n3196), 
        .ZN(n16544) );
  MOAI22 U25450 ( .A1(n29206), .A2(n3197), .B1(ram[12304]), .B2(n3198), 
        .ZN(n16545) );
  MOAI22 U25451 ( .A1(n28971), .A2(n3197), .B1(ram[12305]), .B2(n3198), 
        .ZN(n16546) );
  MOAI22 U25452 ( .A1(n28736), .A2(n3197), .B1(ram[12306]), .B2(n3198), 
        .ZN(n16547) );
  MOAI22 U25453 ( .A1(n28501), .A2(n3197), .B1(ram[12307]), .B2(n3198), 
        .ZN(n16548) );
  MOAI22 U25454 ( .A1(n28266), .A2(n3197), .B1(ram[12308]), .B2(n3198), 
        .ZN(n16549) );
  MOAI22 U25455 ( .A1(n28031), .A2(n3197), .B1(ram[12309]), .B2(n3198), 
        .ZN(n16550) );
  MOAI22 U25456 ( .A1(n27796), .A2(n3197), .B1(ram[12310]), .B2(n3198), 
        .ZN(n16551) );
  MOAI22 U25457 ( .A1(n27561), .A2(n3197), .B1(ram[12311]), .B2(n3198), 
        .ZN(n16552) );
  MOAI22 U25458 ( .A1(n29206), .A2(n3199), .B1(ram[12312]), .B2(n3200), 
        .ZN(n16553) );
  MOAI22 U25459 ( .A1(n28971), .A2(n3199), .B1(ram[12313]), .B2(n3200), 
        .ZN(n16554) );
  MOAI22 U25460 ( .A1(n28736), .A2(n3199), .B1(ram[12314]), .B2(n3200), 
        .ZN(n16555) );
  MOAI22 U25461 ( .A1(n28501), .A2(n3199), .B1(ram[12315]), .B2(n3200), 
        .ZN(n16556) );
  MOAI22 U25462 ( .A1(n28266), .A2(n3199), .B1(ram[12316]), .B2(n3200), 
        .ZN(n16557) );
  MOAI22 U25463 ( .A1(n28031), .A2(n3199), .B1(ram[12317]), .B2(n3200), 
        .ZN(n16558) );
  MOAI22 U25464 ( .A1(n27796), .A2(n3199), .B1(ram[12318]), .B2(n3200), 
        .ZN(n16559) );
  MOAI22 U25465 ( .A1(n27561), .A2(n3199), .B1(ram[12319]), .B2(n3200), 
        .ZN(n16560) );
  MOAI22 U25466 ( .A1(n29206), .A2(n3201), .B1(ram[12320]), .B2(n3202), 
        .ZN(n16561) );
  MOAI22 U25467 ( .A1(n28971), .A2(n3201), .B1(ram[12321]), .B2(n3202), 
        .ZN(n16562) );
  MOAI22 U25468 ( .A1(n28736), .A2(n3201), .B1(ram[12322]), .B2(n3202), 
        .ZN(n16563) );
  MOAI22 U25469 ( .A1(n28501), .A2(n3201), .B1(ram[12323]), .B2(n3202), 
        .ZN(n16564) );
  MOAI22 U25470 ( .A1(n28266), .A2(n3201), .B1(ram[12324]), .B2(n3202), 
        .ZN(n16565) );
  MOAI22 U25471 ( .A1(n28031), .A2(n3201), .B1(ram[12325]), .B2(n3202), 
        .ZN(n16566) );
  MOAI22 U25472 ( .A1(n27796), .A2(n3201), .B1(ram[12326]), .B2(n3202), 
        .ZN(n16567) );
  MOAI22 U25473 ( .A1(n27561), .A2(n3201), .B1(ram[12327]), .B2(n3202), 
        .ZN(n16568) );
  MOAI22 U25474 ( .A1(n29206), .A2(n3203), .B1(ram[12328]), .B2(n3204), 
        .ZN(n16569) );
  MOAI22 U25475 ( .A1(n28971), .A2(n3203), .B1(ram[12329]), .B2(n3204), 
        .ZN(n16570) );
  MOAI22 U25476 ( .A1(n28736), .A2(n3203), .B1(ram[12330]), .B2(n3204), 
        .ZN(n16571) );
  MOAI22 U25477 ( .A1(n28501), .A2(n3203), .B1(ram[12331]), .B2(n3204), 
        .ZN(n16572) );
  MOAI22 U25478 ( .A1(n28266), .A2(n3203), .B1(ram[12332]), .B2(n3204), 
        .ZN(n16573) );
  MOAI22 U25479 ( .A1(n28031), .A2(n3203), .B1(ram[12333]), .B2(n3204), 
        .ZN(n16574) );
  MOAI22 U25480 ( .A1(n27796), .A2(n3203), .B1(ram[12334]), .B2(n3204), 
        .ZN(n16575) );
  MOAI22 U25481 ( .A1(n27561), .A2(n3203), .B1(ram[12335]), .B2(n3204), 
        .ZN(n16576) );
  MOAI22 U25482 ( .A1(n29206), .A2(n3205), .B1(ram[12336]), .B2(n3206), 
        .ZN(n16577) );
  MOAI22 U25483 ( .A1(n28971), .A2(n3205), .B1(ram[12337]), .B2(n3206), 
        .ZN(n16578) );
  MOAI22 U25484 ( .A1(n28736), .A2(n3205), .B1(ram[12338]), .B2(n3206), 
        .ZN(n16579) );
  MOAI22 U25485 ( .A1(n28501), .A2(n3205), .B1(ram[12339]), .B2(n3206), 
        .ZN(n16580) );
  MOAI22 U25486 ( .A1(n28266), .A2(n3205), .B1(ram[12340]), .B2(n3206), 
        .ZN(n16581) );
  MOAI22 U25487 ( .A1(n28031), .A2(n3205), .B1(ram[12341]), .B2(n3206), 
        .ZN(n16582) );
  MOAI22 U25488 ( .A1(n27796), .A2(n3205), .B1(ram[12342]), .B2(n3206), 
        .ZN(n16583) );
  MOAI22 U25489 ( .A1(n27561), .A2(n3205), .B1(ram[12343]), .B2(n3206), 
        .ZN(n16584) );
  MOAI22 U25490 ( .A1(n29206), .A2(n3207), .B1(ram[12344]), .B2(n3208), 
        .ZN(n16585) );
  MOAI22 U25491 ( .A1(n28971), .A2(n3207), .B1(ram[12345]), .B2(n3208), 
        .ZN(n16586) );
  MOAI22 U25492 ( .A1(n28736), .A2(n3207), .B1(ram[12346]), .B2(n3208), 
        .ZN(n16587) );
  MOAI22 U25493 ( .A1(n28501), .A2(n3207), .B1(ram[12347]), .B2(n3208), 
        .ZN(n16588) );
  MOAI22 U25494 ( .A1(n28266), .A2(n3207), .B1(ram[12348]), .B2(n3208), 
        .ZN(n16589) );
  MOAI22 U25495 ( .A1(n28031), .A2(n3207), .B1(ram[12349]), .B2(n3208), 
        .ZN(n16590) );
  MOAI22 U25496 ( .A1(n27796), .A2(n3207), .B1(ram[12350]), .B2(n3208), 
        .ZN(n16591) );
  MOAI22 U25497 ( .A1(n27561), .A2(n3207), .B1(ram[12351]), .B2(n3208), 
        .ZN(n16592) );
  MOAI22 U25498 ( .A1(n29206), .A2(n3209), .B1(ram[12352]), .B2(n3210), 
        .ZN(n16593) );
  MOAI22 U25499 ( .A1(n28971), .A2(n3209), .B1(ram[12353]), .B2(n3210), 
        .ZN(n16594) );
  MOAI22 U25500 ( .A1(n28736), .A2(n3209), .B1(ram[12354]), .B2(n3210), 
        .ZN(n16595) );
  MOAI22 U25501 ( .A1(n28501), .A2(n3209), .B1(ram[12355]), .B2(n3210), 
        .ZN(n16596) );
  MOAI22 U25502 ( .A1(n28266), .A2(n3209), .B1(ram[12356]), .B2(n3210), 
        .ZN(n16597) );
  MOAI22 U25503 ( .A1(n28031), .A2(n3209), .B1(ram[12357]), .B2(n3210), 
        .ZN(n16598) );
  MOAI22 U25504 ( .A1(n27796), .A2(n3209), .B1(ram[12358]), .B2(n3210), 
        .ZN(n16599) );
  MOAI22 U25505 ( .A1(n27561), .A2(n3209), .B1(ram[12359]), .B2(n3210), 
        .ZN(n16600) );
  MOAI22 U25506 ( .A1(n29206), .A2(n3211), .B1(ram[12360]), .B2(n3212), 
        .ZN(n16601) );
  MOAI22 U25507 ( .A1(n28971), .A2(n3211), .B1(ram[12361]), .B2(n3212), 
        .ZN(n16602) );
  MOAI22 U25508 ( .A1(n28736), .A2(n3211), .B1(ram[12362]), .B2(n3212), 
        .ZN(n16603) );
  MOAI22 U25509 ( .A1(n28501), .A2(n3211), .B1(ram[12363]), .B2(n3212), 
        .ZN(n16604) );
  MOAI22 U25510 ( .A1(n28266), .A2(n3211), .B1(ram[12364]), .B2(n3212), 
        .ZN(n16605) );
  MOAI22 U25511 ( .A1(n28031), .A2(n3211), .B1(ram[12365]), .B2(n3212), 
        .ZN(n16606) );
  MOAI22 U25512 ( .A1(n27796), .A2(n3211), .B1(ram[12366]), .B2(n3212), 
        .ZN(n16607) );
  MOAI22 U25513 ( .A1(n27561), .A2(n3211), .B1(ram[12367]), .B2(n3212), 
        .ZN(n16608) );
  MOAI22 U25514 ( .A1(n29206), .A2(n3213), .B1(ram[12368]), .B2(n3214), 
        .ZN(n16609) );
  MOAI22 U25515 ( .A1(n28971), .A2(n3213), .B1(ram[12369]), .B2(n3214), 
        .ZN(n16610) );
  MOAI22 U25516 ( .A1(n28736), .A2(n3213), .B1(ram[12370]), .B2(n3214), 
        .ZN(n16611) );
  MOAI22 U25517 ( .A1(n28501), .A2(n3213), .B1(ram[12371]), .B2(n3214), 
        .ZN(n16612) );
  MOAI22 U25518 ( .A1(n28266), .A2(n3213), .B1(ram[12372]), .B2(n3214), 
        .ZN(n16613) );
  MOAI22 U25519 ( .A1(n28031), .A2(n3213), .B1(ram[12373]), .B2(n3214), 
        .ZN(n16614) );
  MOAI22 U25520 ( .A1(n27796), .A2(n3213), .B1(ram[12374]), .B2(n3214), 
        .ZN(n16615) );
  MOAI22 U25521 ( .A1(n27561), .A2(n3213), .B1(ram[12375]), .B2(n3214), 
        .ZN(n16616) );
  MOAI22 U25522 ( .A1(n29207), .A2(n3215), .B1(ram[12376]), .B2(n3216), 
        .ZN(n16617) );
  MOAI22 U25523 ( .A1(n28972), .A2(n3215), .B1(ram[12377]), .B2(n3216), 
        .ZN(n16618) );
  MOAI22 U25524 ( .A1(n28737), .A2(n3215), .B1(ram[12378]), .B2(n3216), 
        .ZN(n16619) );
  MOAI22 U25525 ( .A1(n28502), .A2(n3215), .B1(ram[12379]), .B2(n3216), 
        .ZN(n16620) );
  MOAI22 U25526 ( .A1(n28267), .A2(n3215), .B1(ram[12380]), .B2(n3216), 
        .ZN(n16621) );
  MOAI22 U25527 ( .A1(n28032), .A2(n3215), .B1(ram[12381]), .B2(n3216), 
        .ZN(n16622) );
  MOAI22 U25528 ( .A1(n27797), .A2(n3215), .B1(ram[12382]), .B2(n3216), 
        .ZN(n16623) );
  MOAI22 U25529 ( .A1(n27562), .A2(n3215), .B1(ram[12383]), .B2(n3216), 
        .ZN(n16624) );
  MOAI22 U25530 ( .A1(n29207), .A2(n3217), .B1(ram[12384]), .B2(n3218), 
        .ZN(n16625) );
  MOAI22 U25531 ( .A1(n28972), .A2(n3217), .B1(ram[12385]), .B2(n3218), 
        .ZN(n16626) );
  MOAI22 U25532 ( .A1(n28737), .A2(n3217), .B1(ram[12386]), .B2(n3218), 
        .ZN(n16627) );
  MOAI22 U25533 ( .A1(n28502), .A2(n3217), .B1(ram[12387]), .B2(n3218), 
        .ZN(n16628) );
  MOAI22 U25534 ( .A1(n28267), .A2(n3217), .B1(ram[12388]), .B2(n3218), 
        .ZN(n16629) );
  MOAI22 U25535 ( .A1(n28032), .A2(n3217), .B1(ram[12389]), .B2(n3218), 
        .ZN(n16630) );
  MOAI22 U25536 ( .A1(n27797), .A2(n3217), .B1(ram[12390]), .B2(n3218), 
        .ZN(n16631) );
  MOAI22 U25537 ( .A1(n27562), .A2(n3217), .B1(ram[12391]), .B2(n3218), 
        .ZN(n16632) );
  MOAI22 U25538 ( .A1(n29207), .A2(n3219), .B1(ram[12392]), .B2(n3220), 
        .ZN(n16633) );
  MOAI22 U25539 ( .A1(n28972), .A2(n3219), .B1(ram[12393]), .B2(n3220), 
        .ZN(n16634) );
  MOAI22 U25540 ( .A1(n28737), .A2(n3219), .B1(ram[12394]), .B2(n3220), 
        .ZN(n16635) );
  MOAI22 U25541 ( .A1(n28502), .A2(n3219), .B1(ram[12395]), .B2(n3220), 
        .ZN(n16636) );
  MOAI22 U25542 ( .A1(n28267), .A2(n3219), .B1(ram[12396]), .B2(n3220), 
        .ZN(n16637) );
  MOAI22 U25543 ( .A1(n28032), .A2(n3219), .B1(ram[12397]), .B2(n3220), 
        .ZN(n16638) );
  MOAI22 U25544 ( .A1(n27797), .A2(n3219), .B1(ram[12398]), .B2(n3220), 
        .ZN(n16639) );
  MOAI22 U25545 ( .A1(n27562), .A2(n3219), .B1(ram[12399]), .B2(n3220), 
        .ZN(n16640) );
  MOAI22 U25546 ( .A1(n29207), .A2(n3221), .B1(ram[12400]), .B2(n3222), 
        .ZN(n16641) );
  MOAI22 U25547 ( .A1(n28972), .A2(n3221), .B1(ram[12401]), .B2(n3222), 
        .ZN(n16642) );
  MOAI22 U25548 ( .A1(n28737), .A2(n3221), .B1(ram[12402]), .B2(n3222), 
        .ZN(n16643) );
  MOAI22 U25549 ( .A1(n28502), .A2(n3221), .B1(ram[12403]), .B2(n3222), 
        .ZN(n16644) );
  MOAI22 U25550 ( .A1(n28267), .A2(n3221), .B1(ram[12404]), .B2(n3222), 
        .ZN(n16645) );
  MOAI22 U25551 ( .A1(n28032), .A2(n3221), .B1(ram[12405]), .B2(n3222), 
        .ZN(n16646) );
  MOAI22 U25552 ( .A1(n27797), .A2(n3221), .B1(ram[12406]), .B2(n3222), 
        .ZN(n16647) );
  MOAI22 U25553 ( .A1(n27562), .A2(n3221), .B1(ram[12407]), .B2(n3222), 
        .ZN(n16648) );
  MOAI22 U25554 ( .A1(n29207), .A2(n3223), .B1(ram[12408]), .B2(n3224), 
        .ZN(n16649) );
  MOAI22 U25555 ( .A1(n28972), .A2(n3223), .B1(ram[12409]), .B2(n3224), 
        .ZN(n16650) );
  MOAI22 U25556 ( .A1(n28737), .A2(n3223), .B1(ram[12410]), .B2(n3224), 
        .ZN(n16651) );
  MOAI22 U25557 ( .A1(n28502), .A2(n3223), .B1(ram[12411]), .B2(n3224), 
        .ZN(n16652) );
  MOAI22 U25558 ( .A1(n28267), .A2(n3223), .B1(ram[12412]), .B2(n3224), 
        .ZN(n16653) );
  MOAI22 U25559 ( .A1(n28032), .A2(n3223), .B1(ram[12413]), .B2(n3224), 
        .ZN(n16654) );
  MOAI22 U25560 ( .A1(n27797), .A2(n3223), .B1(ram[12414]), .B2(n3224), 
        .ZN(n16655) );
  MOAI22 U25561 ( .A1(n27562), .A2(n3223), .B1(ram[12415]), .B2(n3224), 
        .ZN(n16656) );
  MOAI22 U25562 ( .A1(n29207), .A2(n3225), .B1(ram[12416]), .B2(n3226), 
        .ZN(n16657) );
  MOAI22 U25563 ( .A1(n28972), .A2(n3225), .B1(ram[12417]), .B2(n3226), 
        .ZN(n16658) );
  MOAI22 U25564 ( .A1(n28737), .A2(n3225), .B1(ram[12418]), .B2(n3226), 
        .ZN(n16659) );
  MOAI22 U25565 ( .A1(n28502), .A2(n3225), .B1(ram[12419]), .B2(n3226), 
        .ZN(n16660) );
  MOAI22 U25566 ( .A1(n28267), .A2(n3225), .B1(ram[12420]), .B2(n3226), 
        .ZN(n16661) );
  MOAI22 U25567 ( .A1(n28032), .A2(n3225), .B1(ram[12421]), .B2(n3226), 
        .ZN(n16662) );
  MOAI22 U25568 ( .A1(n27797), .A2(n3225), .B1(ram[12422]), .B2(n3226), 
        .ZN(n16663) );
  MOAI22 U25569 ( .A1(n27562), .A2(n3225), .B1(ram[12423]), .B2(n3226), 
        .ZN(n16664) );
  MOAI22 U25570 ( .A1(n29207), .A2(n3227), .B1(ram[12424]), .B2(n3228), 
        .ZN(n16665) );
  MOAI22 U25571 ( .A1(n28972), .A2(n3227), .B1(ram[12425]), .B2(n3228), 
        .ZN(n16666) );
  MOAI22 U25572 ( .A1(n28737), .A2(n3227), .B1(ram[12426]), .B2(n3228), 
        .ZN(n16667) );
  MOAI22 U25573 ( .A1(n28502), .A2(n3227), .B1(ram[12427]), .B2(n3228), 
        .ZN(n16668) );
  MOAI22 U25574 ( .A1(n28267), .A2(n3227), .B1(ram[12428]), .B2(n3228), 
        .ZN(n16669) );
  MOAI22 U25575 ( .A1(n28032), .A2(n3227), .B1(ram[12429]), .B2(n3228), 
        .ZN(n16670) );
  MOAI22 U25576 ( .A1(n27797), .A2(n3227), .B1(ram[12430]), .B2(n3228), 
        .ZN(n16671) );
  MOAI22 U25577 ( .A1(n27562), .A2(n3227), .B1(ram[12431]), .B2(n3228), 
        .ZN(n16672) );
  MOAI22 U25578 ( .A1(n29207), .A2(n3229), .B1(ram[12432]), .B2(n3230), 
        .ZN(n16673) );
  MOAI22 U25579 ( .A1(n28972), .A2(n3229), .B1(ram[12433]), .B2(n3230), 
        .ZN(n16674) );
  MOAI22 U25580 ( .A1(n28737), .A2(n3229), .B1(ram[12434]), .B2(n3230), 
        .ZN(n16675) );
  MOAI22 U25581 ( .A1(n28502), .A2(n3229), .B1(ram[12435]), .B2(n3230), 
        .ZN(n16676) );
  MOAI22 U25582 ( .A1(n28267), .A2(n3229), .B1(ram[12436]), .B2(n3230), 
        .ZN(n16677) );
  MOAI22 U25583 ( .A1(n28032), .A2(n3229), .B1(ram[12437]), .B2(n3230), 
        .ZN(n16678) );
  MOAI22 U25584 ( .A1(n27797), .A2(n3229), .B1(ram[12438]), .B2(n3230), 
        .ZN(n16679) );
  MOAI22 U25585 ( .A1(n27562), .A2(n3229), .B1(ram[12439]), .B2(n3230), 
        .ZN(n16680) );
  MOAI22 U25586 ( .A1(n29207), .A2(n3231), .B1(ram[12440]), .B2(n3232), 
        .ZN(n16681) );
  MOAI22 U25587 ( .A1(n28972), .A2(n3231), .B1(ram[12441]), .B2(n3232), 
        .ZN(n16682) );
  MOAI22 U25588 ( .A1(n28737), .A2(n3231), .B1(ram[12442]), .B2(n3232), 
        .ZN(n16683) );
  MOAI22 U25589 ( .A1(n28502), .A2(n3231), .B1(ram[12443]), .B2(n3232), 
        .ZN(n16684) );
  MOAI22 U25590 ( .A1(n28267), .A2(n3231), .B1(ram[12444]), .B2(n3232), 
        .ZN(n16685) );
  MOAI22 U25591 ( .A1(n28032), .A2(n3231), .B1(ram[12445]), .B2(n3232), 
        .ZN(n16686) );
  MOAI22 U25592 ( .A1(n27797), .A2(n3231), .B1(ram[12446]), .B2(n3232), 
        .ZN(n16687) );
  MOAI22 U25593 ( .A1(n27562), .A2(n3231), .B1(ram[12447]), .B2(n3232), 
        .ZN(n16688) );
  MOAI22 U25594 ( .A1(n29207), .A2(n3233), .B1(ram[12448]), .B2(n3234), 
        .ZN(n16689) );
  MOAI22 U25595 ( .A1(n28972), .A2(n3233), .B1(ram[12449]), .B2(n3234), 
        .ZN(n16690) );
  MOAI22 U25596 ( .A1(n28737), .A2(n3233), .B1(ram[12450]), .B2(n3234), 
        .ZN(n16691) );
  MOAI22 U25597 ( .A1(n28502), .A2(n3233), .B1(ram[12451]), .B2(n3234), 
        .ZN(n16692) );
  MOAI22 U25598 ( .A1(n28267), .A2(n3233), .B1(ram[12452]), .B2(n3234), 
        .ZN(n16693) );
  MOAI22 U25599 ( .A1(n28032), .A2(n3233), .B1(ram[12453]), .B2(n3234), 
        .ZN(n16694) );
  MOAI22 U25600 ( .A1(n27797), .A2(n3233), .B1(ram[12454]), .B2(n3234), 
        .ZN(n16695) );
  MOAI22 U25601 ( .A1(n27562), .A2(n3233), .B1(ram[12455]), .B2(n3234), 
        .ZN(n16696) );
  MOAI22 U25602 ( .A1(n29207), .A2(n3235), .B1(ram[12456]), .B2(n3236), 
        .ZN(n16697) );
  MOAI22 U25603 ( .A1(n28972), .A2(n3235), .B1(ram[12457]), .B2(n3236), 
        .ZN(n16698) );
  MOAI22 U25604 ( .A1(n28737), .A2(n3235), .B1(ram[12458]), .B2(n3236), 
        .ZN(n16699) );
  MOAI22 U25605 ( .A1(n28502), .A2(n3235), .B1(ram[12459]), .B2(n3236), 
        .ZN(n16700) );
  MOAI22 U25606 ( .A1(n28267), .A2(n3235), .B1(ram[12460]), .B2(n3236), 
        .ZN(n16701) );
  MOAI22 U25607 ( .A1(n28032), .A2(n3235), .B1(ram[12461]), .B2(n3236), 
        .ZN(n16702) );
  MOAI22 U25608 ( .A1(n27797), .A2(n3235), .B1(ram[12462]), .B2(n3236), 
        .ZN(n16703) );
  MOAI22 U25609 ( .A1(n27562), .A2(n3235), .B1(ram[12463]), .B2(n3236), 
        .ZN(n16704) );
  MOAI22 U25610 ( .A1(n29207), .A2(n3237), .B1(ram[12464]), .B2(n3238), 
        .ZN(n16705) );
  MOAI22 U25611 ( .A1(n28972), .A2(n3237), .B1(ram[12465]), .B2(n3238), 
        .ZN(n16706) );
  MOAI22 U25612 ( .A1(n28737), .A2(n3237), .B1(ram[12466]), .B2(n3238), 
        .ZN(n16707) );
  MOAI22 U25613 ( .A1(n28502), .A2(n3237), .B1(ram[12467]), .B2(n3238), 
        .ZN(n16708) );
  MOAI22 U25614 ( .A1(n28267), .A2(n3237), .B1(ram[12468]), .B2(n3238), 
        .ZN(n16709) );
  MOAI22 U25615 ( .A1(n28032), .A2(n3237), .B1(ram[12469]), .B2(n3238), 
        .ZN(n16710) );
  MOAI22 U25616 ( .A1(n27797), .A2(n3237), .B1(ram[12470]), .B2(n3238), 
        .ZN(n16711) );
  MOAI22 U25617 ( .A1(n27562), .A2(n3237), .B1(ram[12471]), .B2(n3238), 
        .ZN(n16712) );
  MOAI22 U25618 ( .A1(n29207), .A2(n3239), .B1(ram[12472]), .B2(n3240), 
        .ZN(n16713) );
  MOAI22 U25619 ( .A1(n28972), .A2(n3239), .B1(ram[12473]), .B2(n3240), 
        .ZN(n16714) );
  MOAI22 U25620 ( .A1(n28737), .A2(n3239), .B1(ram[12474]), .B2(n3240), 
        .ZN(n16715) );
  MOAI22 U25621 ( .A1(n28502), .A2(n3239), .B1(ram[12475]), .B2(n3240), 
        .ZN(n16716) );
  MOAI22 U25622 ( .A1(n28267), .A2(n3239), .B1(ram[12476]), .B2(n3240), 
        .ZN(n16717) );
  MOAI22 U25623 ( .A1(n28032), .A2(n3239), .B1(ram[12477]), .B2(n3240), 
        .ZN(n16718) );
  MOAI22 U25624 ( .A1(n27797), .A2(n3239), .B1(ram[12478]), .B2(n3240), 
        .ZN(n16719) );
  MOAI22 U25625 ( .A1(n27562), .A2(n3239), .B1(ram[12479]), .B2(n3240), 
        .ZN(n16720) );
  MOAI22 U25626 ( .A1(n29208), .A2(n3241), .B1(ram[12480]), .B2(n3242), 
        .ZN(n16721) );
  MOAI22 U25627 ( .A1(n28973), .A2(n3241), .B1(ram[12481]), .B2(n3242), 
        .ZN(n16722) );
  MOAI22 U25628 ( .A1(n28738), .A2(n3241), .B1(ram[12482]), .B2(n3242), 
        .ZN(n16723) );
  MOAI22 U25629 ( .A1(n28503), .A2(n3241), .B1(ram[12483]), .B2(n3242), 
        .ZN(n16724) );
  MOAI22 U25630 ( .A1(n28268), .A2(n3241), .B1(ram[12484]), .B2(n3242), 
        .ZN(n16725) );
  MOAI22 U25631 ( .A1(n28033), .A2(n3241), .B1(ram[12485]), .B2(n3242), 
        .ZN(n16726) );
  MOAI22 U25632 ( .A1(n27798), .A2(n3241), .B1(ram[12486]), .B2(n3242), 
        .ZN(n16727) );
  MOAI22 U25633 ( .A1(n27563), .A2(n3241), .B1(ram[12487]), .B2(n3242), 
        .ZN(n16728) );
  MOAI22 U25634 ( .A1(n29208), .A2(n3243), .B1(ram[12488]), .B2(n3244), 
        .ZN(n16729) );
  MOAI22 U25635 ( .A1(n28973), .A2(n3243), .B1(ram[12489]), .B2(n3244), 
        .ZN(n16730) );
  MOAI22 U25636 ( .A1(n28738), .A2(n3243), .B1(ram[12490]), .B2(n3244), 
        .ZN(n16731) );
  MOAI22 U25637 ( .A1(n28503), .A2(n3243), .B1(ram[12491]), .B2(n3244), 
        .ZN(n16732) );
  MOAI22 U25638 ( .A1(n28268), .A2(n3243), .B1(ram[12492]), .B2(n3244), 
        .ZN(n16733) );
  MOAI22 U25639 ( .A1(n28033), .A2(n3243), .B1(ram[12493]), .B2(n3244), 
        .ZN(n16734) );
  MOAI22 U25640 ( .A1(n27798), .A2(n3243), .B1(ram[12494]), .B2(n3244), 
        .ZN(n16735) );
  MOAI22 U25641 ( .A1(n27563), .A2(n3243), .B1(ram[12495]), .B2(n3244), 
        .ZN(n16736) );
  MOAI22 U25642 ( .A1(n29208), .A2(n3245), .B1(ram[12496]), .B2(n3246), 
        .ZN(n16737) );
  MOAI22 U25643 ( .A1(n28973), .A2(n3245), .B1(ram[12497]), .B2(n3246), 
        .ZN(n16738) );
  MOAI22 U25644 ( .A1(n28738), .A2(n3245), .B1(ram[12498]), .B2(n3246), 
        .ZN(n16739) );
  MOAI22 U25645 ( .A1(n28503), .A2(n3245), .B1(ram[12499]), .B2(n3246), 
        .ZN(n16740) );
  MOAI22 U25646 ( .A1(n28268), .A2(n3245), .B1(ram[12500]), .B2(n3246), 
        .ZN(n16741) );
  MOAI22 U25647 ( .A1(n28033), .A2(n3245), .B1(ram[12501]), .B2(n3246), 
        .ZN(n16742) );
  MOAI22 U25648 ( .A1(n27798), .A2(n3245), .B1(ram[12502]), .B2(n3246), 
        .ZN(n16743) );
  MOAI22 U25649 ( .A1(n27563), .A2(n3245), .B1(ram[12503]), .B2(n3246), 
        .ZN(n16744) );
  MOAI22 U25650 ( .A1(n29208), .A2(n3247), .B1(ram[12504]), .B2(n3248), 
        .ZN(n16745) );
  MOAI22 U25651 ( .A1(n28973), .A2(n3247), .B1(ram[12505]), .B2(n3248), 
        .ZN(n16746) );
  MOAI22 U25652 ( .A1(n28738), .A2(n3247), .B1(ram[12506]), .B2(n3248), 
        .ZN(n16747) );
  MOAI22 U25653 ( .A1(n28503), .A2(n3247), .B1(ram[12507]), .B2(n3248), 
        .ZN(n16748) );
  MOAI22 U25654 ( .A1(n28268), .A2(n3247), .B1(ram[12508]), .B2(n3248), 
        .ZN(n16749) );
  MOAI22 U25655 ( .A1(n28033), .A2(n3247), .B1(ram[12509]), .B2(n3248), 
        .ZN(n16750) );
  MOAI22 U25656 ( .A1(n27798), .A2(n3247), .B1(ram[12510]), .B2(n3248), 
        .ZN(n16751) );
  MOAI22 U25657 ( .A1(n27563), .A2(n3247), .B1(ram[12511]), .B2(n3248), 
        .ZN(n16752) );
  MOAI22 U25658 ( .A1(n29208), .A2(n3249), .B1(ram[12512]), .B2(n3250), 
        .ZN(n16753) );
  MOAI22 U25659 ( .A1(n28973), .A2(n3249), .B1(ram[12513]), .B2(n3250), 
        .ZN(n16754) );
  MOAI22 U25660 ( .A1(n28738), .A2(n3249), .B1(ram[12514]), .B2(n3250), 
        .ZN(n16755) );
  MOAI22 U25661 ( .A1(n28503), .A2(n3249), .B1(ram[12515]), .B2(n3250), 
        .ZN(n16756) );
  MOAI22 U25662 ( .A1(n28268), .A2(n3249), .B1(ram[12516]), .B2(n3250), 
        .ZN(n16757) );
  MOAI22 U25663 ( .A1(n28033), .A2(n3249), .B1(ram[12517]), .B2(n3250), 
        .ZN(n16758) );
  MOAI22 U25664 ( .A1(n27798), .A2(n3249), .B1(ram[12518]), .B2(n3250), 
        .ZN(n16759) );
  MOAI22 U25665 ( .A1(n27563), .A2(n3249), .B1(ram[12519]), .B2(n3250), 
        .ZN(n16760) );
  MOAI22 U25666 ( .A1(n29208), .A2(n3251), .B1(ram[12520]), .B2(n3252), 
        .ZN(n16761) );
  MOAI22 U25667 ( .A1(n28973), .A2(n3251), .B1(ram[12521]), .B2(n3252), 
        .ZN(n16762) );
  MOAI22 U25668 ( .A1(n28738), .A2(n3251), .B1(ram[12522]), .B2(n3252), 
        .ZN(n16763) );
  MOAI22 U25669 ( .A1(n28503), .A2(n3251), .B1(ram[12523]), .B2(n3252), 
        .ZN(n16764) );
  MOAI22 U25670 ( .A1(n28268), .A2(n3251), .B1(ram[12524]), .B2(n3252), 
        .ZN(n16765) );
  MOAI22 U25671 ( .A1(n28033), .A2(n3251), .B1(ram[12525]), .B2(n3252), 
        .ZN(n16766) );
  MOAI22 U25672 ( .A1(n27798), .A2(n3251), .B1(ram[12526]), .B2(n3252), 
        .ZN(n16767) );
  MOAI22 U25673 ( .A1(n27563), .A2(n3251), .B1(ram[12527]), .B2(n3252), 
        .ZN(n16768) );
  MOAI22 U25674 ( .A1(n29208), .A2(n3253), .B1(ram[12528]), .B2(n3254), 
        .ZN(n16769) );
  MOAI22 U25675 ( .A1(n28973), .A2(n3253), .B1(ram[12529]), .B2(n3254), 
        .ZN(n16770) );
  MOAI22 U25676 ( .A1(n28738), .A2(n3253), .B1(ram[12530]), .B2(n3254), 
        .ZN(n16771) );
  MOAI22 U25677 ( .A1(n28503), .A2(n3253), .B1(ram[12531]), .B2(n3254), 
        .ZN(n16772) );
  MOAI22 U25678 ( .A1(n28268), .A2(n3253), .B1(ram[12532]), .B2(n3254), 
        .ZN(n16773) );
  MOAI22 U25679 ( .A1(n28033), .A2(n3253), .B1(ram[12533]), .B2(n3254), 
        .ZN(n16774) );
  MOAI22 U25680 ( .A1(n27798), .A2(n3253), .B1(ram[12534]), .B2(n3254), 
        .ZN(n16775) );
  MOAI22 U25681 ( .A1(n27563), .A2(n3253), .B1(ram[12535]), .B2(n3254), 
        .ZN(n16776) );
  MOAI22 U25682 ( .A1(n29208), .A2(n3255), .B1(ram[12536]), .B2(n3256), 
        .ZN(n16777) );
  MOAI22 U25683 ( .A1(n28973), .A2(n3255), .B1(ram[12537]), .B2(n3256), 
        .ZN(n16778) );
  MOAI22 U25684 ( .A1(n28738), .A2(n3255), .B1(ram[12538]), .B2(n3256), 
        .ZN(n16779) );
  MOAI22 U25685 ( .A1(n28503), .A2(n3255), .B1(ram[12539]), .B2(n3256), 
        .ZN(n16780) );
  MOAI22 U25686 ( .A1(n28268), .A2(n3255), .B1(ram[12540]), .B2(n3256), 
        .ZN(n16781) );
  MOAI22 U25687 ( .A1(n28033), .A2(n3255), .B1(ram[12541]), .B2(n3256), 
        .ZN(n16782) );
  MOAI22 U25688 ( .A1(n27798), .A2(n3255), .B1(ram[12542]), .B2(n3256), 
        .ZN(n16783) );
  MOAI22 U25689 ( .A1(n27563), .A2(n3255), .B1(ram[12543]), .B2(n3256), 
        .ZN(n16784) );
  MOAI22 U25690 ( .A1(n29208), .A2(n3257), .B1(ram[12544]), .B2(n3258), 
        .ZN(n16785) );
  MOAI22 U25691 ( .A1(n28973), .A2(n3257), .B1(ram[12545]), .B2(n3258), 
        .ZN(n16786) );
  MOAI22 U25692 ( .A1(n28738), .A2(n3257), .B1(ram[12546]), .B2(n3258), 
        .ZN(n16787) );
  MOAI22 U25693 ( .A1(n28503), .A2(n3257), .B1(ram[12547]), .B2(n3258), 
        .ZN(n16788) );
  MOAI22 U25694 ( .A1(n28268), .A2(n3257), .B1(ram[12548]), .B2(n3258), 
        .ZN(n16789) );
  MOAI22 U25695 ( .A1(n28033), .A2(n3257), .B1(ram[12549]), .B2(n3258), 
        .ZN(n16790) );
  MOAI22 U25696 ( .A1(n27798), .A2(n3257), .B1(ram[12550]), .B2(n3258), 
        .ZN(n16791) );
  MOAI22 U25697 ( .A1(n27563), .A2(n3257), .B1(ram[12551]), .B2(n3258), 
        .ZN(n16792) );
  MOAI22 U25698 ( .A1(n29208), .A2(n3259), .B1(ram[12552]), .B2(n3260), 
        .ZN(n16793) );
  MOAI22 U25699 ( .A1(n28973), .A2(n3259), .B1(ram[12553]), .B2(n3260), 
        .ZN(n16794) );
  MOAI22 U25700 ( .A1(n28738), .A2(n3259), .B1(ram[12554]), .B2(n3260), 
        .ZN(n16795) );
  MOAI22 U25701 ( .A1(n28503), .A2(n3259), .B1(ram[12555]), .B2(n3260), 
        .ZN(n16796) );
  MOAI22 U25702 ( .A1(n28268), .A2(n3259), .B1(ram[12556]), .B2(n3260), 
        .ZN(n16797) );
  MOAI22 U25703 ( .A1(n28033), .A2(n3259), .B1(ram[12557]), .B2(n3260), 
        .ZN(n16798) );
  MOAI22 U25704 ( .A1(n27798), .A2(n3259), .B1(ram[12558]), .B2(n3260), 
        .ZN(n16799) );
  MOAI22 U25705 ( .A1(n27563), .A2(n3259), .B1(ram[12559]), .B2(n3260), 
        .ZN(n16800) );
  MOAI22 U25706 ( .A1(n29208), .A2(n3261), .B1(ram[12560]), .B2(n3262), 
        .ZN(n16801) );
  MOAI22 U25707 ( .A1(n28973), .A2(n3261), .B1(ram[12561]), .B2(n3262), 
        .ZN(n16802) );
  MOAI22 U25708 ( .A1(n28738), .A2(n3261), .B1(ram[12562]), .B2(n3262), 
        .ZN(n16803) );
  MOAI22 U25709 ( .A1(n28503), .A2(n3261), .B1(ram[12563]), .B2(n3262), 
        .ZN(n16804) );
  MOAI22 U25710 ( .A1(n28268), .A2(n3261), .B1(ram[12564]), .B2(n3262), 
        .ZN(n16805) );
  MOAI22 U25711 ( .A1(n28033), .A2(n3261), .B1(ram[12565]), .B2(n3262), 
        .ZN(n16806) );
  MOAI22 U25712 ( .A1(n27798), .A2(n3261), .B1(ram[12566]), .B2(n3262), 
        .ZN(n16807) );
  MOAI22 U25713 ( .A1(n27563), .A2(n3261), .B1(ram[12567]), .B2(n3262), 
        .ZN(n16808) );
  MOAI22 U25714 ( .A1(n29208), .A2(n3263), .B1(ram[12568]), .B2(n3264), 
        .ZN(n16809) );
  MOAI22 U25715 ( .A1(n28973), .A2(n3263), .B1(ram[12569]), .B2(n3264), 
        .ZN(n16810) );
  MOAI22 U25716 ( .A1(n28738), .A2(n3263), .B1(ram[12570]), .B2(n3264), 
        .ZN(n16811) );
  MOAI22 U25717 ( .A1(n28503), .A2(n3263), .B1(ram[12571]), .B2(n3264), 
        .ZN(n16812) );
  MOAI22 U25718 ( .A1(n28268), .A2(n3263), .B1(ram[12572]), .B2(n3264), 
        .ZN(n16813) );
  MOAI22 U25719 ( .A1(n28033), .A2(n3263), .B1(ram[12573]), .B2(n3264), 
        .ZN(n16814) );
  MOAI22 U25720 ( .A1(n27798), .A2(n3263), .B1(ram[12574]), .B2(n3264), 
        .ZN(n16815) );
  MOAI22 U25721 ( .A1(n27563), .A2(n3263), .B1(ram[12575]), .B2(n3264), 
        .ZN(n16816) );
  MOAI22 U25722 ( .A1(n29208), .A2(n3265), .B1(ram[12576]), .B2(n3266), 
        .ZN(n16817) );
  MOAI22 U25723 ( .A1(n28973), .A2(n3265), .B1(ram[12577]), .B2(n3266), 
        .ZN(n16818) );
  MOAI22 U25724 ( .A1(n28738), .A2(n3265), .B1(ram[12578]), .B2(n3266), 
        .ZN(n16819) );
  MOAI22 U25725 ( .A1(n28503), .A2(n3265), .B1(ram[12579]), .B2(n3266), 
        .ZN(n16820) );
  MOAI22 U25726 ( .A1(n28268), .A2(n3265), .B1(ram[12580]), .B2(n3266), 
        .ZN(n16821) );
  MOAI22 U25727 ( .A1(n28033), .A2(n3265), .B1(ram[12581]), .B2(n3266), 
        .ZN(n16822) );
  MOAI22 U25728 ( .A1(n27798), .A2(n3265), .B1(ram[12582]), .B2(n3266), 
        .ZN(n16823) );
  MOAI22 U25729 ( .A1(n27563), .A2(n3265), .B1(ram[12583]), .B2(n3266), 
        .ZN(n16824) );
  MOAI22 U25730 ( .A1(n29209), .A2(n3267), .B1(ram[12584]), .B2(n3268), 
        .ZN(n16825) );
  MOAI22 U25731 ( .A1(n28974), .A2(n3267), .B1(ram[12585]), .B2(n3268), 
        .ZN(n16826) );
  MOAI22 U25732 ( .A1(n28739), .A2(n3267), .B1(ram[12586]), .B2(n3268), 
        .ZN(n16827) );
  MOAI22 U25733 ( .A1(n28504), .A2(n3267), .B1(ram[12587]), .B2(n3268), 
        .ZN(n16828) );
  MOAI22 U25734 ( .A1(n28269), .A2(n3267), .B1(ram[12588]), .B2(n3268), 
        .ZN(n16829) );
  MOAI22 U25735 ( .A1(n28034), .A2(n3267), .B1(ram[12589]), .B2(n3268), 
        .ZN(n16830) );
  MOAI22 U25736 ( .A1(n27799), .A2(n3267), .B1(ram[12590]), .B2(n3268), 
        .ZN(n16831) );
  MOAI22 U25737 ( .A1(n27564), .A2(n3267), .B1(ram[12591]), .B2(n3268), 
        .ZN(n16832) );
  MOAI22 U25738 ( .A1(n29209), .A2(n3269), .B1(ram[12592]), .B2(n3270), 
        .ZN(n16833) );
  MOAI22 U25739 ( .A1(n28974), .A2(n3269), .B1(ram[12593]), .B2(n3270), 
        .ZN(n16834) );
  MOAI22 U25740 ( .A1(n28739), .A2(n3269), .B1(ram[12594]), .B2(n3270), 
        .ZN(n16835) );
  MOAI22 U25741 ( .A1(n28504), .A2(n3269), .B1(ram[12595]), .B2(n3270), 
        .ZN(n16836) );
  MOAI22 U25742 ( .A1(n28269), .A2(n3269), .B1(ram[12596]), .B2(n3270), 
        .ZN(n16837) );
  MOAI22 U25743 ( .A1(n28034), .A2(n3269), .B1(ram[12597]), .B2(n3270), 
        .ZN(n16838) );
  MOAI22 U25744 ( .A1(n27799), .A2(n3269), .B1(ram[12598]), .B2(n3270), 
        .ZN(n16839) );
  MOAI22 U25745 ( .A1(n27564), .A2(n3269), .B1(ram[12599]), .B2(n3270), 
        .ZN(n16840) );
  MOAI22 U25746 ( .A1(n29209), .A2(n3271), .B1(ram[12600]), .B2(n3272), 
        .ZN(n16841) );
  MOAI22 U25747 ( .A1(n28974), .A2(n3271), .B1(ram[12601]), .B2(n3272), 
        .ZN(n16842) );
  MOAI22 U25748 ( .A1(n28739), .A2(n3271), .B1(ram[12602]), .B2(n3272), 
        .ZN(n16843) );
  MOAI22 U25749 ( .A1(n28504), .A2(n3271), .B1(ram[12603]), .B2(n3272), 
        .ZN(n16844) );
  MOAI22 U25750 ( .A1(n28269), .A2(n3271), .B1(ram[12604]), .B2(n3272), 
        .ZN(n16845) );
  MOAI22 U25751 ( .A1(n28034), .A2(n3271), .B1(ram[12605]), .B2(n3272), 
        .ZN(n16846) );
  MOAI22 U25752 ( .A1(n27799), .A2(n3271), .B1(ram[12606]), .B2(n3272), 
        .ZN(n16847) );
  MOAI22 U25753 ( .A1(n27564), .A2(n3271), .B1(ram[12607]), .B2(n3272), 
        .ZN(n16848) );
  MOAI22 U25754 ( .A1(n29209), .A2(n3273), .B1(ram[12608]), .B2(n3274), 
        .ZN(n16849) );
  MOAI22 U25755 ( .A1(n28974), .A2(n3273), .B1(ram[12609]), .B2(n3274), 
        .ZN(n16850) );
  MOAI22 U25756 ( .A1(n28739), .A2(n3273), .B1(ram[12610]), .B2(n3274), 
        .ZN(n16851) );
  MOAI22 U25757 ( .A1(n28504), .A2(n3273), .B1(ram[12611]), .B2(n3274), 
        .ZN(n16852) );
  MOAI22 U25758 ( .A1(n28269), .A2(n3273), .B1(ram[12612]), .B2(n3274), 
        .ZN(n16853) );
  MOAI22 U25759 ( .A1(n28034), .A2(n3273), .B1(ram[12613]), .B2(n3274), 
        .ZN(n16854) );
  MOAI22 U25760 ( .A1(n27799), .A2(n3273), .B1(ram[12614]), .B2(n3274), 
        .ZN(n16855) );
  MOAI22 U25761 ( .A1(n27564), .A2(n3273), .B1(ram[12615]), .B2(n3274), 
        .ZN(n16856) );
  MOAI22 U25762 ( .A1(n29209), .A2(n3275), .B1(ram[12616]), .B2(n3276), 
        .ZN(n16857) );
  MOAI22 U25763 ( .A1(n28974), .A2(n3275), .B1(ram[12617]), .B2(n3276), 
        .ZN(n16858) );
  MOAI22 U25764 ( .A1(n28739), .A2(n3275), .B1(ram[12618]), .B2(n3276), 
        .ZN(n16859) );
  MOAI22 U25765 ( .A1(n28504), .A2(n3275), .B1(ram[12619]), .B2(n3276), 
        .ZN(n16860) );
  MOAI22 U25766 ( .A1(n28269), .A2(n3275), .B1(ram[12620]), .B2(n3276), 
        .ZN(n16861) );
  MOAI22 U25767 ( .A1(n28034), .A2(n3275), .B1(ram[12621]), .B2(n3276), 
        .ZN(n16862) );
  MOAI22 U25768 ( .A1(n27799), .A2(n3275), .B1(ram[12622]), .B2(n3276), 
        .ZN(n16863) );
  MOAI22 U25769 ( .A1(n27564), .A2(n3275), .B1(ram[12623]), .B2(n3276), 
        .ZN(n16864) );
  MOAI22 U25770 ( .A1(n29209), .A2(n3277), .B1(ram[12624]), .B2(n3278), 
        .ZN(n16865) );
  MOAI22 U25771 ( .A1(n28974), .A2(n3277), .B1(ram[12625]), .B2(n3278), 
        .ZN(n16866) );
  MOAI22 U25772 ( .A1(n28739), .A2(n3277), .B1(ram[12626]), .B2(n3278), 
        .ZN(n16867) );
  MOAI22 U25773 ( .A1(n28504), .A2(n3277), .B1(ram[12627]), .B2(n3278), 
        .ZN(n16868) );
  MOAI22 U25774 ( .A1(n28269), .A2(n3277), .B1(ram[12628]), .B2(n3278), 
        .ZN(n16869) );
  MOAI22 U25775 ( .A1(n28034), .A2(n3277), .B1(ram[12629]), .B2(n3278), 
        .ZN(n16870) );
  MOAI22 U25776 ( .A1(n27799), .A2(n3277), .B1(ram[12630]), .B2(n3278), 
        .ZN(n16871) );
  MOAI22 U25777 ( .A1(n27564), .A2(n3277), .B1(ram[12631]), .B2(n3278), 
        .ZN(n16872) );
  MOAI22 U25778 ( .A1(n29209), .A2(n3279), .B1(ram[12632]), .B2(n3280), 
        .ZN(n16873) );
  MOAI22 U25779 ( .A1(n28974), .A2(n3279), .B1(ram[12633]), .B2(n3280), 
        .ZN(n16874) );
  MOAI22 U25780 ( .A1(n28739), .A2(n3279), .B1(ram[12634]), .B2(n3280), 
        .ZN(n16875) );
  MOAI22 U25781 ( .A1(n28504), .A2(n3279), .B1(ram[12635]), .B2(n3280), 
        .ZN(n16876) );
  MOAI22 U25782 ( .A1(n28269), .A2(n3279), .B1(ram[12636]), .B2(n3280), 
        .ZN(n16877) );
  MOAI22 U25783 ( .A1(n28034), .A2(n3279), .B1(ram[12637]), .B2(n3280), 
        .ZN(n16878) );
  MOAI22 U25784 ( .A1(n27799), .A2(n3279), .B1(ram[12638]), .B2(n3280), 
        .ZN(n16879) );
  MOAI22 U25785 ( .A1(n27564), .A2(n3279), .B1(ram[12639]), .B2(n3280), 
        .ZN(n16880) );
  MOAI22 U25786 ( .A1(n29209), .A2(n3281), .B1(ram[12640]), .B2(n3282), 
        .ZN(n16881) );
  MOAI22 U25787 ( .A1(n28974), .A2(n3281), .B1(ram[12641]), .B2(n3282), 
        .ZN(n16882) );
  MOAI22 U25788 ( .A1(n28739), .A2(n3281), .B1(ram[12642]), .B2(n3282), 
        .ZN(n16883) );
  MOAI22 U25789 ( .A1(n28504), .A2(n3281), .B1(ram[12643]), .B2(n3282), 
        .ZN(n16884) );
  MOAI22 U25790 ( .A1(n28269), .A2(n3281), .B1(ram[12644]), .B2(n3282), 
        .ZN(n16885) );
  MOAI22 U25791 ( .A1(n28034), .A2(n3281), .B1(ram[12645]), .B2(n3282), 
        .ZN(n16886) );
  MOAI22 U25792 ( .A1(n27799), .A2(n3281), .B1(ram[12646]), .B2(n3282), 
        .ZN(n16887) );
  MOAI22 U25793 ( .A1(n27564), .A2(n3281), .B1(ram[12647]), .B2(n3282), 
        .ZN(n16888) );
  MOAI22 U25794 ( .A1(n29209), .A2(n3283), .B1(ram[12648]), .B2(n3284), 
        .ZN(n16889) );
  MOAI22 U25795 ( .A1(n28974), .A2(n3283), .B1(ram[12649]), .B2(n3284), 
        .ZN(n16890) );
  MOAI22 U25796 ( .A1(n28739), .A2(n3283), .B1(ram[12650]), .B2(n3284), 
        .ZN(n16891) );
  MOAI22 U25797 ( .A1(n28504), .A2(n3283), .B1(ram[12651]), .B2(n3284), 
        .ZN(n16892) );
  MOAI22 U25798 ( .A1(n28269), .A2(n3283), .B1(ram[12652]), .B2(n3284), 
        .ZN(n16893) );
  MOAI22 U25799 ( .A1(n28034), .A2(n3283), .B1(ram[12653]), .B2(n3284), 
        .ZN(n16894) );
  MOAI22 U25800 ( .A1(n27799), .A2(n3283), .B1(ram[12654]), .B2(n3284), 
        .ZN(n16895) );
  MOAI22 U25801 ( .A1(n27564), .A2(n3283), .B1(ram[12655]), .B2(n3284), 
        .ZN(n16896) );
  MOAI22 U25802 ( .A1(n29209), .A2(n3285), .B1(ram[12656]), .B2(n3286), 
        .ZN(n16897) );
  MOAI22 U25803 ( .A1(n28974), .A2(n3285), .B1(ram[12657]), .B2(n3286), 
        .ZN(n16898) );
  MOAI22 U25804 ( .A1(n28739), .A2(n3285), .B1(ram[12658]), .B2(n3286), 
        .ZN(n16899) );
  MOAI22 U25805 ( .A1(n28504), .A2(n3285), .B1(ram[12659]), .B2(n3286), 
        .ZN(n16900) );
  MOAI22 U25806 ( .A1(n28269), .A2(n3285), .B1(ram[12660]), .B2(n3286), 
        .ZN(n16901) );
  MOAI22 U25807 ( .A1(n28034), .A2(n3285), .B1(ram[12661]), .B2(n3286), 
        .ZN(n16902) );
  MOAI22 U25808 ( .A1(n27799), .A2(n3285), .B1(ram[12662]), .B2(n3286), 
        .ZN(n16903) );
  MOAI22 U25809 ( .A1(n27564), .A2(n3285), .B1(ram[12663]), .B2(n3286), 
        .ZN(n16904) );
  MOAI22 U25810 ( .A1(n29209), .A2(n3287), .B1(ram[12664]), .B2(n3288), 
        .ZN(n16905) );
  MOAI22 U25811 ( .A1(n28974), .A2(n3287), .B1(ram[12665]), .B2(n3288), 
        .ZN(n16906) );
  MOAI22 U25812 ( .A1(n28739), .A2(n3287), .B1(ram[12666]), .B2(n3288), 
        .ZN(n16907) );
  MOAI22 U25813 ( .A1(n28504), .A2(n3287), .B1(ram[12667]), .B2(n3288), 
        .ZN(n16908) );
  MOAI22 U25814 ( .A1(n28269), .A2(n3287), .B1(ram[12668]), .B2(n3288), 
        .ZN(n16909) );
  MOAI22 U25815 ( .A1(n28034), .A2(n3287), .B1(ram[12669]), .B2(n3288), 
        .ZN(n16910) );
  MOAI22 U25816 ( .A1(n27799), .A2(n3287), .B1(ram[12670]), .B2(n3288), 
        .ZN(n16911) );
  MOAI22 U25817 ( .A1(n27564), .A2(n3287), .B1(ram[12671]), .B2(n3288), 
        .ZN(n16912) );
  MOAI22 U25818 ( .A1(n29209), .A2(n3289), .B1(ram[12672]), .B2(n3290), 
        .ZN(n16913) );
  MOAI22 U25819 ( .A1(n28974), .A2(n3289), .B1(ram[12673]), .B2(n3290), 
        .ZN(n16914) );
  MOAI22 U25820 ( .A1(n28739), .A2(n3289), .B1(ram[12674]), .B2(n3290), 
        .ZN(n16915) );
  MOAI22 U25821 ( .A1(n28504), .A2(n3289), .B1(ram[12675]), .B2(n3290), 
        .ZN(n16916) );
  MOAI22 U25822 ( .A1(n28269), .A2(n3289), .B1(ram[12676]), .B2(n3290), 
        .ZN(n16917) );
  MOAI22 U25823 ( .A1(n28034), .A2(n3289), .B1(ram[12677]), .B2(n3290), 
        .ZN(n16918) );
  MOAI22 U25824 ( .A1(n27799), .A2(n3289), .B1(ram[12678]), .B2(n3290), 
        .ZN(n16919) );
  MOAI22 U25825 ( .A1(n27564), .A2(n3289), .B1(ram[12679]), .B2(n3290), 
        .ZN(n16920) );
  MOAI22 U25826 ( .A1(n29209), .A2(n3291), .B1(ram[12680]), .B2(n3292), 
        .ZN(n16921) );
  MOAI22 U25827 ( .A1(n28974), .A2(n3291), .B1(ram[12681]), .B2(n3292), 
        .ZN(n16922) );
  MOAI22 U25828 ( .A1(n28739), .A2(n3291), .B1(ram[12682]), .B2(n3292), 
        .ZN(n16923) );
  MOAI22 U25829 ( .A1(n28504), .A2(n3291), .B1(ram[12683]), .B2(n3292), 
        .ZN(n16924) );
  MOAI22 U25830 ( .A1(n28269), .A2(n3291), .B1(ram[12684]), .B2(n3292), 
        .ZN(n16925) );
  MOAI22 U25831 ( .A1(n28034), .A2(n3291), .B1(ram[12685]), .B2(n3292), 
        .ZN(n16926) );
  MOAI22 U25832 ( .A1(n27799), .A2(n3291), .B1(ram[12686]), .B2(n3292), 
        .ZN(n16927) );
  MOAI22 U25833 ( .A1(n27564), .A2(n3291), .B1(ram[12687]), .B2(n3292), 
        .ZN(n16928) );
  MOAI22 U25834 ( .A1(n29210), .A2(n3293), .B1(ram[12688]), .B2(n3294), 
        .ZN(n16929) );
  MOAI22 U25835 ( .A1(n28975), .A2(n3293), .B1(ram[12689]), .B2(n3294), 
        .ZN(n16930) );
  MOAI22 U25836 ( .A1(n28740), .A2(n3293), .B1(ram[12690]), .B2(n3294), 
        .ZN(n16931) );
  MOAI22 U25837 ( .A1(n28505), .A2(n3293), .B1(ram[12691]), .B2(n3294), 
        .ZN(n16932) );
  MOAI22 U25838 ( .A1(n28270), .A2(n3293), .B1(ram[12692]), .B2(n3294), 
        .ZN(n16933) );
  MOAI22 U25839 ( .A1(n28035), .A2(n3293), .B1(ram[12693]), .B2(n3294), 
        .ZN(n16934) );
  MOAI22 U25840 ( .A1(n27800), .A2(n3293), .B1(ram[12694]), .B2(n3294), 
        .ZN(n16935) );
  MOAI22 U25841 ( .A1(n27565), .A2(n3293), .B1(ram[12695]), .B2(n3294), 
        .ZN(n16936) );
  MOAI22 U25842 ( .A1(n29210), .A2(n3295), .B1(ram[12696]), .B2(n3296), 
        .ZN(n16937) );
  MOAI22 U25843 ( .A1(n28975), .A2(n3295), .B1(ram[12697]), .B2(n3296), 
        .ZN(n16938) );
  MOAI22 U25844 ( .A1(n28740), .A2(n3295), .B1(ram[12698]), .B2(n3296), 
        .ZN(n16939) );
  MOAI22 U25845 ( .A1(n28505), .A2(n3295), .B1(ram[12699]), .B2(n3296), 
        .ZN(n16940) );
  MOAI22 U25846 ( .A1(n28270), .A2(n3295), .B1(ram[12700]), .B2(n3296), 
        .ZN(n16941) );
  MOAI22 U25847 ( .A1(n28035), .A2(n3295), .B1(ram[12701]), .B2(n3296), 
        .ZN(n16942) );
  MOAI22 U25848 ( .A1(n27800), .A2(n3295), .B1(ram[12702]), .B2(n3296), 
        .ZN(n16943) );
  MOAI22 U25849 ( .A1(n27565), .A2(n3295), .B1(ram[12703]), .B2(n3296), 
        .ZN(n16944) );
  MOAI22 U25850 ( .A1(n29210), .A2(n3297), .B1(ram[12704]), .B2(n3298), 
        .ZN(n16945) );
  MOAI22 U25851 ( .A1(n28975), .A2(n3297), .B1(ram[12705]), .B2(n3298), 
        .ZN(n16946) );
  MOAI22 U25852 ( .A1(n28740), .A2(n3297), .B1(ram[12706]), .B2(n3298), 
        .ZN(n16947) );
  MOAI22 U25853 ( .A1(n28505), .A2(n3297), .B1(ram[12707]), .B2(n3298), 
        .ZN(n16948) );
  MOAI22 U25854 ( .A1(n28270), .A2(n3297), .B1(ram[12708]), .B2(n3298), 
        .ZN(n16949) );
  MOAI22 U25855 ( .A1(n28035), .A2(n3297), .B1(ram[12709]), .B2(n3298), 
        .ZN(n16950) );
  MOAI22 U25856 ( .A1(n27800), .A2(n3297), .B1(ram[12710]), .B2(n3298), 
        .ZN(n16951) );
  MOAI22 U25857 ( .A1(n27565), .A2(n3297), .B1(ram[12711]), .B2(n3298), 
        .ZN(n16952) );
  MOAI22 U25858 ( .A1(n29210), .A2(n3299), .B1(ram[12712]), .B2(n3300), 
        .ZN(n16953) );
  MOAI22 U25859 ( .A1(n28975), .A2(n3299), .B1(ram[12713]), .B2(n3300), 
        .ZN(n16954) );
  MOAI22 U25860 ( .A1(n28740), .A2(n3299), .B1(ram[12714]), .B2(n3300), 
        .ZN(n16955) );
  MOAI22 U25861 ( .A1(n28505), .A2(n3299), .B1(ram[12715]), .B2(n3300), 
        .ZN(n16956) );
  MOAI22 U25862 ( .A1(n28270), .A2(n3299), .B1(ram[12716]), .B2(n3300), 
        .ZN(n16957) );
  MOAI22 U25863 ( .A1(n28035), .A2(n3299), .B1(ram[12717]), .B2(n3300), 
        .ZN(n16958) );
  MOAI22 U25864 ( .A1(n27800), .A2(n3299), .B1(ram[12718]), .B2(n3300), 
        .ZN(n16959) );
  MOAI22 U25865 ( .A1(n27565), .A2(n3299), .B1(ram[12719]), .B2(n3300), 
        .ZN(n16960) );
  MOAI22 U25866 ( .A1(n29210), .A2(n3301), .B1(ram[12720]), .B2(n3302), 
        .ZN(n16961) );
  MOAI22 U25867 ( .A1(n28975), .A2(n3301), .B1(ram[12721]), .B2(n3302), 
        .ZN(n16962) );
  MOAI22 U25868 ( .A1(n28740), .A2(n3301), .B1(ram[12722]), .B2(n3302), 
        .ZN(n16963) );
  MOAI22 U25869 ( .A1(n28505), .A2(n3301), .B1(ram[12723]), .B2(n3302), 
        .ZN(n16964) );
  MOAI22 U25870 ( .A1(n28270), .A2(n3301), .B1(ram[12724]), .B2(n3302), 
        .ZN(n16965) );
  MOAI22 U25871 ( .A1(n28035), .A2(n3301), .B1(ram[12725]), .B2(n3302), 
        .ZN(n16966) );
  MOAI22 U25872 ( .A1(n27800), .A2(n3301), .B1(ram[12726]), .B2(n3302), 
        .ZN(n16967) );
  MOAI22 U25873 ( .A1(n27565), .A2(n3301), .B1(ram[12727]), .B2(n3302), 
        .ZN(n16968) );
  MOAI22 U25874 ( .A1(n29210), .A2(n3303), .B1(ram[12728]), .B2(n3304), 
        .ZN(n16969) );
  MOAI22 U25875 ( .A1(n28975), .A2(n3303), .B1(ram[12729]), .B2(n3304), 
        .ZN(n16970) );
  MOAI22 U25876 ( .A1(n28740), .A2(n3303), .B1(ram[12730]), .B2(n3304), 
        .ZN(n16971) );
  MOAI22 U25877 ( .A1(n28505), .A2(n3303), .B1(ram[12731]), .B2(n3304), 
        .ZN(n16972) );
  MOAI22 U25878 ( .A1(n28270), .A2(n3303), .B1(ram[12732]), .B2(n3304), 
        .ZN(n16973) );
  MOAI22 U25879 ( .A1(n28035), .A2(n3303), .B1(ram[12733]), .B2(n3304), 
        .ZN(n16974) );
  MOAI22 U25880 ( .A1(n27800), .A2(n3303), .B1(ram[12734]), .B2(n3304), 
        .ZN(n16975) );
  MOAI22 U25881 ( .A1(n27565), .A2(n3303), .B1(ram[12735]), .B2(n3304), 
        .ZN(n16976) );
  MOAI22 U25882 ( .A1(n29210), .A2(n3305), .B1(ram[12736]), .B2(n3306), 
        .ZN(n16977) );
  MOAI22 U25883 ( .A1(n28975), .A2(n3305), .B1(ram[12737]), .B2(n3306), 
        .ZN(n16978) );
  MOAI22 U25884 ( .A1(n28740), .A2(n3305), .B1(ram[12738]), .B2(n3306), 
        .ZN(n16979) );
  MOAI22 U25885 ( .A1(n28505), .A2(n3305), .B1(ram[12739]), .B2(n3306), 
        .ZN(n16980) );
  MOAI22 U25886 ( .A1(n28270), .A2(n3305), .B1(ram[12740]), .B2(n3306), 
        .ZN(n16981) );
  MOAI22 U25887 ( .A1(n28035), .A2(n3305), .B1(ram[12741]), .B2(n3306), 
        .ZN(n16982) );
  MOAI22 U25888 ( .A1(n27800), .A2(n3305), .B1(ram[12742]), .B2(n3306), 
        .ZN(n16983) );
  MOAI22 U25889 ( .A1(n27565), .A2(n3305), .B1(ram[12743]), .B2(n3306), 
        .ZN(n16984) );
  MOAI22 U25890 ( .A1(n29210), .A2(n3307), .B1(ram[12744]), .B2(n3308), 
        .ZN(n16985) );
  MOAI22 U25891 ( .A1(n28975), .A2(n3307), .B1(ram[12745]), .B2(n3308), 
        .ZN(n16986) );
  MOAI22 U25892 ( .A1(n28740), .A2(n3307), .B1(ram[12746]), .B2(n3308), 
        .ZN(n16987) );
  MOAI22 U25893 ( .A1(n28505), .A2(n3307), .B1(ram[12747]), .B2(n3308), 
        .ZN(n16988) );
  MOAI22 U25894 ( .A1(n28270), .A2(n3307), .B1(ram[12748]), .B2(n3308), 
        .ZN(n16989) );
  MOAI22 U25895 ( .A1(n28035), .A2(n3307), .B1(ram[12749]), .B2(n3308), 
        .ZN(n16990) );
  MOAI22 U25896 ( .A1(n27800), .A2(n3307), .B1(ram[12750]), .B2(n3308), 
        .ZN(n16991) );
  MOAI22 U25897 ( .A1(n27565), .A2(n3307), .B1(ram[12751]), .B2(n3308), 
        .ZN(n16992) );
  MOAI22 U25898 ( .A1(n29210), .A2(n3309), .B1(ram[12752]), .B2(n3310), 
        .ZN(n16993) );
  MOAI22 U25899 ( .A1(n28975), .A2(n3309), .B1(ram[12753]), .B2(n3310), 
        .ZN(n16994) );
  MOAI22 U25900 ( .A1(n28740), .A2(n3309), .B1(ram[12754]), .B2(n3310), 
        .ZN(n16995) );
  MOAI22 U25901 ( .A1(n28505), .A2(n3309), .B1(ram[12755]), .B2(n3310), 
        .ZN(n16996) );
  MOAI22 U25902 ( .A1(n28270), .A2(n3309), .B1(ram[12756]), .B2(n3310), 
        .ZN(n16997) );
  MOAI22 U25903 ( .A1(n28035), .A2(n3309), .B1(ram[12757]), .B2(n3310), 
        .ZN(n16998) );
  MOAI22 U25904 ( .A1(n27800), .A2(n3309), .B1(ram[12758]), .B2(n3310), 
        .ZN(n16999) );
  MOAI22 U25905 ( .A1(n27565), .A2(n3309), .B1(ram[12759]), .B2(n3310), 
        .ZN(n17000) );
  MOAI22 U25906 ( .A1(n29210), .A2(n3311), .B1(ram[12760]), .B2(n3312), 
        .ZN(n17001) );
  MOAI22 U25907 ( .A1(n28975), .A2(n3311), .B1(ram[12761]), .B2(n3312), 
        .ZN(n17002) );
  MOAI22 U25908 ( .A1(n28740), .A2(n3311), .B1(ram[12762]), .B2(n3312), 
        .ZN(n17003) );
  MOAI22 U25909 ( .A1(n28505), .A2(n3311), .B1(ram[12763]), .B2(n3312), 
        .ZN(n17004) );
  MOAI22 U25910 ( .A1(n28270), .A2(n3311), .B1(ram[12764]), .B2(n3312), 
        .ZN(n17005) );
  MOAI22 U25911 ( .A1(n28035), .A2(n3311), .B1(ram[12765]), .B2(n3312), 
        .ZN(n17006) );
  MOAI22 U25912 ( .A1(n27800), .A2(n3311), .B1(ram[12766]), .B2(n3312), 
        .ZN(n17007) );
  MOAI22 U25913 ( .A1(n27565), .A2(n3311), .B1(ram[12767]), .B2(n3312), 
        .ZN(n17008) );
  MOAI22 U25914 ( .A1(n29210), .A2(n3313), .B1(ram[12768]), .B2(n3314), 
        .ZN(n17009) );
  MOAI22 U25915 ( .A1(n28975), .A2(n3313), .B1(ram[12769]), .B2(n3314), 
        .ZN(n17010) );
  MOAI22 U25916 ( .A1(n28740), .A2(n3313), .B1(ram[12770]), .B2(n3314), 
        .ZN(n17011) );
  MOAI22 U25917 ( .A1(n28505), .A2(n3313), .B1(ram[12771]), .B2(n3314), 
        .ZN(n17012) );
  MOAI22 U25918 ( .A1(n28270), .A2(n3313), .B1(ram[12772]), .B2(n3314), 
        .ZN(n17013) );
  MOAI22 U25919 ( .A1(n28035), .A2(n3313), .B1(ram[12773]), .B2(n3314), 
        .ZN(n17014) );
  MOAI22 U25920 ( .A1(n27800), .A2(n3313), .B1(ram[12774]), .B2(n3314), 
        .ZN(n17015) );
  MOAI22 U25921 ( .A1(n27565), .A2(n3313), .B1(ram[12775]), .B2(n3314), 
        .ZN(n17016) );
  MOAI22 U25922 ( .A1(n29210), .A2(n3315), .B1(ram[12776]), .B2(n3316), 
        .ZN(n17017) );
  MOAI22 U25923 ( .A1(n28975), .A2(n3315), .B1(ram[12777]), .B2(n3316), 
        .ZN(n17018) );
  MOAI22 U25924 ( .A1(n28740), .A2(n3315), .B1(ram[12778]), .B2(n3316), 
        .ZN(n17019) );
  MOAI22 U25925 ( .A1(n28505), .A2(n3315), .B1(ram[12779]), .B2(n3316), 
        .ZN(n17020) );
  MOAI22 U25926 ( .A1(n28270), .A2(n3315), .B1(ram[12780]), .B2(n3316), 
        .ZN(n17021) );
  MOAI22 U25927 ( .A1(n28035), .A2(n3315), .B1(ram[12781]), .B2(n3316), 
        .ZN(n17022) );
  MOAI22 U25928 ( .A1(n27800), .A2(n3315), .B1(ram[12782]), .B2(n3316), 
        .ZN(n17023) );
  MOAI22 U25929 ( .A1(n27565), .A2(n3315), .B1(ram[12783]), .B2(n3316), 
        .ZN(n17024) );
  MOAI22 U25930 ( .A1(n29210), .A2(n3317), .B1(ram[12784]), .B2(n3318), 
        .ZN(n17025) );
  MOAI22 U25931 ( .A1(n28975), .A2(n3317), .B1(ram[12785]), .B2(n3318), 
        .ZN(n17026) );
  MOAI22 U25932 ( .A1(n28740), .A2(n3317), .B1(ram[12786]), .B2(n3318), 
        .ZN(n17027) );
  MOAI22 U25933 ( .A1(n28505), .A2(n3317), .B1(ram[12787]), .B2(n3318), 
        .ZN(n17028) );
  MOAI22 U25934 ( .A1(n28270), .A2(n3317), .B1(ram[12788]), .B2(n3318), 
        .ZN(n17029) );
  MOAI22 U25935 ( .A1(n28035), .A2(n3317), .B1(ram[12789]), .B2(n3318), 
        .ZN(n17030) );
  MOAI22 U25936 ( .A1(n27800), .A2(n3317), .B1(ram[12790]), .B2(n3318), 
        .ZN(n17031) );
  MOAI22 U25937 ( .A1(n27565), .A2(n3317), .B1(ram[12791]), .B2(n3318), 
        .ZN(n17032) );
  MOAI22 U25938 ( .A1(n29211), .A2(n3319), .B1(ram[12792]), .B2(n3320), 
        .ZN(n17033) );
  MOAI22 U25939 ( .A1(n28976), .A2(n3319), .B1(ram[12793]), .B2(n3320), 
        .ZN(n17034) );
  MOAI22 U25940 ( .A1(n28741), .A2(n3319), .B1(ram[12794]), .B2(n3320), 
        .ZN(n17035) );
  MOAI22 U25941 ( .A1(n28506), .A2(n3319), .B1(ram[12795]), .B2(n3320), 
        .ZN(n17036) );
  MOAI22 U25942 ( .A1(n28271), .A2(n3319), .B1(ram[12796]), .B2(n3320), 
        .ZN(n17037) );
  MOAI22 U25943 ( .A1(n28036), .A2(n3319), .B1(ram[12797]), .B2(n3320), 
        .ZN(n17038) );
  MOAI22 U25944 ( .A1(n27801), .A2(n3319), .B1(ram[12798]), .B2(n3320), 
        .ZN(n17039) );
  MOAI22 U25945 ( .A1(n27566), .A2(n3319), .B1(ram[12799]), .B2(n3320), 
        .ZN(n17040) );
  MOAI22 U25946 ( .A1(n29211), .A2(n3322), .B1(ram[12800]), .B2(n3323), 
        .ZN(n17041) );
  MOAI22 U25947 ( .A1(n28976), .A2(n3322), .B1(ram[12801]), .B2(n3323), 
        .ZN(n17042) );
  MOAI22 U25948 ( .A1(n28741), .A2(n3322), .B1(ram[12802]), .B2(n3323), 
        .ZN(n17043) );
  MOAI22 U25949 ( .A1(n28506), .A2(n3322), .B1(ram[12803]), .B2(n3323), 
        .ZN(n17044) );
  MOAI22 U25950 ( .A1(n28271), .A2(n3322), .B1(ram[12804]), .B2(n3323), 
        .ZN(n17045) );
  MOAI22 U25951 ( .A1(n28036), .A2(n3322), .B1(ram[12805]), .B2(n3323), 
        .ZN(n17046) );
  MOAI22 U25952 ( .A1(n27801), .A2(n3322), .B1(ram[12806]), .B2(n3323), 
        .ZN(n17047) );
  MOAI22 U25953 ( .A1(n27566), .A2(n3322), .B1(ram[12807]), .B2(n3323), 
        .ZN(n17048) );
  MOAI22 U25954 ( .A1(n29211), .A2(n3325), .B1(ram[12808]), .B2(n3326), 
        .ZN(n17049) );
  MOAI22 U25955 ( .A1(n28976), .A2(n3325), .B1(ram[12809]), .B2(n3326), 
        .ZN(n17050) );
  MOAI22 U25956 ( .A1(n28741), .A2(n3325), .B1(ram[12810]), .B2(n3326), 
        .ZN(n17051) );
  MOAI22 U25957 ( .A1(n28506), .A2(n3325), .B1(ram[12811]), .B2(n3326), 
        .ZN(n17052) );
  MOAI22 U25958 ( .A1(n28271), .A2(n3325), .B1(ram[12812]), .B2(n3326), 
        .ZN(n17053) );
  MOAI22 U25959 ( .A1(n28036), .A2(n3325), .B1(ram[12813]), .B2(n3326), 
        .ZN(n17054) );
  MOAI22 U25960 ( .A1(n27801), .A2(n3325), .B1(ram[12814]), .B2(n3326), 
        .ZN(n17055) );
  MOAI22 U25961 ( .A1(n27566), .A2(n3325), .B1(ram[12815]), .B2(n3326), 
        .ZN(n17056) );
  MOAI22 U25962 ( .A1(n29211), .A2(n3327), .B1(ram[12816]), .B2(n3328), 
        .ZN(n17057) );
  MOAI22 U25963 ( .A1(n28976), .A2(n3327), .B1(ram[12817]), .B2(n3328), 
        .ZN(n17058) );
  MOAI22 U25964 ( .A1(n28741), .A2(n3327), .B1(ram[12818]), .B2(n3328), 
        .ZN(n17059) );
  MOAI22 U25965 ( .A1(n28506), .A2(n3327), .B1(ram[12819]), .B2(n3328), 
        .ZN(n17060) );
  MOAI22 U25966 ( .A1(n28271), .A2(n3327), .B1(ram[12820]), .B2(n3328), 
        .ZN(n17061) );
  MOAI22 U25967 ( .A1(n28036), .A2(n3327), .B1(ram[12821]), .B2(n3328), 
        .ZN(n17062) );
  MOAI22 U25968 ( .A1(n27801), .A2(n3327), .B1(ram[12822]), .B2(n3328), 
        .ZN(n17063) );
  MOAI22 U25969 ( .A1(n27566), .A2(n3327), .B1(ram[12823]), .B2(n3328), 
        .ZN(n17064) );
  MOAI22 U25970 ( .A1(n29211), .A2(n3329), .B1(ram[12824]), .B2(n3330), 
        .ZN(n17065) );
  MOAI22 U25971 ( .A1(n28976), .A2(n3329), .B1(ram[12825]), .B2(n3330), 
        .ZN(n17066) );
  MOAI22 U25972 ( .A1(n28741), .A2(n3329), .B1(ram[12826]), .B2(n3330), 
        .ZN(n17067) );
  MOAI22 U25973 ( .A1(n28506), .A2(n3329), .B1(ram[12827]), .B2(n3330), 
        .ZN(n17068) );
  MOAI22 U25974 ( .A1(n28271), .A2(n3329), .B1(ram[12828]), .B2(n3330), 
        .ZN(n17069) );
  MOAI22 U25975 ( .A1(n28036), .A2(n3329), .B1(ram[12829]), .B2(n3330), 
        .ZN(n17070) );
  MOAI22 U25976 ( .A1(n27801), .A2(n3329), .B1(ram[12830]), .B2(n3330), 
        .ZN(n17071) );
  MOAI22 U25977 ( .A1(n27566), .A2(n3329), .B1(ram[12831]), .B2(n3330), 
        .ZN(n17072) );
  MOAI22 U25978 ( .A1(n29211), .A2(n3331), .B1(ram[12832]), .B2(n3332), 
        .ZN(n17073) );
  MOAI22 U25979 ( .A1(n28976), .A2(n3331), .B1(ram[12833]), .B2(n3332), 
        .ZN(n17074) );
  MOAI22 U25980 ( .A1(n28741), .A2(n3331), .B1(ram[12834]), .B2(n3332), 
        .ZN(n17075) );
  MOAI22 U25981 ( .A1(n28506), .A2(n3331), .B1(ram[12835]), .B2(n3332), 
        .ZN(n17076) );
  MOAI22 U25982 ( .A1(n28271), .A2(n3331), .B1(ram[12836]), .B2(n3332), 
        .ZN(n17077) );
  MOAI22 U25983 ( .A1(n28036), .A2(n3331), .B1(ram[12837]), .B2(n3332), 
        .ZN(n17078) );
  MOAI22 U25984 ( .A1(n27801), .A2(n3331), .B1(ram[12838]), .B2(n3332), 
        .ZN(n17079) );
  MOAI22 U25985 ( .A1(n27566), .A2(n3331), .B1(ram[12839]), .B2(n3332), 
        .ZN(n17080) );
  MOAI22 U25986 ( .A1(n29211), .A2(n3333), .B1(ram[12840]), .B2(n3334), 
        .ZN(n17081) );
  MOAI22 U25987 ( .A1(n28976), .A2(n3333), .B1(ram[12841]), .B2(n3334), 
        .ZN(n17082) );
  MOAI22 U25988 ( .A1(n28741), .A2(n3333), .B1(ram[12842]), .B2(n3334), 
        .ZN(n17083) );
  MOAI22 U25989 ( .A1(n28506), .A2(n3333), .B1(ram[12843]), .B2(n3334), 
        .ZN(n17084) );
  MOAI22 U25990 ( .A1(n28271), .A2(n3333), .B1(ram[12844]), .B2(n3334), 
        .ZN(n17085) );
  MOAI22 U25991 ( .A1(n28036), .A2(n3333), .B1(ram[12845]), .B2(n3334), 
        .ZN(n17086) );
  MOAI22 U25992 ( .A1(n27801), .A2(n3333), .B1(ram[12846]), .B2(n3334), 
        .ZN(n17087) );
  MOAI22 U25993 ( .A1(n27566), .A2(n3333), .B1(ram[12847]), .B2(n3334), 
        .ZN(n17088) );
  MOAI22 U25994 ( .A1(n29211), .A2(n3335), .B1(ram[12848]), .B2(n3336), 
        .ZN(n17089) );
  MOAI22 U25995 ( .A1(n28976), .A2(n3335), .B1(ram[12849]), .B2(n3336), 
        .ZN(n17090) );
  MOAI22 U25996 ( .A1(n28741), .A2(n3335), .B1(ram[12850]), .B2(n3336), 
        .ZN(n17091) );
  MOAI22 U25997 ( .A1(n28506), .A2(n3335), .B1(ram[12851]), .B2(n3336), 
        .ZN(n17092) );
  MOAI22 U25998 ( .A1(n28271), .A2(n3335), .B1(ram[12852]), .B2(n3336), 
        .ZN(n17093) );
  MOAI22 U25999 ( .A1(n28036), .A2(n3335), .B1(ram[12853]), .B2(n3336), 
        .ZN(n17094) );
  MOAI22 U26000 ( .A1(n27801), .A2(n3335), .B1(ram[12854]), .B2(n3336), 
        .ZN(n17095) );
  MOAI22 U26001 ( .A1(n27566), .A2(n3335), .B1(ram[12855]), .B2(n3336), 
        .ZN(n17096) );
  MOAI22 U26002 ( .A1(n29211), .A2(n3337), .B1(ram[12856]), .B2(n3338), 
        .ZN(n17097) );
  MOAI22 U26003 ( .A1(n28976), .A2(n3337), .B1(ram[12857]), .B2(n3338), 
        .ZN(n17098) );
  MOAI22 U26004 ( .A1(n28741), .A2(n3337), .B1(ram[12858]), .B2(n3338), 
        .ZN(n17099) );
  MOAI22 U26005 ( .A1(n28506), .A2(n3337), .B1(ram[12859]), .B2(n3338), 
        .ZN(n17100) );
  MOAI22 U26006 ( .A1(n28271), .A2(n3337), .B1(ram[12860]), .B2(n3338), 
        .ZN(n17101) );
  MOAI22 U26007 ( .A1(n28036), .A2(n3337), .B1(ram[12861]), .B2(n3338), 
        .ZN(n17102) );
  MOAI22 U26008 ( .A1(n27801), .A2(n3337), .B1(ram[12862]), .B2(n3338), 
        .ZN(n17103) );
  MOAI22 U26009 ( .A1(n27566), .A2(n3337), .B1(ram[12863]), .B2(n3338), 
        .ZN(n17104) );
  MOAI22 U26010 ( .A1(n29211), .A2(n3339), .B1(ram[12864]), .B2(n3340), 
        .ZN(n17105) );
  MOAI22 U26011 ( .A1(n28976), .A2(n3339), .B1(ram[12865]), .B2(n3340), 
        .ZN(n17106) );
  MOAI22 U26012 ( .A1(n28741), .A2(n3339), .B1(ram[12866]), .B2(n3340), 
        .ZN(n17107) );
  MOAI22 U26013 ( .A1(n28506), .A2(n3339), .B1(ram[12867]), .B2(n3340), 
        .ZN(n17108) );
  MOAI22 U26014 ( .A1(n28271), .A2(n3339), .B1(ram[12868]), .B2(n3340), 
        .ZN(n17109) );
  MOAI22 U26015 ( .A1(n28036), .A2(n3339), .B1(ram[12869]), .B2(n3340), 
        .ZN(n17110) );
  MOAI22 U26016 ( .A1(n27801), .A2(n3339), .B1(ram[12870]), .B2(n3340), 
        .ZN(n17111) );
  MOAI22 U26017 ( .A1(n27566), .A2(n3339), .B1(ram[12871]), .B2(n3340), 
        .ZN(n17112) );
  MOAI22 U26018 ( .A1(n29211), .A2(n3341), .B1(ram[12872]), .B2(n3342), 
        .ZN(n17113) );
  MOAI22 U26019 ( .A1(n28976), .A2(n3341), .B1(ram[12873]), .B2(n3342), 
        .ZN(n17114) );
  MOAI22 U26020 ( .A1(n28741), .A2(n3341), .B1(ram[12874]), .B2(n3342), 
        .ZN(n17115) );
  MOAI22 U26021 ( .A1(n28506), .A2(n3341), .B1(ram[12875]), .B2(n3342), 
        .ZN(n17116) );
  MOAI22 U26022 ( .A1(n28271), .A2(n3341), .B1(ram[12876]), .B2(n3342), 
        .ZN(n17117) );
  MOAI22 U26023 ( .A1(n28036), .A2(n3341), .B1(ram[12877]), .B2(n3342), 
        .ZN(n17118) );
  MOAI22 U26024 ( .A1(n27801), .A2(n3341), .B1(ram[12878]), .B2(n3342), 
        .ZN(n17119) );
  MOAI22 U26025 ( .A1(n27566), .A2(n3341), .B1(ram[12879]), .B2(n3342), 
        .ZN(n17120) );
  MOAI22 U26026 ( .A1(n29211), .A2(n3343), .B1(ram[12880]), .B2(n3344), 
        .ZN(n17121) );
  MOAI22 U26027 ( .A1(n28976), .A2(n3343), .B1(ram[12881]), .B2(n3344), 
        .ZN(n17122) );
  MOAI22 U26028 ( .A1(n28741), .A2(n3343), .B1(ram[12882]), .B2(n3344), 
        .ZN(n17123) );
  MOAI22 U26029 ( .A1(n28506), .A2(n3343), .B1(ram[12883]), .B2(n3344), 
        .ZN(n17124) );
  MOAI22 U26030 ( .A1(n28271), .A2(n3343), .B1(ram[12884]), .B2(n3344), 
        .ZN(n17125) );
  MOAI22 U26031 ( .A1(n28036), .A2(n3343), .B1(ram[12885]), .B2(n3344), 
        .ZN(n17126) );
  MOAI22 U26032 ( .A1(n27801), .A2(n3343), .B1(ram[12886]), .B2(n3344), 
        .ZN(n17127) );
  MOAI22 U26033 ( .A1(n27566), .A2(n3343), .B1(ram[12887]), .B2(n3344), 
        .ZN(n17128) );
  MOAI22 U26034 ( .A1(n29211), .A2(n3345), .B1(ram[12888]), .B2(n3346), 
        .ZN(n17129) );
  MOAI22 U26035 ( .A1(n28976), .A2(n3345), .B1(ram[12889]), .B2(n3346), 
        .ZN(n17130) );
  MOAI22 U26036 ( .A1(n28741), .A2(n3345), .B1(ram[12890]), .B2(n3346), 
        .ZN(n17131) );
  MOAI22 U26037 ( .A1(n28506), .A2(n3345), .B1(ram[12891]), .B2(n3346), 
        .ZN(n17132) );
  MOAI22 U26038 ( .A1(n28271), .A2(n3345), .B1(ram[12892]), .B2(n3346), 
        .ZN(n17133) );
  MOAI22 U26039 ( .A1(n28036), .A2(n3345), .B1(ram[12893]), .B2(n3346), 
        .ZN(n17134) );
  MOAI22 U26040 ( .A1(n27801), .A2(n3345), .B1(ram[12894]), .B2(n3346), 
        .ZN(n17135) );
  MOAI22 U26041 ( .A1(n27566), .A2(n3345), .B1(ram[12895]), .B2(n3346), 
        .ZN(n17136) );
  MOAI22 U26042 ( .A1(n29212), .A2(n3347), .B1(ram[12896]), .B2(n3348), 
        .ZN(n17137) );
  MOAI22 U26043 ( .A1(n28977), .A2(n3347), .B1(ram[12897]), .B2(n3348), 
        .ZN(n17138) );
  MOAI22 U26044 ( .A1(n28742), .A2(n3347), .B1(ram[12898]), .B2(n3348), 
        .ZN(n17139) );
  MOAI22 U26045 ( .A1(n28507), .A2(n3347), .B1(ram[12899]), .B2(n3348), 
        .ZN(n17140) );
  MOAI22 U26046 ( .A1(n28272), .A2(n3347), .B1(ram[12900]), .B2(n3348), 
        .ZN(n17141) );
  MOAI22 U26047 ( .A1(n28037), .A2(n3347), .B1(ram[12901]), .B2(n3348), 
        .ZN(n17142) );
  MOAI22 U26048 ( .A1(n27802), .A2(n3347), .B1(ram[12902]), .B2(n3348), 
        .ZN(n17143) );
  MOAI22 U26049 ( .A1(n27567), .A2(n3347), .B1(ram[12903]), .B2(n3348), 
        .ZN(n17144) );
  MOAI22 U26050 ( .A1(n29212), .A2(n3349), .B1(ram[12904]), .B2(n3350), 
        .ZN(n17145) );
  MOAI22 U26051 ( .A1(n28977), .A2(n3349), .B1(ram[12905]), .B2(n3350), 
        .ZN(n17146) );
  MOAI22 U26052 ( .A1(n28742), .A2(n3349), .B1(ram[12906]), .B2(n3350), 
        .ZN(n17147) );
  MOAI22 U26053 ( .A1(n28507), .A2(n3349), .B1(ram[12907]), .B2(n3350), 
        .ZN(n17148) );
  MOAI22 U26054 ( .A1(n28272), .A2(n3349), .B1(ram[12908]), .B2(n3350), 
        .ZN(n17149) );
  MOAI22 U26055 ( .A1(n28037), .A2(n3349), .B1(ram[12909]), .B2(n3350), 
        .ZN(n17150) );
  MOAI22 U26056 ( .A1(n27802), .A2(n3349), .B1(ram[12910]), .B2(n3350), 
        .ZN(n17151) );
  MOAI22 U26057 ( .A1(n27567), .A2(n3349), .B1(ram[12911]), .B2(n3350), 
        .ZN(n17152) );
  MOAI22 U26058 ( .A1(n29212), .A2(n3351), .B1(ram[12912]), .B2(n3352), 
        .ZN(n17153) );
  MOAI22 U26059 ( .A1(n28977), .A2(n3351), .B1(ram[12913]), .B2(n3352), 
        .ZN(n17154) );
  MOAI22 U26060 ( .A1(n28742), .A2(n3351), .B1(ram[12914]), .B2(n3352), 
        .ZN(n17155) );
  MOAI22 U26061 ( .A1(n28507), .A2(n3351), .B1(ram[12915]), .B2(n3352), 
        .ZN(n17156) );
  MOAI22 U26062 ( .A1(n28272), .A2(n3351), .B1(ram[12916]), .B2(n3352), 
        .ZN(n17157) );
  MOAI22 U26063 ( .A1(n28037), .A2(n3351), .B1(ram[12917]), .B2(n3352), 
        .ZN(n17158) );
  MOAI22 U26064 ( .A1(n27802), .A2(n3351), .B1(ram[12918]), .B2(n3352), 
        .ZN(n17159) );
  MOAI22 U26065 ( .A1(n27567), .A2(n3351), .B1(ram[12919]), .B2(n3352), 
        .ZN(n17160) );
  MOAI22 U26066 ( .A1(n29212), .A2(n3353), .B1(ram[12920]), .B2(n3354), 
        .ZN(n17161) );
  MOAI22 U26067 ( .A1(n28977), .A2(n3353), .B1(ram[12921]), .B2(n3354), 
        .ZN(n17162) );
  MOAI22 U26068 ( .A1(n28742), .A2(n3353), .B1(ram[12922]), .B2(n3354), 
        .ZN(n17163) );
  MOAI22 U26069 ( .A1(n28507), .A2(n3353), .B1(ram[12923]), .B2(n3354), 
        .ZN(n17164) );
  MOAI22 U26070 ( .A1(n28272), .A2(n3353), .B1(ram[12924]), .B2(n3354), 
        .ZN(n17165) );
  MOAI22 U26071 ( .A1(n28037), .A2(n3353), .B1(ram[12925]), .B2(n3354), 
        .ZN(n17166) );
  MOAI22 U26072 ( .A1(n27802), .A2(n3353), .B1(ram[12926]), .B2(n3354), 
        .ZN(n17167) );
  MOAI22 U26073 ( .A1(n27567), .A2(n3353), .B1(ram[12927]), .B2(n3354), 
        .ZN(n17168) );
  MOAI22 U26074 ( .A1(n29212), .A2(n3355), .B1(ram[12928]), .B2(n3356), 
        .ZN(n17169) );
  MOAI22 U26075 ( .A1(n28977), .A2(n3355), .B1(ram[12929]), .B2(n3356), 
        .ZN(n17170) );
  MOAI22 U26076 ( .A1(n28742), .A2(n3355), .B1(ram[12930]), .B2(n3356), 
        .ZN(n17171) );
  MOAI22 U26077 ( .A1(n28507), .A2(n3355), .B1(ram[12931]), .B2(n3356), 
        .ZN(n17172) );
  MOAI22 U26078 ( .A1(n28272), .A2(n3355), .B1(ram[12932]), .B2(n3356), 
        .ZN(n17173) );
  MOAI22 U26079 ( .A1(n28037), .A2(n3355), .B1(ram[12933]), .B2(n3356), 
        .ZN(n17174) );
  MOAI22 U26080 ( .A1(n27802), .A2(n3355), .B1(ram[12934]), .B2(n3356), 
        .ZN(n17175) );
  MOAI22 U26081 ( .A1(n27567), .A2(n3355), .B1(ram[12935]), .B2(n3356), 
        .ZN(n17176) );
  MOAI22 U26082 ( .A1(n29212), .A2(n3357), .B1(ram[12936]), .B2(n3358), 
        .ZN(n17177) );
  MOAI22 U26083 ( .A1(n28977), .A2(n3357), .B1(ram[12937]), .B2(n3358), 
        .ZN(n17178) );
  MOAI22 U26084 ( .A1(n28742), .A2(n3357), .B1(ram[12938]), .B2(n3358), 
        .ZN(n17179) );
  MOAI22 U26085 ( .A1(n28507), .A2(n3357), .B1(ram[12939]), .B2(n3358), 
        .ZN(n17180) );
  MOAI22 U26086 ( .A1(n28272), .A2(n3357), .B1(ram[12940]), .B2(n3358), 
        .ZN(n17181) );
  MOAI22 U26087 ( .A1(n28037), .A2(n3357), .B1(ram[12941]), .B2(n3358), 
        .ZN(n17182) );
  MOAI22 U26088 ( .A1(n27802), .A2(n3357), .B1(ram[12942]), .B2(n3358), 
        .ZN(n17183) );
  MOAI22 U26089 ( .A1(n27567), .A2(n3357), .B1(ram[12943]), .B2(n3358), 
        .ZN(n17184) );
  MOAI22 U26090 ( .A1(n29212), .A2(n3359), .B1(ram[12944]), .B2(n3360), 
        .ZN(n17185) );
  MOAI22 U26091 ( .A1(n28977), .A2(n3359), .B1(ram[12945]), .B2(n3360), 
        .ZN(n17186) );
  MOAI22 U26092 ( .A1(n28742), .A2(n3359), .B1(ram[12946]), .B2(n3360), 
        .ZN(n17187) );
  MOAI22 U26093 ( .A1(n28507), .A2(n3359), .B1(ram[12947]), .B2(n3360), 
        .ZN(n17188) );
  MOAI22 U26094 ( .A1(n28272), .A2(n3359), .B1(ram[12948]), .B2(n3360), 
        .ZN(n17189) );
  MOAI22 U26095 ( .A1(n28037), .A2(n3359), .B1(ram[12949]), .B2(n3360), 
        .ZN(n17190) );
  MOAI22 U26096 ( .A1(n27802), .A2(n3359), .B1(ram[12950]), .B2(n3360), 
        .ZN(n17191) );
  MOAI22 U26097 ( .A1(n27567), .A2(n3359), .B1(ram[12951]), .B2(n3360), 
        .ZN(n17192) );
  MOAI22 U26098 ( .A1(n29212), .A2(n3361), .B1(ram[12952]), .B2(n3362), 
        .ZN(n17193) );
  MOAI22 U26099 ( .A1(n28977), .A2(n3361), .B1(ram[12953]), .B2(n3362), 
        .ZN(n17194) );
  MOAI22 U26100 ( .A1(n28742), .A2(n3361), .B1(ram[12954]), .B2(n3362), 
        .ZN(n17195) );
  MOAI22 U26101 ( .A1(n28507), .A2(n3361), .B1(ram[12955]), .B2(n3362), 
        .ZN(n17196) );
  MOAI22 U26102 ( .A1(n28272), .A2(n3361), .B1(ram[12956]), .B2(n3362), 
        .ZN(n17197) );
  MOAI22 U26103 ( .A1(n28037), .A2(n3361), .B1(ram[12957]), .B2(n3362), 
        .ZN(n17198) );
  MOAI22 U26104 ( .A1(n27802), .A2(n3361), .B1(ram[12958]), .B2(n3362), 
        .ZN(n17199) );
  MOAI22 U26105 ( .A1(n27567), .A2(n3361), .B1(ram[12959]), .B2(n3362), 
        .ZN(n17200) );
  MOAI22 U26106 ( .A1(n29212), .A2(n3363), .B1(ram[12960]), .B2(n3364), 
        .ZN(n17201) );
  MOAI22 U26107 ( .A1(n28977), .A2(n3363), .B1(ram[12961]), .B2(n3364), 
        .ZN(n17202) );
  MOAI22 U26108 ( .A1(n28742), .A2(n3363), .B1(ram[12962]), .B2(n3364), 
        .ZN(n17203) );
  MOAI22 U26109 ( .A1(n28507), .A2(n3363), .B1(ram[12963]), .B2(n3364), 
        .ZN(n17204) );
  MOAI22 U26110 ( .A1(n28272), .A2(n3363), .B1(ram[12964]), .B2(n3364), 
        .ZN(n17205) );
  MOAI22 U26111 ( .A1(n28037), .A2(n3363), .B1(ram[12965]), .B2(n3364), 
        .ZN(n17206) );
  MOAI22 U26112 ( .A1(n27802), .A2(n3363), .B1(ram[12966]), .B2(n3364), 
        .ZN(n17207) );
  MOAI22 U26113 ( .A1(n27567), .A2(n3363), .B1(ram[12967]), .B2(n3364), 
        .ZN(n17208) );
  MOAI22 U26114 ( .A1(n29212), .A2(n3365), .B1(ram[12968]), .B2(n3366), 
        .ZN(n17209) );
  MOAI22 U26115 ( .A1(n28977), .A2(n3365), .B1(ram[12969]), .B2(n3366), 
        .ZN(n17210) );
  MOAI22 U26116 ( .A1(n28742), .A2(n3365), .B1(ram[12970]), .B2(n3366), 
        .ZN(n17211) );
  MOAI22 U26117 ( .A1(n28507), .A2(n3365), .B1(ram[12971]), .B2(n3366), 
        .ZN(n17212) );
  MOAI22 U26118 ( .A1(n28272), .A2(n3365), .B1(ram[12972]), .B2(n3366), 
        .ZN(n17213) );
  MOAI22 U26119 ( .A1(n28037), .A2(n3365), .B1(ram[12973]), .B2(n3366), 
        .ZN(n17214) );
  MOAI22 U26120 ( .A1(n27802), .A2(n3365), .B1(ram[12974]), .B2(n3366), 
        .ZN(n17215) );
  MOAI22 U26121 ( .A1(n27567), .A2(n3365), .B1(ram[12975]), .B2(n3366), 
        .ZN(n17216) );
  MOAI22 U26122 ( .A1(n29212), .A2(n3367), .B1(ram[12976]), .B2(n3368), 
        .ZN(n17217) );
  MOAI22 U26123 ( .A1(n28977), .A2(n3367), .B1(ram[12977]), .B2(n3368), 
        .ZN(n17218) );
  MOAI22 U26124 ( .A1(n28742), .A2(n3367), .B1(ram[12978]), .B2(n3368), 
        .ZN(n17219) );
  MOAI22 U26125 ( .A1(n28507), .A2(n3367), .B1(ram[12979]), .B2(n3368), 
        .ZN(n17220) );
  MOAI22 U26126 ( .A1(n28272), .A2(n3367), .B1(ram[12980]), .B2(n3368), 
        .ZN(n17221) );
  MOAI22 U26127 ( .A1(n28037), .A2(n3367), .B1(ram[12981]), .B2(n3368), 
        .ZN(n17222) );
  MOAI22 U26128 ( .A1(n27802), .A2(n3367), .B1(ram[12982]), .B2(n3368), 
        .ZN(n17223) );
  MOAI22 U26129 ( .A1(n27567), .A2(n3367), .B1(ram[12983]), .B2(n3368), 
        .ZN(n17224) );
  MOAI22 U26130 ( .A1(n29212), .A2(n3369), .B1(ram[12984]), .B2(n3370), 
        .ZN(n17225) );
  MOAI22 U26131 ( .A1(n28977), .A2(n3369), .B1(ram[12985]), .B2(n3370), 
        .ZN(n17226) );
  MOAI22 U26132 ( .A1(n28742), .A2(n3369), .B1(ram[12986]), .B2(n3370), 
        .ZN(n17227) );
  MOAI22 U26133 ( .A1(n28507), .A2(n3369), .B1(ram[12987]), .B2(n3370), 
        .ZN(n17228) );
  MOAI22 U26134 ( .A1(n28272), .A2(n3369), .B1(ram[12988]), .B2(n3370), 
        .ZN(n17229) );
  MOAI22 U26135 ( .A1(n28037), .A2(n3369), .B1(ram[12989]), .B2(n3370), 
        .ZN(n17230) );
  MOAI22 U26136 ( .A1(n27802), .A2(n3369), .B1(ram[12990]), .B2(n3370), 
        .ZN(n17231) );
  MOAI22 U26137 ( .A1(n27567), .A2(n3369), .B1(ram[12991]), .B2(n3370), 
        .ZN(n17232) );
  MOAI22 U26138 ( .A1(n29212), .A2(n3371), .B1(ram[12992]), .B2(n3372), 
        .ZN(n17233) );
  MOAI22 U26139 ( .A1(n28977), .A2(n3371), .B1(ram[12993]), .B2(n3372), 
        .ZN(n17234) );
  MOAI22 U26140 ( .A1(n28742), .A2(n3371), .B1(ram[12994]), .B2(n3372), 
        .ZN(n17235) );
  MOAI22 U26141 ( .A1(n28507), .A2(n3371), .B1(ram[12995]), .B2(n3372), 
        .ZN(n17236) );
  MOAI22 U26142 ( .A1(n28272), .A2(n3371), .B1(ram[12996]), .B2(n3372), 
        .ZN(n17237) );
  MOAI22 U26143 ( .A1(n28037), .A2(n3371), .B1(ram[12997]), .B2(n3372), 
        .ZN(n17238) );
  MOAI22 U26144 ( .A1(n27802), .A2(n3371), .B1(ram[12998]), .B2(n3372), 
        .ZN(n17239) );
  MOAI22 U26145 ( .A1(n27567), .A2(n3371), .B1(ram[12999]), .B2(n3372), 
        .ZN(n17240) );
  MOAI22 U26146 ( .A1(n29213), .A2(n3373), .B1(ram[13000]), .B2(n3374), 
        .ZN(n17241) );
  MOAI22 U26147 ( .A1(n28978), .A2(n3373), .B1(ram[13001]), .B2(n3374), 
        .ZN(n17242) );
  MOAI22 U26148 ( .A1(n28743), .A2(n3373), .B1(ram[13002]), .B2(n3374), 
        .ZN(n17243) );
  MOAI22 U26149 ( .A1(n28508), .A2(n3373), .B1(ram[13003]), .B2(n3374), 
        .ZN(n17244) );
  MOAI22 U26150 ( .A1(n28273), .A2(n3373), .B1(ram[13004]), .B2(n3374), 
        .ZN(n17245) );
  MOAI22 U26151 ( .A1(n28038), .A2(n3373), .B1(ram[13005]), .B2(n3374), 
        .ZN(n17246) );
  MOAI22 U26152 ( .A1(n27803), .A2(n3373), .B1(ram[13006]), .B2(n3374), 
        .ZN(n17247) );
  MOAI22 U26153 ( .A1(n27568), .A2(n3373), .B1(ram[13007]), .B2(n3374), 
        .ZN(n17248) );
  MOAI22 U26154 ( .A1(n29213), .A2(n3375), .B1(ram[13008]), .B2(n3376), 
        .ZN(n17249) );
  MOAI22 U26155 ( .A1(n28978), .A2(n3375), .B1(ram[13009]), .B2(n3376), 
        .ZN(n17250) );
  MOAI22 U26156 ( .A1(n28743), .A2(n3375), .B1(ram[13010]), .B2(n3376), 
        .ZN(n17251) );
  MOAI22 U26157 ( .A1(n28508), .A2(n3375), .B1(ram[13011]), .B2(n3376), 
        .ZN(n17252) );
  MOAI22 U26158 ( .A1(n28273), .A2(n3375), .B1(ram[13012]), .B2(n3376), 
        .ZN(n17253) );
  MOAI22 U26159 ( .A1(n28038), .A2(n3375), .B1(ram[13013]), .B2(n3376), 
        .ZN(n17254) );
  MOAI22 U26160 ( .A1(n27803), .A2(n3375), .B1(ram[13014]), .B2(n3376), 
        .ZN(n17255) );
  MOAI22 U26161 ( .A1(n27568), .A2(n3375), .B1(ram[13015]), .B2(n3376), 
        .ZN(n17256) );
  MOAI22 U26162 ( .A1(n29213), .A2(n3377), .B1(ram[13016]), .B2(n3378), 
        .ZN(n17257) );
  MOAI22 U26163 ( .A1(n28978), .A2(n3377), .B1(ram[13017]), .B2(n3378), 
        .ZN(n17258) );
  MOAI22 U26164 ( .A1(n28743), .A2(n3377), .B1(ram[13018]), .B2(n3378), 
        .ZN(n17259) );
  MOAI22 U26165 ( .A1(n28508), .A2(n3377), .B1(ram[13019]), .B2(n3378), 
        .ZN(n17260) );
  MOAI22 U26166 ( .A1(n28273), .A2(n3377), .B1(ram[13020]), .B2(n3378), 
        .ZN(n17261) );
  MOAI22 U26167 ( .A1(n28038), .A2(n3377), .B1(ram[13021]), .B2(n3378), 
        .ZN(n17262) );
  MOAI22 U26168 ( .A1(n27803), .A2(n3377), .B1(ram[13022]), .B2(n3378), 
        .ZN(n17263) );
  MOAI22 U26169 ( .A1(n27568), .A2(n3377), .B1(ram[13023]), .B2(n3378), 
        .ZN(n17264) );
  MOAI22 U26170 ( .A1(n29213), .A2(n3379), .B1(ram[13024]), .B2(n3380), 
        .ZN(n17265) );
  MOAI22 U26171 ( .A1(n28978), .A2(n3379), .B1(ram[13025]), .B2(n3380), 
        .ZN(n17266) );
  MOAI22 U26172 ( .A1(n28743), .A2(n3379), .B1(ram[13026]), .B2(n3380), 
        .ZN(n17267) );
  MOAI22 U26173 ( .A1(n28508), .A2(n3379), .B1(ram[13027]), .B2(n3380), 
        .ZN(n17268) );
  MOAI22 U26174 ( .A1(n28273), .A2(n3379), .B1(ram[13028]), .B2(n3380), 
        .ZN(n17269) );
  MOAI22 U26175 ( .A1(n28038), .A2(n3379), .B1(ram[13029]), .B2(n3380), 
        .ZN(n17270) );
  MOAI22 U26176 ( .A1(n27803), .A2(n3379), .B1(ram[13030]), .B2(n3380), 
        .ZN(n17271) );
  MOAI22 U26177 ( .A1(n27568), .A2(n3379), .B1(ram[13031]), .B2(n3380), 
        .ZN(n17272) );
  MOAI22 U26178 ( .A1(n29213), .A2(n3381), .B1(ram[13032]), .B2(n3382), 
        .ZN(n17273) );
  MOAI22 U26179 ( .A1(n28978), .A2(n3381), .B1(ram[13033]), .B2(n3382), 
        .ZN(n17274) );
  MOAI22 U26180 ( .A1(n28743), .A2(n3381), .B1(ram[13034]), .B2(n3382), 
        .ZN(n17275) );
  MOAI22 U26181 ( .A1(n28508), .A2(n3381), .B1(ram[13035]), .B2(n3382), 
        .ZN(n17276) );
  MOAI22 U26182 ( .A1(n28273), .A2(n3381), .B1(ram[13036]), .B2(n3382), 
        .ZN(n17277) );
  MOAI22 U26183 ( .A1(n28038), .A2(n3381), .B1(ram[13037]), .B2(n3382), 
        .ZN(n17278) );
  MOAI22 U26184 ( .A1(n27803), .A2(n3381), .B1(ram[13038]), .B2(n3382), 
        .ZN(n17279) );
  MOAI22 U26185 ( .A1(n27568), .A2(n3381), .B1(ram[13039]), .B2(n3382), 
        .ZN(n17280) );
  MOAI22 U26186 ( .A1(n29213), .A2(n3383), .B1(ram[13040]), .B2(n3384), 
        .ZN(n17281) );
  MOAI22 U26187 ( .A1(n28978), .A2(n3383), .B1(ram[13041]), .B2(n3384), 
        .ZN(n17282) );
  MOAI22 U26188 ( .A1(n28743), .A2(n3383), .B1(ram[13042]), .B2(n3384), 
        .ZN(n17283) );
  MOAI22 U26189 ( .A1(n28508), .A2(n3383), .B1(ram[13043]), .B2(n3384), 
        .ZN(n17284) );
  MOAI22 U26190 ( .A1(n28273), .A2(n3383), .B1(ram[13044]), .B2(n3384), 
        .ZN(n17285) );
  MOAI22 U26191 ( .A1(n28038), .A2(n3383), .B1(ram[13045]), .B2(n3384), 
        .ZN(n17286) );
  MOAI22 U26192 ( .A1(n27803), .A2(n3383), .B1(ram[13046]), .B2(n3384), 
        .ZN(n17287) );
  MOAI22 U26193 ( .A1(n27568), .A2(n3383), .B1(ram[13047]), .B2(n3384), 
        .ZN(n17288) );
  MOAI22 U26194 ( .A1(n29213), .A2(n3385), .B1(ram[13048]), .B2(n3386), 
        .ZN(n17289) );
  MOAI22 U26195 ( .A1(n28978), .A2(n3385), .B1(ram[13049]), .B2(n3386), 
        .ZN(n17290) );
  MOAI22 U26196 ( .A1(n28743), .A2(n3385), .B1(ram[13050]), .B2(n3386), 
        .ZN(n17291) );
  MOAI22 U26197 ( .A1(n28508), .A2(n3385), .B1(ram[13051]), .B2(n3386), 
        .ZN(n17292) );
  MOAI22 U26198 ( .A1(n28273), .A2(n3385), .B1(ram[13052]), .B2(n3386), 
        .ZN(n17293) );
  MOAI22 U26199 ( .A1(n28038), .A2(n3385), .B1(ram[13053]), .B2(n3386), 
        .ZN(n17294) );
  MOAI22 U26200 ( .A1(n27803), .A2(n3385), .B1(ram[13054]), .B2(n3386), 
        .ZN(n17295) );
  MOAI22 U26201 ( .A1(n27568), .A2(n3385), .B1(ram[13055]), .B2(n3386), 
        .ZN(n17296) );
  MOAI22 U26202 ( .A1(n29213), .A2(n3387), .B1(ram[13056]), .B2(n3388), 
        .ZN(n17297) );
  MOAI22 U26203 ( .A1(n28978), .A2(n3387), .B1(ram[13057]), .B2(n3388), 
        .ZN(n17298) );
  MOAI22 U26204 ( .A1(n28743), .A2(n3387), .B1(ram[13058]), .B2(n3388), 
        .ZN(n17299) );
  MOAI22 U26205 ( .A1(n28508), .A2(n3387), .B1(ram[13059]), .B2(n3388), 
        .ZN(n17300) );
  MOAI22 U26206 ( .A1(n28273), .A2(n3387), .B1(ram[13060]), .B2(n3388), 
        .ZN(n17301) );
  MOAI22 U26207 ( .A1(n28038), .A2(n3387), .B1(ram[13061]), .B2(n3388), 
        .ZN(n17302) );
  MOAI22 U26208 ( .A1(n27803), .A2(n3387), .B1(ram[13062]), .B2(n3388), 
        .ZN(n17303) );
  MOAI22 U26209 ( .A1(n27568), .A2(n3387), .B1(ram[13063]), .B2(n3388), 
        .ZN(n17304) );
  MOAI22 U26210 ( .A1(n29213), .A2(n3389), .B1(ram[13064]), .B2(n3390), 
        .ZN(n17305) );
  MOAI22 U26211 ( .A1(n28978), .A2(n3389), .B1(ram[13065]), .B2(n3390), 
        .ZN(n17306) );
  MOAI22 U26212 ( .A1(n28743), .A2(n3389), .B1(ram[13066]), .B2(n3390), 
        .ZN(n17307) );
  MOAI22 U26213 ( .A1(n28508), .A2(n3389), .B1(ram[13067]), .B2(n3390), 
        .ZN(n17308) );
  MOAI22 U26214 ( .A1(n28273), .A2(n3389), .B1(ram[13068]), .B2(n3390), 
        .ZN(n17309) );
  MOAI22 U26215 ( .A1(n28038), .A2(n3389), .B1(ram[13069]), .B2(n3390), 
        .ZN(n17310) );
  MOAI22 U26216 ( .A1(n27803), .A2(n3389), .B1(ram[13070]), .B2(n3390), 
        .ZN(n17311) );
  MOAI22 U26217 ( .A1(n27568), .A2(n3389), .B1(ram[13071]), .B2(n3390), 
        .ZN(n17312) );
  MOAI22 U26218 ( .A1(n29213), .A2(n3391), .B1(ram[13072]), .B2(n3392), 
        .ZN(n17313) );
  MOAI22 U26219 ( .A1(n28978), .A2(n3391), .B1(ram[13073]), .B2(n3392), 
        .ZN(n17314) );
  MOAI22 U26220 ( .A1(n28743), .A2(n3391), .B1(ram[13074]), .B2(n3392), 
        .ZN(n17315) );
  MOAI22 U26221 ( .A1(n28508), .A2(n3391), .B1(ram[13075]), .B2(n3392), 
        .ZN(n17316) );
  MOAI22 U26222 ( .A1(n28273), .A2(n3391), .B1(ram[13076]), .B2(n3392), 
        .ZN(n17317) );
  MOAI22 U26223 ( .A1(n28038), .A2(n3391), .B1(ram[13077]), .B2(n3392), 
        .ZN(n17318) );
  MOAI22 U26224 ( .A1(n27803), .A2(n3391), .B1(ram[13078]), .B2(n3392), 
        .ZN(n17319) );
  MOAI22 U26225 ( .A1(n27568), .A2(n3391), .B1(ram[13079]), .B2(n3392), 
        .ZN(n17320) );
  MOAI22 U26226 ( .A1(n29213), .A2(n3393), .B1(ram[13080]), .B2(n3394), 
        .ZN(n17321) );
  MOAI22 U26227 ( .A1(n28978), .A2(n3393), .B1(ram[13081]), .B2(n3394), 
        .ZN(n17322) );
  MOAI22 U26228 ( .A1(n28743), .A2(n3393), .B1(ram[13082]), .B2(n3394), 
        .ZN(n17323) );
  MOAI22 U26229 ( .A1(n28508), .A2(n3393), .B1(ram[13083]), .B2(n3394), 
        .ZN(n17324) );
  MOAI22 U26230 ( .A1(n28273), .A2(n3393), .B1(ram[13084]), .B2(n3394), 
        .ZN(n17325) );
  MOAI22 U26231 ( .A1(n28038), .A2(n3393), .B1(ram[13085]), .B2(n3394), 
        .ZN(n17326) );
  MOAI22 U26232 ( .A1(n27803), .A2(n3393), .B1(ram[13086]), .B2(n3394), 
        .ZN(n17327) );
  MOAI22 U26233 ( .A1(n27568), .A2(n3393), .B1(ram[13087]), .B2(n3394), 
        .ZN(n17328) );
  MOAI22 U26234 ( .A1(n29213), .A2(n3395), .B1(ram[13088]), .B2(n3396), 
        .ZN(n17329) );
  MOAI22 U26235 ( .A1(n28978), .A2(n3395), .B1(ram[13089]), .B2(n3396), 
        .ZN(n17330) );
  MOAI22 U26236 ( .A1(n28743), .A2(n3395), .B1(ram[13090]), .B2(n3396), 
        .ZN(n17331) );
  MOAI22 U26237 ( .A1(n28508), .A2(n3395), .B1(ram[13091]), .B2(n3396), 
        .ZN(n17332) );
  MOAI22 U26238 ( .A1(n28273), .A2(n3395), .B1(ram[13092]), .B2(n3396), 
        .ZN(n17333) );
  MOAI22 U26239 ( .A1(n28038), .A2(n3395), .B1(ram[13093]), .B2(n3396), 
        .ZN(n17334) );
  MOAI22 U26240 ( .A1(n27803), .A2(n3395), .B1(ram[13094]), .B2(n3396), 
        .ZN(n17335) );
  MOAI22 U26241 ( .A1(n27568), .A2(n3395), .B1(ram[13095]), .B2(n3396), 
        .ZN(n17336) );
  MOAI22 U26242 ( .A1(n29213), .A2(n3397), .B1(ram[13096]), .B2(n3398), 
        .ZN(n17337) );
  MOAI22 U26243 ( .A1(n28978), .A2(n3397), .B1(ram[13097]), .B2(n3398), 
        .ZN(n17338) );
  MOAI22 U26244 ( .A1(n28743), .A2(n3397), .B1(ram[13098]), .B2(n3398), 
        .ZN(n17339) );
  MOAI22 U26245 ( .A1(n28508), .A2(n3397), .B1(ram[13099]), .B2(n3398), 
        .ZN(n17340) );
  MOAI22 U26246 ( .A1(n28273), .A2(n3397), .B1(ram[13100]), .B2(n3398), 
        .ZN(n17341) );
  MOAI22 U26247 ( .A1(n28038), .A2(n3397), .B1(ram[13101]), .B2(n3398), 
        .ZN(n17342) );
  MOAI22 U26248 ( .A1(n27803), .A2(n3397), .B1(ram[13102]), .B2(n3398), 
        .ZN(n17343) );
  MOAI22 U26249 ( .A1(n27568), .A2(n3397), .B1(ram[13103]), .B2(n3398), 
        .ZN(n17344) );
  MOAI22 U26250 ( .A1(n29214), .A2(n3399), .B1(ram[13104]), .B2(n3400), 
        .ZN(n17345) );
  MOAI22 U26251 ( .A1(n28979), .A2(n3399), .B1(ram[13105]), .B2(n3400), 
        .ZN(n17346) );
  MOAI22 U26252 ( .A1(n28744), .A2(n3399), .B1(ram[13106]), .B2(n3400), 
        .ZN(n17347) );
  MOAI22 U26253 ( .A1(n28509), .A2(n3399), .B1(ram[13107]), .B2(n3400), 
        .ZN(n17348) );
  MOAI22 U26254 ( .A1(n28274), .A2(n3399), .B1(ram[13108]), .B2(n3400), 
        .ZN(n17349) );
  MOAI22 U26255 ( .A1(n28039), .A2(n3399), .B1(ram[13109]), .B2(n3400), 
        .ZN(n17350) );
  MOAI22 U26256 ( .A1(n27804), .A2(n3399), .B1(ram[13110]), .B2(n3400), 
        .ZN(n17351) );
  MOAI22 U26257 ( .A1(n27569), .A2(n3399), .B1(ram[13111]), .B2(n3400), 
        .ZN(n17352) );
  MOAI22 U26258 ( .A1(n29214), .A2(n3401), .B1(ram[13112]), .B2(n3402), 
        .ZN(n17353) );
  MOAI22 U26259 ( .A1(n28979), .A2(n3401), .B1(ram[13113]), .B2(n3402), 
        .ZN(n17354) );
  MOAI22 U26260 ( .A1(n28744), .A2(n3401), .B1(ram[13114]), .B2(n3402), 
        .ZN(n17355) );
  MOAI22 U26261 ( .A1(n28509), .A2(n3401), .B1(ram[13115]), .B2(n3402), 
        .ZN(n17356) );
  MOAI22 U26262 ( .A1(n28274), .A2(n3401), .B1(ram[13116]), .B2(n3402), 
        .ZN(n17357) );
  MOAI22 U26263 ( .A1(n28039), .A2(n3401), .B1(ram[13117]), .B2(n3402), 
        .ZN(n17358) );
  MOAI22 U26264 ( .A1(n27804), .A2(n3401), .B1(ram[13118]), .B2(n3402), 
        .ZN(n17359) );
  MOAI22 U26265 ( .A1(n27569), .A2(n3401), .B1(ram[13119]), .B2(n3402), 
        .ZN(n17360) );
  MOAI22 U26266 ( .A1(n29214), .A2(n3403), .B1(ram[13120]), .B2(n3404), 
        .ZN(n17361) );
  MOAI22 U26267 ( .A1(n28979), .A2(n3403), .B1(ram[13121]), .B2(n3404), 
        .ZN(n17362) );
  MOAI22 U26268 ( .A1(n28744), .A2(n3403), .B1(ram[13122]), .B2(n3404), 
        .ZN(n17363) );
  MOAI22 U26269 ( .A1(n28509), .A2(n3403), .B1(ram[13123]), .B2(n3404), 
        .ZN(n17364) );
  MOAI22 U26270 ( .A1(n28274), .A2(n3403), .B1(ram[13124]), .B2(n3404), 
        .ZN(n17365) );
  MOAI22 U26271 ( .A1(n28039), .A2(n3403), .B1(ram[13125]), .B2(n3404), 
        .ZN(n17366) );
  MOAI22 U26272 ( .A1(n27804), .A2(n3403), .B1(ram[13126]), .B2(n3404), 
        .ZN(n17367) );
  MOAI22 U26273 ( .A1(n27569), .A2(n3403), .B1(ram[13127]), .B2(n3404), 
        .ZN(n17368) );
  MOAI22 U26274 ( .A1(n29214), .A2(n3405), .B1(ram[13128]), .B2(n3406), 
        .ZN(n17369) );
  MOAI22 U26275 ( .A1(n28979), .A2(n3405), .B1(ram[13129]), .B2(n3406), 
        .ZN(n17370) );
  MOAI22 U26276 ( .A1(n28744), .A2(n3405), .B1(ram[13130]), .B2(n3406), 
        .ZN(n17371) );
  MOAI22 U26277 ( .A1(n28509), .A2(n3405), .B1(ram[13131]), .B2(n3406), 
        .ZN(n17372) );
  MOAI22 U26278 ( .A1(n28274), .A2(n3405), .B1(ram[13132]), .B2(n3406), 
        .ZN(n17373) );
  MOAI22 U26279 ( .A1(n28039), .A2(n3405), .B1(ram[13133]), .B2(n3406), 
        .ZN(n17374) );
  MOAI22 U26280 ( .A1(n27804), .A2(n3405), .B1(ram[13134]), .B2(n3406), 
        .ZN(n17375) );
  MOAI22 U26281 ( .A1(n27569), .A2(n3405), .B1(ram[13135]), .B2(n3406), 
        .ZN(n17376) );
  MOAI22 U26282 ( .A1(n29214), .A2(n3407), .B1(ram[13136]), .B2(n3408), 
        .ZN(n17377) );
  MOAI22 U26283 ( .A1(n28979), .A2(n3407), .B1(ram[13137]), .B2(n3408), 
        .ZN(n17378) );
  MOAI22 U26284 ( .A1(n28744), .A2(n3407), .B1(ram[13138]), .B2(n3408), 
        .ZN(n17379) );
  MOAI22 U26285 ( .A1(n28509), .A2(n3407), .B1(ram[13139]), .B2(n3408), 
        .ZN(n17380) );
  MOAI22 U26286 ( .A1(n28274), .A2(n3407), .B1(ram[13140]), .B2(n3408), 
        .ZN(n17381) );
  MOAI22 U26287 ( .A1(n28039), .A2(n3407), .B1(ram[13141]), .B2(n3408), 
        .ZN(n17382) );
  MOAI22 U26288 ( .A1(n27804), .A2(n3407), .B1(ram[13142]), .B2(n3408), 
        .ZN(n17383) );
  MOAI22 U26289 ( .A1(n27569), .A2(n3407), .B1(ram[13143]), .B2(n3408), 
        .ZN(n17384) );
  MOAI22 U26290 ( .A1(n29214), .A2(n3409), .B1(ram[13144]), .B2(n3410), 
        .ZN(n17385) );
  MOAI22 U26291 ( .A1(n28979), .A2(n3409), .B1(ram[13145]), .B2(n3410), 
        .ZN(n17386) );
  MOAI22 U26292 ( .A1(n28744), .A2(n3409), .B1(ram[13146]), .B2(n3410), 
        .ZN(n17387) );
  MOAI22 U26293 ( .A1(n28509), .A2(n3409), .B1(ram[13147]), .B2(n3410), 
        .ZN(n17388) );
  MOAI22 U26294 ( .A1(n28274), .A2(n3409), .B1(ram[13148]), .B2(n3410), 
        .ZN(n17389) );
  MOAI22 U26295 ( .A1(n28039), .A2(n3409), .B1(ram[13149]), .B2(n3410), 
        .ZN(n17390) );
  MOAI22 U26296 ( .A1(n27804), .A2(n3409), .B1(ram[13150]), .B2(n3410), 
        .ZN(n17391) );
  MOAI22 U26297 ( .A1(n27569), .A2(n3409), .B1(ram[13151]), .B2(n3410), 
        .ZN(n17392) );
  MOAI22 U26298 ( .A1(n29214), .A2(n3411), .B1(ram[13152]), .B2(n3412), 
        .ZN(n17393) );
  MOAI22 U26299 ( .A1(n28979), .A2(n3411), .B1(ram[13153]), .B2(n3412), 
        .ZN(n17394) );
  MOAI22 U26300 ( .A1(n28744), .A2(n3411), .B1(ram[13154]), .B2(n3412), 
        .ZN(n17395) );
  MOAI22 U26301 ( .A1(n28509), .A2(n3411), .B1(ram[13155]), .B2(n3412), 
        .ZN(n17396) );
  MOAI22 U26302 ( .A1(n28274), .A2(n3411), .B1(ram[13156]), .B2(n3412), 
        .ZN(n17397) );
  MOAI22 U26303 ( .A1(n28039), .A2(n3411), .B1(ram[13157]), .B2(n3412), 
        .ZN(n17398) );
  MOAI22 U26304 ( .A1(n27804), .A2(n3411), .B1(ram[13158]), .B2(n3412), 
        .ZN(n17399) );
  MOAI22 U26305 ( .A1(n27569), .A2(n3411), .B1(ram[13159]), .B2(n3412), 
        .ZN(n17400) );
  MOAI22 U26306 ( .A1(n29214), .A2(n3413), .B1(ram[13160]), .B2(n3414), 
        .ZN(n17401) );
  MOAI22 U26307 ( .A1(n28979), .A2(n3413), .B1(ram[13161]), .B2(n3414), 
        .ZN(n17402) );
  MOAI22 U26308 ( .A1(n28744), .A2(n3413), .B1(ram[13162]), .B2(n3414), 
        .ZN(n17403) );
  MOAI22 U26309 ( .A1(n28509), .A2(n3413), .B1(ram[13163]), .B2(n3414), 
        .ZN(n17404) );
  MOAI22 U26310 ( .A1(n28274), .A2(n3413), .B1(ram[13164]), .B2(n3414), 
        .ZN(n17405) );
  MOAI22 U26311 ( .A1(n28039), .A2(n3413), .B1(ram[13165]), .B2(n3414), 
        .ZN(n17406) );
  MOAI22 U26312 ( .A1(n27804), .A2(n3413), .B1(ram[13166]), .B2(n3414), 
        .ZN(n17407) );
  MOAI22 U26313 ( .A1(n27569), .A2(n3413), .B1(ram[13167]), .B2(n3414), 
        .ZN(n17408) );
  MOAI22 U26314 ( .A1(n29214), .A2(n3415), .B1(ram[13168]), .B2(n3416), 
        .ZN(n17409) );
  MOAI22 U26315 ( .A1(n28979), .A2(n3415), .B1(ram[13169]), .B2(n3416), 
        .ZN(n17410) );
  MOAI22 U26316 ( .A1(n28744), .A2(n3415), .B1(ram[13170]), .B2(n3416), 
        .ZN(n17411) );
  MOAI22 U26317 ( .A1(n28509), .A2(n3415), .B1(ram[13171]), .B2(n3416), 
        .ZN(n17412) );
  MOAI22 U26318 ( .A1(n28274), .A2(n3415), .B1(ram[13172]), .B2(n3416), 
        .ZN(n17413) );
  MOAI22 U26319 ( .A1(n28039), .A2(n3415), .B1(ram[13173]), .B2(n3416), 
        .ZN(n17414) );
  MOAI22 U26320 ( .A1(n27804), .A2(n3415), .B1(ram[13174]), .B2(n3416), 
        .ZN(n17415) );
  MOAI22 U26321 ( .A1(n27569), .A2(n3415), .B1(ram[13175]), .B2(n3416), 
        .ZN(n17416) );
  MOAI22 U26322 ( .A1(n29214), .A2(n3417), .B1(ram[13176]), .B2(n3418), 
        .ZN(n17417) );
  MOAI22 U26323 ( .A1(n28979), .A2(n3417), .B1(ram[13177]), .B2(n3418), 
        .ZN(n17418) );
  MOAI22 U26324 ( .A1(n28744), .A2(n3417), .B1(ram[13178]), .B2(n3418), 
        .ZN(n17419) );
  MOAI22 U26325 ( .A1(n28509), .A2(n3417), .B1(ram[13179]), .B2(n3418), 
        .ZN(n17420) );
  MOAI22 U26326 ( .A1(n28274), .A2(n3417), .B1(ram[13180]), .B2(n3418), 
        .ZN(n17421) );
  MOAI22 U26327 ( .A1(n28039), .A2(n3417), .B1(ram[13181]), .B2(n3418), 
        .ZN(n17422) );
  MOAI22 U26328 ( .A1(n27804), .A2(n3417), .B1(ram[13182]), .B2(n3418), 
        .ZN(n17423) );
  MOAI22 U26329 ( .A1(n27569), .A2(n3417), .B1(ram[13183]), .B2(n3418), 
        .ZN(n17424) );
  MOAI22 U26330 ( .A1(n29214), .A2(n3419), .B1(ram[13184]), .B2(n3420), 
        .ZN(n17425) );
  MOAI22 U26331 ( .A1(n28979), .A2(n3419), .B1(ram[13185]), .B2(n3420), 
        .ZN(n17426) );
  MOAI22 U26332 ( .A1(n28744), .A2(n3419), .B1(ram[13186]), .B2(n3420), 
        .ZN(n17427) );
  MOAI22 U26333 ( .A1(n28509), .A2(n3419), .B1(ram[13187]), .B2(n3420), 
        .ZN(n17428) );
  MOAI22 U26334 ( .A1(n28274), .A2(n3419), .B1(ram[13188]), .B2(n3420), 
        .ZN(n17429) );
  MOAI22 U26335 ( .A1(n28039), .A2(n3419), .B1(ram[13189]), .B2(n3420), 
        .ZN(n17430) );
  MOAI22 U26336 ( .A1(n27804), .A2(n3419), .B1(ram[13190]), .B2(n3420), 
        .ZN(n17431) );
  MOAI22 U26337 ( .A1(n27569), .A2(n3419), .B1(ram[13191]), .B2(n3420), 
        .ZN(n17432) );
  MOAI22 U26338 ( .A1(n29214), .A2(n3421), .B1(ram[13192]), .B2(n3422), 
        .ZN(n17433) );
  MOAI22 U26339 ( .A1(n28979), .A2(n3421), .B1(ram[13193]), .B2(n3422), 
        .ZN(n17434) );
  MOAI22 U26340 ( .A1(n28744), .A2(n3421), .B1(ram[13194]), .B2(n3422), 
        .ZN(n17435) );
  MOAI22 U26341 ( .A1(n28509), .A2(n3421), .B1(ram[13195]), .B2(n3422), 
        .ZN(n17436) );
  MOAI22 U26342 ( .A1(n28274), .A2(n3421), .B1(ram[13196]), .B2(n3422), 
        .ZN(n17437) );
  MOAI22 U26343 ( .A1(n28039), .A2(n3421), .B1(ram[13197]), .B2(n3422), 
        .ZN(n17438) );
  MOAI22 U26344 ( .A1(n27804), .A2(n3421), .B1(ram[13198]), .B2(n3422), 
        .ZN(n17439) );
  MOAI22 U26345 ( .A1(n27569), .A2(n3421), .B1(ram[13199]), .B2(n3422), 
        .ZN(n17440) );
  MOAI22 U26346 ( .A1(n29214), .A2(n3423), .B1(ram[13200]), .B2(n3424), 
        .ZN(n17441) );
  MOAI22 U26347 ( .A1(n28979), .A2(n3423), .B1(ram[13201]), .B2(n3424), 
        .ZN(n17442) );
  MOAI22 U26348 ( .A1(n28744), .A2(n3423), .B1(ram[13202]), .B2(n3424), 
        .ZN(n17443) );
  MOAI22 U26349 ( .A1(n28509), .A2(n3423), .B1(ram[13203]), .B2(n3424), 
        .ZN(n17444) );
  MOAI22 U26350 ( .A1(n28274), .A2(n3423), .B1(ram[13204]), .B2(n3424), 
        .ZN(n17445) );
  MOAI22 U26351 ( .A1(n28039), .A2(n3423), .B1(ram[13205]), .B2(n3424), 
        .ZN(n17446) );
  MOAI22 U26352 ( .A1(n27804), .A2(n3423), .B1(ram[13206]), .B2(n3424), 
        .ZN(n17447) );
  MOAI22 U26353 ( .A1(n27569), .A2(n3423), .B1(ram[13207]), .B2(n3424), 
        .ZN(n17448) );
  MOAI22 U26354 ( .A1(n29215), .A2(n3425), .B1(ram[13208]), .B2(n3426), 
        .ZN(n17449) );
  MOAI22 U26355 ( .A1(n28980), .A2(n3425), .B1(ram[13209]), .B2(n3426), 
        .ZN(n17450) );
  MOAI22 U26356 ( .A1(n28745), .A2(n3425), .B1(ram[13210]), .B2(n3426), 
        .ZN(n17451) );
  MOAI22 U26357 ( .A1(n28510), .A2(n3425), .B1(ram[13211]), .B2(n3426), 
        .ZN(n17452) );
  MOAI22 U26358 ( .A1(n28275), .A2(n3425), .B1(ram[13212]), .B2(n3426), 
        .ZN(n17453) );
  MOAI22 U26359 ( .A1(n28040), .A2(n3425), .B1(ram[13213]), .B2(n3426), 
        .ZN(n17454) );
  MOAI22 U26360 ( .A1(n27805), .A2(n3425), .B1(ram[13214]), .B2(n3426), 
        .ZN(n17455) );
  MOAI22 U26361 ( .A1(n27570), .A2(n3425), .B1(ram[13215]), .B2(n3426), 
        .ZN(n17456) );
  MOAI22 U26362 ( .A1(n29215), .A2(n3427), .B1(ram[13216]), .B2(n3428), 
        .ZN(n17457) );
  MOAI22 U26363 ( .A1(n28980), .A2(n3427), .B1(ram[13217]), .B2(n3428), 
        .ZN(n17458) );
  MOAI22 U26364 ( .A1(n28745), .A2(n3427), .B1(ram[13218]), .B2(n3428), 
        .ZN(n17459) );
  MOAI22 U26365 ( .A1(n28510), .A2(n3427), .B1(ram[13219]), .B2(n3428), 
        .ZN(n17460) );
  MOAI22 U26366 ( .A1(n28275), .A2(n3427), .B1(ram[13220]), .B2(n3428), 
        .ZN(n17461) );
  MOAI22 U26367 ( .A1(n28040), .A2(n3427), .B1(ram[13221]), .B2(n3428), 
        .ZN(n17462) );
  MOAI22 U26368 ( .A1(n27805), .A2(n3427), .B1(ram[13222]), .B2(n3428), 
        .ZN(n17463) );
  MOAI22 U26369 ( .A1(n27570), .A2(n3427), .B1(ram[13223]), .B2(n3428), 
        .ZN(n17464) );
  MOAI22 U26370 ( .A1(n29215), .A2(n3429), .B1(ram[13224]), .B2(n3430), 
        .ZN(n17465) );
  MOAI22 U26371 ( .A1(n28980), .A2(n3429), .B1(ram[13225]), .B2(n3430), 
        .ZN(n17466) );
  MOAI22 U26372 ( .A1(n28745), .A2(n3429), .B1(ram[13226]), .B2(n3430), 
        .ZN(n17467) );
  MOAI22 U26373 ( .A1(n28510), .A2(n3429), .B1(ram[13227]), .B2(n3430), 
        .ZN(n17468) );
  MOAI22 U26374 ( .A1(n28275), .A2(n3429), .B1(ram[13228]), .B2(n3430), 
        .ZN(n17469) );
  MOAI22 U26375 ( .A1(n28040), .A2(n3429), .B1(ram[13229]), .B2(n3430), 
        .ZN(n17470) );
  MOAI22 U26376 ( .A1(n27805), .A2(n3429), .B1(ram[13230]), .B2(n3430), 
        .ZN(n17471) );
  MOAI22 U26377 ( .A1(n27570), .A2(n3429), .B1(ram[13231]), .B2(n3430), 
        .ZN(n17472) );
  MOAI22 U26378 ( .A1(n29215), .A2(n3431), .B1(ram[13232]), .B2(n3432), 
        .ZN(n17473) );
  MOAI22 U26379 ( .A1(n28980), .A2(n3431), .B1(ram[13233]), .B2(n3432), 
        .ZN(n17474) );
  MOAI22 U26380 ( .A1(n28745), .A2(n3431), .B1(ram[13234]), .B2(n3432), 
        .ZN(n17475) );
  MOAI22 U26381 ( .A1(n28510), .A2(n3431), .B1(ram[13235]), .B2(n3432), 
        .ZN(n17476) );
  MOAI22 U26382 ( .A1(n28275), .A2(n3431), .B1(ram[13236]), .B2(n3432), 
        .ZN(n17477) );
  MOAI22 U26383 ( .A1(n28040), .A2(n3431), .B1(ram[13237]), .B2(n3432), 
        .ZN(n17478) );
  MOAI22 U26384 ( .A1(n27805), .A2(n3431), .B1(ram[13238]), .B2(n3432), 
        .ZN(n17479) );
  MOAI22 U26385 ( .A1(n27570), .A2(n3431), .B1(ram[13239]), .B2(n3432), 
        .ZN(n17480) );
  MOAI22 U26386 ( .A1(n29215), .A2(n3433), .B1(ram[13240]), .B2(n3434), 
        .ZN(n17481) );
  MOAI22 U26387 ( .A1(n28980), .A2(n3433), .B1(ram[13241]), .B2(n3434), 
        .ZN(n17482) );
  MOAI22 U26388 ( .A1(n28745), .A2(n3433), .B1(ram[13242]), .B2(n3434), 
        .ZN(n17483) );
  MOAI22 U26389 ( .A1(n28510), .A2(n3433), .B1(ram[13243]), .B2(n3434), 
        .ZN(n17484) );
  MOAI22 U26390 ( .A1(n28275), .A2(n3433), .B1(ram[13244]), .B2(n3434), 
        .ZN(n17485) );
  MOAI22 U26391 ( .A1(n28040), .A2(n3433), .B1(ram[13245]), .B2(n3434), 
        .ZN(n17486) );
  MOAI22 U26392 ( .A1(n27805), .A2(n3433), .B1(ram[13246]), .B2(n3434), 
        .ZN(n17487) );
  MOAI22 U26393 ( .A1(n27570), .A2(n3433), .B1(ram[13247]), .B2(n3434), 
        .ZN(n17488) );
  MOAI22 U26394 ( .A1(n29215), .A2(n3435), .B1(ram[13248]), .B2(n3436), 
        .ZN(n17489) );
  MOAI22 U26395 ( .A1(n28980), .A2(n3435), .B1(ram[13249]), .B2(n3436), 
        .ZN(n17490) );
  MOAI22 U26396 ( .A1(n28745), .A2(n3435), .B1(ram[13250]), .B2(n3436), 
        .ZN(n17491) );
  MOAI22 U26397 ( .A1(n28510), .A2(n3435), .B1(ram[13251]), .B2(n3436), 
        .ZN(n17492) );
  MOAI22 U26398 ( .A1(n28275), .A2(n3435), .B1(ram[13252]), .B2(n3436), 
        .ZN(n17493) );
  MOAI22 U26399 ( .A1(n28040), .A2(n3435), .B1(ram[13253]), .B2(n3436), 
        .ZN(n17494) );
  MOAI22 U26400 ( .A1(n27805), .A2(n3435), .B1(ram[13254]), .B2(n3436), 
        .ZN(n17495) );
  MOAI22 U26401 ( .A1(n27570), .A2(n3435), .B1(ram[13255]), .B2(n3436), 
        .ZN(n17496) );
  MOAI22 U26402 ( .A1(n29215), .A2(n3437), .B1(ram[13256]), .B2(n3438), 
        .ZN(n17497) );
  MOAI22 U26403 ( .A1(n28980), .A2(n3437), .B1(ram[13257]), .B2(n3438), 
        .ZN(n17498) );
  MOAI22 U26404 ( .A1(n28745), .A2(n3437), .B1(ram[13258]), .B2(n3438), 
        .ZN(n17499) );
  MOAI22 U26405 ( .A1(n28510), .A2(n3437), .B1(ram[13259]), .B2(n3438), 
        .ZN(n17500) );
  MOAI22 U26406 ( .A1(n28275), .A2(n3437), .B1(ram[13260]), .B2(n3438), 
        .ZN(n17501) );
  MOAI22 U26407 ( .A1(n28040), .A2(n3437), .B1(ram[13261]), .B2(n3438), 
        .ZN(n17502) );
  MOAI22 U26408 ( .A1(n27805), .A2(n3437), .B1(ram[13262]), .B2(n3438), 
        .ZN(n17503) );
  MOAI22 U26409 ( .A1(n27570), .A2(n3437), .B1(ram[13263]), .B2(n3438), 
        .ZN(n17504) );
  MOAI22 U26410 ( .A1(n29215), .A2(n3439), .B1(ram[13264]), .B2(n3440), 
        .ZN(n17505) );
  MOAI22 U26411 ( .A1(n28980), .A2(n3439), .B1(ram[13265]), .B2(n3440), 
        .ZN(n17506) );
  MOAI22 U26412 ( .A1(n28745), .A2(n3439), .B1(ram[13266]), .B2(n3440), 
        .ZN(n17507) );
  MOAI22 U26413 ( .A1(n28510), .A2(n3439), .B1(ram[13267]), .B2(n3440), 
        .ZN(n17508) );
  MOAI22 U26414 ( .A1(n28275), .A2(n3439), .B1(ram[13268]), .B2(n3440), 
        .ZN(n17509) );
  MOAI22 U26415 ( .A1(n28040), .A2(n3439), .B1(ram[13269]), .B2(n3440), 
        .ZN(n17510) );
  MOAI22 U26416 ( .A1(n27805), .A2(n3439), .B1(ram[13270]), .B2(n3440), 
        .ZN(n17511) );
  MOAI22 U26417 ( .A1(n27570), .A2(n3439), .B1(ram[13271]), .B2(n3440), 
        .ZN(n17512) );
  MOAI22 U26418 ( .A1(n29215), .A2(n3441), .B1(ram[13272]), .B2(n3442), 
        .ZN(n17513) );
  MOAI22 U26419 ( .A1(n28980), .A2(n3441), .B1(ram[13273]), .B2(n3442), 
        .ZN(n17514) );
  MOAI22 U26420 ( .A1(n28745), .A2(n3441), .B1(ram[13274]), .B2(n3442), 
        .ZN(n17515) );
  MOAI22 U26421 ( .A1(n28510), .A2(n3441), .B1(ram[13275]), .B2(n3442), 
        .ZN(n17516) );
  MOAI22 U26422 ( .A1(n28275), .A2(n3441), .B1(ram[13276]), .B2(n3442), 
        .ZN(n17517) );
  MOAI22 U26423 ( .A1(n28040), .A2(n3441), .B1(ram[13277]), .B2(n3442), 
        .ZN(n17518) );
  MOAI22 U26424 ( .A1(n27805), .A2(n3441), .B1(ram[13278]), .B2(n3442), 
        .ZN(n17519) );
  MOAI22 U26425 ( .A1(n27570), .A2(n3441), .B1(ram[13279]), .B2(n3442), 
        .ZN(n17520) );
  MOAI22 U26426 ( .A1(n29215), .A2(n3443), .B1(ram[13280]), .B2(n3444), 
        .ZN(n17521) );
  MOAI22 U26427 ( .A1(n28980), .A2(n3443), .B1(ram[13281]), .B2(n3444), 
        .ZN(n17522) );
  MOAI22 U26428 ( .A1(n28745), .A2(n3443), .B1(ram[13282]), .B2(n3444), 
        .ZN(n17523) );
  MOAI22 U26429 ( .A1(n28510), .A2(n3443), .B1(ram[13283]), .B2(n3444), 
        .ZN(n17524) );
  MOAI22 U26430 ( .A1(n28275), .A2(n3443), .B1(ram[13284]), .B2(n3444), 
        .ZN(n17525) );
  MOAI22 U26431 ( .A1(n28040), .A2(n3443), .B1(ram[13285]), .B2(n3444), 
        .ZN(n17526) );
  MOAI22 U26432 ( .A1(n27805), .A2(n3443), .B1(ram[13286]), .B2(n3444), 
        .ZN(n17527) );
  MOAI22 U26433 ( .A1(n27570), .A2(n3443), .B1(ram[13287]), .B2(n3444), 
        .ZN(n17528) );
  MOAI22 U26434 ( .A1(n29215), .A2(n3445), .B1(ram[13288]), .B2(n3446), 
        .ZN(n17529) );
  MOAI22 U26435 ( .A1(n28980), .A2(n3445), .B1(ram[13289]), .B2(n3446), 
        .ZN(n17530) );
  MOAI22 U26436 ( .A1(n28745), .A2(n3445), .B1(ram[13290]), .B2(n3446), 
        .ZN(n17531) );
  MOAI22 U26437 ( .A1(n28510), .A2(n3445), .B1(ram[13291]), .B2(n3446), 
        .ZN(n17532) );
  MOAI22 U26438 ( .A1(n28275), .A2(n3445), .B1(ram[13292]), .B2(n3446), 
        .ZN(n17533) );
  MOAI22 U26439 ( .A1(n28040), .A2(n3445), .B1(ram[13293]), .B2(n3446), 
        .ZN(n17534) );
  MOAI22 U26440 ( .A1(n27805), .A2(n3445), .B1(ram[13294]), .B2(n3446), 
        .ZN(n17535) );
  MOAI22 U26441 ( .A1(n27570), .A2(n3445), .B1(ram[13295]), .B2(n3446), 
        .ZN(n17536) );
  MOAI22 U26442 ( .A1(n29215), .A2(n3447), .B1(ram[13296]), .B2(n3448), 
        .ZN(n17537) );
  MOAI22 U26443 ( .A1(n28980), .A2(n3447), .B1(ram[13297]), .B2(n3448), 
        .ZN(n17538) );
  MOAI22 U26444 ( .A1(n28745), .A2(n3447), .B1(ram[13298]), .B2(n3448), 
        .ZN(n17539) );
  MOAI22 U26445 ( .A1(n28510), .A2(n3447), .B1(ram[13299]), .B2(n3448), 
        .ZN(n17540) );
  MOAI22 U26446 ( .A1(n28275), .A2(n3447), .B1(ram[13300]), .B2(n3448), 
        .ZN(n17541) );
  MOAI22 U26447 ( .A1(n28040), .A2(n3447), .B1(ram[13301]), .B2(n3448), 
        .ZN(n17542) );
  MOAI22 U26448 ( .A1(n27805), .A2(n3447), .B1(ram[13302]), .B2(n3448), 
        .ZN(n17543) );
  MOAI22 U26449 ( .A1(n27570), .A2(n3447), .B1(ram[13303]), .B2(n3448), 
        .ZN(n17544) );
  MOAI22 U26450 ( .A1(n29215), .A2(n3449), .B1(ram[13304]), .B2(n3450), 
        .ZN(n17545) );
  MOAI22 U26451 ( .A1(n28980), .A2(n3449), .B1(ram[13305]), .B2(n3450), 
        .ZN(n17546) );
  MOAI22 U26452 ( .A1(n28745), .A2(n3449), .B1(ram[13306]), .B2(n3450), 
        .ZN(n17547) );
  MOAI22 U26453 ( .A1(n28510), .A2(n3449), .B1(ram[13307]), .B2(n3450), 
        .ZN(n17548) );
  MOAI22 U26454 ( .A1(n28275), .A2(n3449), .B1(ram[13308]), .B2(n3450), 
        .ZN(n17549) );
  MOAI22 U26455 ( .A1(n28040), .A2(n3449), .B1(ram[13309]), .B2(n3450), 
        .ZN(n17550) );
  MOAI22 U26456 ( .A1(n27805), .A2(n3449), .B1(ram[13310]), .B2(n3450), 
        .ZN(n17551) );
  MOAI22 U26457 ( .A1(n27570), .A2(n3449), .B1(ram[13311]), .B2(n3450), 
        .ZN(n17552) );
  MOAI22 U26458 ( .A1(n29216), .A2(n3451), .B1(ram[13312]), .B2(n3452), 
        .ZN(n17553) );
  MOAI22 U26459 ( .A1(n28981), .A2(n3451), .B1(ram[13313]), .B2(n3452), 
        .ZN(n17554) );
  MOAI22 U26460 ( .A1(n28746), .A2(n3451), .B1(ram[13314]), .B2(n3452), 
        .ZN(n17555) );
  MOAI22 U26461 ( .A1(n28511), .A2(n3451), .B1(ram[13315]), .B2(n3452), 
        .ZN(n17556) );
  MOAI22 U26462 ( .A1(n28276), .A2(n3451), .B1(ram[13316]), .B2(n3452), 
        .ZN(n17557) );
  MOAI22 U26463 ( .A1(n28041), .A2(n3451), .B1(ram[13317]), .B2(n3452), 
        .ZN(n17558) );
  MOAI22 U26464 ( .A1(n27806), .A2(n3451), .B1(ram[13318]), .B2(n3452), 
        .ZN(n17559) );
  MOAI22 U26465 ( .A1(n27571), .A2(n3451), .B1(ram[13319]), .B2(n3452), 
        .ZN(n17560) );
  MOAI22 U26466 ( .A1(n29216), .A2(n3454), .B1(ram[13320]), .B2(n3455), 
        .ZN(n17561) );
  MOAI22 U26467 ( .A1(n28981), .A2(n3454), .B1(ram[13321]), .B2(n3455), 
        .ZN(n17562) );
  MOAI22 U26468 ( .A1(n28746), .A2(n3454), .B1(ram[13322]), .B2(n3455), 
        .ZN(n17563) );
  MOAI22 U26469 ( .A1(n28511), .A2(n3454), .B1(ram[13323]), .B2(n3455), 
        .ZN(n17564) );
  MOAI22 U26470 ( .A1(n28276), .A2(n3454), .B1(ram[13324]), .B2(n3455), 
        .ZN(n17565) );
  MOAI22 U26471 ( .A1(n28041), .A2(n3454), .B1(ram[13325]), .B2(n3455), 
        .ZN(n17566) );
  MOAI22 U26472 ( .A1(n27806), .A2(n3454), .B1(ram[13326]), .B2(n3455), 
        .ZN(n17567) );
  MOAI22 U26473 ( .A1(n27571), .A2(n3454), .B1(ram[13327]), .B2(n3455), 
        .ZN(n17568) );
  MOAI22 U26474 ( .A1(n29216), .A2(n3456), .B1(ram[13328]), .B2(n3457), 
        .ZN(n17569) );
  MOAI22 U26475 ( .A1(n28981), .A2(n3456), .B1(ram[13329]), .B2(n3457), 
        .ZN(n17570) );
  MOAI22 U26476 ( .A1(n28746), .A2(n3456), .B1(ram[13330]), .B2(n3457), 
        .ZN(n17571) );
  MOAI22 U26477 ( .A1(n28511), .A2(n3456), .B1(ram[13331]), .B2(n3457), 
        .ZN(n17572) );
  MOAI22 U26478 ( .A1(n28276), .A2(n3456), .B1(ram[13332]), .B2(n3457), 
        .ZN(n17573) );
  MOAI22 U26479 ( .A1(n28041), .A2(n3456), .B1(ram[13333]), .B2(n3457), 
        .ZN(n17574) );
  MOAI22 U26480 ( .A1(n27806), .A2(n3456), .B1(ram[13334]), .B2(n3457), 
        .ZN(n17575) );
  MOAI22 U26481 ( .A1(n27571), .A2(n3456), .B1(ram[13335]), .B2(n3457), 
        .ZN(n17576) );
  MOAI22 U26482 ( .A1(n29216), .A2(n3458), .B1(ram[13336]), .B2(n3459), 
        .ZN(n17577) );
  MOAI22 U26483 ( .A1(n28981), .A2(n3458), .B1(ram[13337]), .B2(n3459), 
        .ZN(n17578) );
  MOAI22 U26484 ( .A1(n28746), .A2(n3458), .B1(ram[13338]), .B2(n3459), 
        .ZN(n17579) );
  MOAI22 U26485 ( .A1(n28511), .A2(n3458), .B1(ram[13339]), .B2(n3459), 
        .ZN(n17580) );
  MOAI22 U26486 ( .A1(n28276), .A2(n3458), .B1(ram[13340]), .B2(n3459), 
        .ZN(n17581) );
  MOAI22 U26487 ( .A1(n28041), .A2(n3458), .B1(ram[13341]), .B2(n3459), 
        .ZN(n17582) );
  MOAI22 U26488 ( .A1(n27806), .A2(n3458), .B1(ram[13342]), .B2(n3459), 
        .ZN(n17583) );
  MOAI22 U26489 ( .A1(n27571), .A2(n3458), .B1(ram[13343]), .B2(n3459), 
        .ZN(n17584) );
  MOAI22 U26490 ( .A1(n29216), .A2(n3460), .B1(ram[13344]), .B2(n3461), 
        .ZN(n17585) );
  MOAI22 U26491 ( .A1(n28981), .A2(n3460), .B1(ram[13345]), .B2(n3461), 
        .ZN(n17586) );
  MOAI22 U26492 ( .A1(n28746), .A2(n3460), .B1(ram[13346]), .B2(n3461), 
        .ZN(n17587) );
  MOAI22 U26493 ( .A1(n28511), .A2(n3460), .B1(ram[13347]), .B2(n3461), 
        .ZN(n17588) );
  MOAI22 U26494 ( .A1(n28276), .A2(n3460), .B1(ram[13348]), .B2(n3461), 
        .ZN(n17589) );
  MOAI22 U26495 ( .A1(n28041), .A2(n3460), .B1(ram[13349]), .B2(n3461), 
        .ZN(n17590) );
  MOAI22 U26496 ( .A1(n27806), .A2(n3460), .B1(ram[13350]), .B2(n3461), 
        .ZN(n17591) );
  MOAI22 U26497 ( .A1(n27571), .A2(n3460), .B1(ram[13351]), .B2(n3461), 
        .ZN(n17592) );
  MOAI22 U26498 ( .A1(n29216), .A2(n3462), .B1(ram[13352]), .B2(n3463), 
        .ZN(n17593) );
  MOAI22 U26499 ( .A1(n28981), .A2(n3462), .B1(ram[13353]), .B2(n3463), 
        .ZN(n17594) );
  MOAI22 U26500 ( .A1(n28746), .A2(n3462), .B1(ram[13354]), .B2(n3463), 
        .ZN(n17595) );
  MOAI22 U26501 ( .A1(n28511), .A2(n3462), .B1(ram[13355]), .B2(n3463), 
        .ZN(n17596) );
  MOAI22 U26502 ( .A1(n28276), .A2(n3462), .B1(ram[13356]), .B2(n3463), 
        .ZN(n17597) );
  MOAI22 U26503 ( .A1(n28041), .A2(n3462), .B1(ram[13357]), .B2(n3463), 
        .ZN(n17598) );
  MOAI22 U26504 ( .A1(n27806), .A2(n3462), .B1(ram[13358]), .B2(n3463), 
        .ZN(n17599) );
  MOAI22 U26505 ( .A1(n27571), .A2(n3462), .B1(ram[13359]), .B2(n3463), 
        .ZN(n17600) );
  MOAI22 U26506 ( .A1(n29216), .A2(n3464), .B1(ram[13360]), .B2(n3465), 
        .ZN(n17601) );
  MOAI22 U26507 ( .A1(n28981), .A2(n3464), .B1(ram[13361]), .B2(n3465), 
        .ZN(n17602) );
  MOAI22 U26508 ( .A1(n28746), .A2(n3464), .B1(ram[13362]), .B2(n3465), 
        .ZN(n17603) );
  MOAI22 U26509 ( .A1(n28511), .A2(n3464), .B1(ram[13363]), .B2(n3465), 
        .ZN(n17604) );
  MOAI22 U26510 ( .A1(n28276), .A2(n3464), .B1(ram[13364]), .B2(n3465), 
        .ZN(n17605) );
  MOAI22 U26511 ( .A1(n28041), .A2(n3464), .B1(ram[13365]), .B2(n3465), 
        .ZN(n17606) );
  MOAI22 U26512 ( .A1(n27806), .A2(n3464), .B1(ram[13366]), .B2(n3465), 
        .ZN(n17607) );
  MOAI22 U26513 ( .A1(n27571), .A2(n3464), .B1(ram[13367]), .B2(n3465), 
        .ZN(n17608) );
  MOAI22 U26514 ( .A1(n29216), .A2(n3466), .B1(ram[13368]), .B2(n3467), 
        .ZN(n17609) );
  MOAI22 U26515 ( .A1(n28981), .A2(n3466), .B1(ram[13369]), .B2(n3467), 
        .ZN(n17610) );
  MOAI22 U26516 ( .A1(n28746), .A2(n3466), .B1(ram[13370]), .B2(n3467), 
        .ZN(n17611) );
  MOAI22 U26517 ( .A1(n28511), .A2(n3466), .B1(ram[13371]), .B2(n3467), 
        .ZN(n17612) );
  MOAI22 U26518 ( .A1(n28276), .A2(n3466), .B1(ram[13372]), .B2(n3467), 
        .ZN(n17613) );
  MOAI22 U26519 ( .A1(n28041), .A2(n3466), .B1(ram[13373]), .B2(n3467), 
        .ZN(n17614) );
  MOAI22 U26520 ( .A1(n27806), .A2(n3466), .B1(ram[13374]), .B2(n3467), 
        .ZN(n17615) );
  MOAI22 U26521 ( .A1(n27571), .A2(n3466), .B1(ram[13375]), .B2(n3467), 
        .ZN(n17616) );
  MOAI22 U26522 ( .A1(n29216), .A2(n3468), .B1(ram[13376]), .B2(n3469), 
        .ZN(n17617) );
  MOAI22 U26523 ( .A1(n28981), .A2(n3468), .B1(ram[13377]), .B2(n3469), 
        .ZN(n17618) );
  MOAI22 U26524 ( .A1(n28746), .A2(n3468), .B1(ram[13378]), .B2(n3469), 
        .ZN(n17619) );
  MOAI22 U26525 ( .A1(n28511), .A2(n3468), .B1(ram[13379]), .B2(n3469), 
        .ZN(n17620) );
  MOAI22 U26526 ( .A1(n28276), .A2(n3468), .B1(ram[13380]), .B2(n3469), 
        .ZN(n17621) );
  MOAI22 U26527 ( .A1(n28041), .A2(n3468), .B1(ram[13381]), .B2(n3469), 
        .ZN(n17622) );
  MOAI22 U26528 ( .A1(n27806), .A2(n3468), .B1(ram[13382]), .B2(n3469), 
        .ZN(n17623) );
  MOAI22 U26529 ( .A1(n27571), .A2(n3468), .B1(ram[13383]), .B2(n3469), 
        .ZN(n17624) );
  MOAI22 U26530 ( .A1(n29216), .A2(n3470), .B1(ram[13384]), .B2(n3471), 
        .ZN(n17625) );
  MOAI22 U26531 ( .A1(n28981), .A2(n3470), .B1(ram[13385]), .B2(n3471), 
        .ZN(n17626) );
  MOAI22 U26532 ( .A1(n28746), .A2(n3470), .B1(ram[13386]), .B2(n3471), 
        .ZN(n17627) );
  MOAI22 U26533 ( .A1(n28511), .A2(n3470), .B1(ram[13387]), .B2(n3471), 
        .ZN(n17628) );
  MOAI22 U26534 ( .A1(n28276), .A2(n3470), .B1(ram[13388]), .B2(n3471), 
        .ZN(n17629) );
  MOAI22 U26535 ( .A1(n28041), .A2(n3470), .B1(ram[13389]), .B2(n3471), 
        .ZN(n17630) );
  MOAI22 U26536 ( .A1(n27806), .A2(n3470), .B1(ram[13390]), .B2(n3471), 
        .ZN(n17631) );
  MOAI22 U26537 ( .A1(n27571), .A2(n3470), .B1(ram[13391]), .B2(n3471), 
        .ZN(n17632) );
  MOAI22 U26538 ( .A1(n29216), .A2(n3472), .B1(ram[13392]), .B2(n3473), 
        .ZN(n17633) );
  MOAI22 U26539 ( .A1(n28981), .A2(n3472), .B1(ram[13393]), .B2(n3473), 
        .ZN(n17634) );
  MOAI22 U26540 ( .A1(n28746), .A2(n3472), .B1(ram[13394]), .B2(n3473), 
        .ZN(n17635) );
  MOAI22 U26541 ( .A1(n28511), .A2(n3472), .B1(ram[13395]), .B2(n3473), 
        .ZN(n17636) );
  MOAI22 U26542 ( .A1(n28276), .A2(n3472), .B1(ram[13396]), .B2(n3473), 
        .ZN(n17637) );
  MOAI22 U26543 ( .A1(n28041), .A2(n3472), .B1(ram[13397]), .B2(n3473), 
        .ZN(n17638) );
  MOAI22 U26544 ( .A1(n27806), .A2(n3472), .B1(ram[13398]), .B2(n3473), 
        .ZN(n17639) );
  MOAI22 U26545 ( .A1(n27571), .A2(n3472), .B1(ram[13399]), .B2(n3473), 
        .ZN(n17640) );
  MOAI22 U26546 ( .A1(n29216), .A2(n3474), .B1(ram[13400]), .B2(n3475), 
        .ZN(n17641) );
  MOAI22 U26547 ( .A1(n28981), .A2(n3474), .B1(ram[13401]), .B2(n3475), 
        .ZN(n17642) );
  MOAI22 U26548 ( .A1(n28746), .A2(n3474), .B1(ram[13402]), .B2(n3475), 
        .ZN(n17643) );
  MOAI22 U26549 ( .A1(n28511), .A2(n3474), .B1(ram[13403]), .B2(n3475), 
        .ZN(n17644) );
  MOAI22 U26550 ( .A1(n28276), .A2(n3474), .B1(ram[13404]), .B2(n3475), 
        .ZN(n17645) );
  MOAI22 U26551 ( .A1(n28041), .A2(n3474), .B1(ram[13405]), .B2(n3475), 
        .ZN(n17646) );
  MOAI22 U26552 ( .A1(n27806), .A2(n3474), .B1(ram[13406]), .B2(n3475), 
        .ZN(n17647) );
  MOAI22 U26553 ( .A1(n27571), .A2(n3474), .B1(ram[13407]), .B2(n3475), 
        .ZN(n17648) );
  MOAI22 U26554 ( .A1(n29216), .A2(n3476), .B1(ram[13408]), .B2(n3477), 
        .ZN(n17649) );
  MOAI22 U26555 ( .A1(n28981), .A2(n3476), .B1(ram[13409]), .B2(n3477), 
        .ZN(n17650) );
  MOAI22 U26556 ( .A1(n28746), .A2(n3476), .B1(ram[13410]), .B2(n3477), 
        .ZN(n17651) );
  MOAI22 U26557 ( .A1(n28511), .A2(n3476), .B1(ram[13411]), .B2(n3477), 
        .ZN(n17652) );
  MOAI22 U26558 ( .A1(n28276), .A2(n3476), .B1(ram[13412]), .B2(n3477), 
        .ZN(n17653) );
  MOAI22 U26559 ( .A1(n28041), .A2(n3476), .B1(ram[13413]), .B2(n3477), 
        .ZN(n17654) );
  MOAI22 U26560 ( .A1(n27806), .A2(n3476), .B1(ram[13414]), .B2(n3477), 
        .ZN(n17655) );
  MOAI22 U26561 ( .A1(n27571), .A2(n3476), .B1(ram[13415]), .B2(n3477), 
        .ZN(n17656) );
  MOAI22 U26562 ( .A1(n29217), .A2(n3478), .B1(ram[13416]), .B2(n3479), 
        .ZN(n17657) );
  MOAI22 U26563 ( .A1(n28982), .A2(n3478), .B1(ram[13417]), .B2(n3479), 
        .ZN(n17658) );
  MOAI22 U26564 ( .A1(n28747), .A2(n3478), .B1(ram[13418]), .B2(n3479), 
        .ZN(n17659) );
  MOAI22 U26565 ( .A1(n28512), .A2(n3478), .B1(ram[13419]), .B2(n3479), 
        .ZN(n17660) );
  MOAI22 U26566 ( .A1(n28277), .A2(n3478), .B1(ram[13420]), .B2(n3479), 
        .ZN(n17661) );
  MOAI22 U26567 ( .A1(n28042), .A2(n3478), .B1(ram[13421]), .B2(n3479), 
        .ZN(n17662) );
  MOAI22 U26568 ( .A1(n27807), .A2(n3478), .B1(ram[13422]), .B2(n3479), 
        .ZN(n17663) );
  MOAI22 U26569 ( .A1(n27572), .A2(n3478), .B1(ram[13423]), .B2(n3479), 
        .ZN(n17664) );
  MOAI22 U26570 ( .A1(n29217), .A2(n3480), .B1(ram[13424]), .B2(n3481), 
        .ZN(n17665) );
  MOAI22 U26571 ( .A1(n28982), .A2(n3480), .B1(ram[13425]), .B2(n3481), 
        .ZN(n17666) );
  MOAI22 U26572 ( .A1(n28747), .A2(n3480), .B1(ram[13426]), .B2(n3481), 
        .ZN(n17667) );
  MOAI22 U26573 ( .A1(n28512), .A2(n3480), .B1(ram[13427]), .B2(n3481), 
        .ZN(n17668) );
  MOAI22 U26574 ( .A1(n28277), .A2(n3480), .B1(ram[13428]), .B2(n3481), 
        .ZN(n17669) );
  MOAI22 U26575 ( .A1(n28042), .A2(n3480), .B1(ram[13429]), .B2(n3481), 
        .ZN(n17670) );
  MOAI22 U26576 ( .A1(n27807), .A2(n3480), .B1(ram[13430]), .B2(n3481), 
        .ZN(n17671) );
  MOAI22 U26577 ( .A1(n27572), .A2(n3480), .B1(ram[13431]), .B2(n3481), 
        .ZN(n17672) );
  MOAI22 U26578 ( .A1(n29217), .A2(n3482), .B1(ram[13432]), .B2(n3483), 
        .ZN(n17673) );
  MOAI22 U26579 ( .A1(n28982), .A2(n3482), .B1(ram[13433]), .B2(n3483), 
        .ZN(n17674) );
  MOAI22 U26580 ( .A1(n28747), .A2(n3482), .B1(ram[13434]), .B2(n3483), 
        .ZN(n17675) );
  MOAI22 U26581 ( .A1(n28512), .A2(n3482), .B1(ram[13435]), .B2(n3483), 
        .ZN(n17676) );
  MOAI22 U26582 ( .A1(n28277), .A2(n3482), .B1(ram[13436]), .B2(n3483), 
        .ZN(n17677) );
  MOAI22 U26583 ( .A1(n28042), .A2(n3482), .B1(ram[13437]), .B2(n3483), 
        .ZN(n17678) );
  MOAI22 U26584 ( .A1(n27807), .A2(n3482), .B1(ram[13438]), .B2(n3483), 
        .ZN(n17679) );
  MOAI22 U26585 ( .A1(n27572), .A2(n3482), .B1(ram[13439]), .B2(n3483), 
        .ZN(n17680) );
  MOAI22 U26586 ( .A1(n29217), .A2(n3484), .B1(ram[13440]), .B2(n3485), 
        .ZN(n17681) );
  MOAI22 U26587 ( .A1(n28982), .A2(n3484), .B1(ram[13441]), .B2(n3485), 
        .ZN(n17682) );
  MOAI22 U26588 ( .A1(n28747), .A2(n3484), .B1(ram[13442]), .B2(n3485), 
        .ZN(n17683) );
  MOAI22 U26589 ( .A1(n28512), .A2(n3484), .B1(ram[13443]), .B2(n3485), 
        .ZN(n17684) );
  MOAI22 U26590 ( .A1(n28277), .A2(n3484), .B1(ram[13444]), .B2(n3485), 
        .ZN(n17685) );
  MOAI22 U26591 ( .A1(n28042), .A2(n3484), .B1(ram[13445]), .B2(n3485), 
        .ZN(n17686) );
  MOAI22 U26592 ( .A1(n27807), .A2(n3484), .B1(ram[13446]), .B2(n3485), 
        .ZN(n17687) );
  MOAI22 U26593 ( .A1(n27572), .A2(n3484), .B1(ram[13447]), .B2(n3485), 
        .ZN(n17688) );
  MOAI22 U26594 ( .A1(n29217), .A2(n3486), .B1(ram[13448]), .B2(n3487), 
        .ZN(n17689) );
  MOAI22 U26595 ( .A1(n28982), .A2(n3486), .B1(ram[13449]), .B2(n3487), 
        .ZN(n17690) );
  MOAI22 U26596 ( .A1(n28747), .A2(n3486), .B1(ram[13450]), .B2(n3487), 
        .ZN(n17691) );
  MOAI22 U26597 ( .A1(n28512), .A2(n3486), .B1(ram[13451]), .B2(n3487), 
        .ZN(n17692) );
  MOAI22 U26598 ( .A1(n28277), .A2(n3486), .B1(ram[13452]), .B2(n3487), 
        .ZN(n17693) );
  MOAI22 U26599 ( .A1(n28042), .A2(n3486), .B1(ram[13453]), .B2(n3487), 
        .ZN(n17694) );
  MOAI22 U26600 ( .A1(n27807), .A2(n3486), .B1(ram[13454]), .B2(n3487), 
        .ZN(n17695) );
  MOAI22 U26601 ( .A1(n27572), .A2(n3486), .B1(ram[13455]), .B2(n3487), 
        .ZN(n17696) );
  MOAI22 U26602 ( .A1(n29217), .A2(n3488), .B1(ram[13456]), .B2(n3489), 
        .ZN(n17697) );
  MOAI22 U26603 ( .A1(n28982), .A2(n3488), .B1(ram[13457]), .B2(n3489), 
        .ZN(n17698) );
  MOAI22 U26604 ( .A1(n28747), .A2(n3488), .B1(ram[13458]), .B2(n3489), 
        .ZN(n17699) );
  MOAI22 U26605 ( .A1(n28512), .A2(n3488), .B1(ram[13459]), .B2(n3489), 
        .ZN(n17700) );
  MOAI22 U26606 ( .A1(n28277), .A2(n3488), .B1(ram[13460]), .B2(n3489), 
        .ZN(n17701) );
  MOAI22 U26607 ( .A1(n28042), .A2(n3488), .B1(ram[13461]), .B2(n3489), 
        .ZN(n17702) );
  MOAI22 U26608 ( .A1(n27807), .A2(n3488), .B1(ram[13462]), .B2(n3489), 
        .ZN(n17703) );
  MOAI22 U26609 ( .A1(n27572), .A2(n3488), .B1(ram[13463]), .B2(n3489), 
        .ZN(n17704) );
  MOAI22 U26610 ( .A1(n29217), .A2(n3490), .B1(ram[13464]), .B2(n3491), 
        .ZN(n17705) );
  MOAI22 U26611 ( .A1(n28982), .A2(n3490), .B1(ram[13465]), .B2(n3491), 
        .ZN(n17706) );
  MOAI22 U26612 ( .A1(n28747), .A2(n3490), .B1(ram[13466]), .B2(n3491), 
        .ZN(n17707) );
  MOAI22 U26613 ( .A1(n28512), .A2(n3490), .B1(ram[13467]), .B2(n3491), 
        .ZN(n17708) );
  MOAI22 U26614 ( .A1(n28277), .A2(n3490), .B1(ram[13468]), .B2(n3491), 
        .ZN(n17709) );
  MOAI22 U26615 ( .A1(n28042), .A2(n3490), .B1(ram[13469]), .B2(n3491), 
        .ZN(n17710) );
  MOAI22 U26616 ( .A1(n27807), .A2(n3490), .B1(ram[13470]), .B2(n3491), 
        .ZN(n17711) );
  MOAI22 U26617 ( .A1(n27572), .A2(n3490), .B1(ram[13471]), .B2(n3491), 
        .ZN(n17712) );
  MOAI22 U26618 ( .A1(n29217), .A2(n3492), .B1(ram[13472]), .B2(n3493), 
        .ZN(n17713) );
  MOAI22 U26619 ( .A1(n28982), .A2(n3492), .B1(ram[13473]), .B2(n3493), 
        .ZN(n17714) );
  MOAI22 U26620 ( .A1(n28747), .A2(n3492), .B1(ram[13474]), .B2(n3493), 
        .ZN(n17715) );
  MOAI22 U26621 ( .A1(n28512), .A2(n3492), .B1(ram[13475]), .B2(n3493), 
        .ZN(n17716) );
  MOAI22 U26622 ( .A1(n28277), .A2(n3492), .B1(ram[13476]), .B2(n3493), 
        .ZN(n17717) );
  MOAI22 U26623 ( .A1(n28042), .A2(n3492), .B1(ram[13477]), .B2(n3493), 
        .ZN(n17718) );
  MOAI22 U26624 ( .A1(n27807), .A2(n3492), .B1(ram[13478]), .B2(n3493), 
        .ZN(n17719) );
  MOAI22 U26625 ( .A1(n27572), .A2(n3492), .B1(ram[13479]), .B2(n3493), 
        .ZN(n17720) );
  MOAI22 U26626 ( .A1(n29217), .A2(n3494), .B1(ram[13480]), .B2(n3495), 
        .ZN(n17721) );
  MOAI22 U26627 ( .A1(n28982), .A2(n3494), .B1(ram[13481]), .B2(n3495), 
        .ZN(n17722) );
  MOAI22 U26628 ( .A1(n28747), .A2(n3494), .B1(ram[13482]), .B2(n3495), 
        .ZN(n17723) );
  MOAI22 U26629 ( .A1(n28512), .A2(n3494), .B1(ram[13483]), .B2(n3495), 
        .ZN(n17724) );
  MOAI22 U26630 ( .A1(n28277), .A2(n3494), .B1(ram[13484]), .B2(n3495), 
        .ZN(n17725) );
  MOAI22 U26631 ( .A1(n28042), .A2(n3494), .B1(ram[13485]), .B2(n3495), 
        .ZN(n17726) );
  MOAI22 U26632 ( .A1(n27807), .A2(n3494), .B1(ram[13486]), .B2(n3495), 
        .ZN(n17727) );
  MOAI22 U26633 ( .A1(n27572), .A2(n3494), .B1(ram[13487]), .B2(n3495), 
        .ZN(n17728) );
  MOAI22 U26634 ( .A1(n29217), .A2(n3496), .B1(ram[13488]), .B2(n3497), 
        .ZN(n17729) );
  MOAI22 U26635 ( .A1(n28982), .A2(n3496), .B1(ram[13489]), .B2(n3497), 
        .ZN(n17730) );
  MOAI22 U26636 ( .A1(n28747), .A2(n3496), .B1(ram[13490]), .B2(n3497), 
        .ZN(n17731) );
  MOAI22 U26637 ( .A1(n28512), .A2(n3496), .B1(ram[13491]), .B2(n3497), 
        .ZN(n17732) );
  MOAI22 U26638 ( .A1(n28277), .A2(n3496), .B1(ram[13492]), .B2(n3497), 
        .ZN(n17733) );
  MOAI22 U26639 ( .A1(n28042), .A2(n3496), .B1(ram[13493]), .B2(n3497), 
        .ZN(n17734) );
  MOAI22 U26640 ( .A1(n27807), .A2(n3496), .B1(ram[13494]), .B2(n3497), 
        .ZN(n17735) );
  MOAI22 U26641 ( .A1(n27572), .A2(n3496), .B1(ram[13495]), .B2(n3497), 
        .ZN(n17736) );
  MOAI22 U26642 ( .A1(n29217), .A2(n3498), .B1(ram[13496]), .B2(n3499), 
        .ZN(n17737) );
  MOAI22 U26643 ( .A1(n28982), .A2(n3498), .B1(ram[13497]), .B2(n3499), 
        .ZN(n17738) );
  MOAI22 U26644 ( .A1(n28747), .A2(n3498), .B1(ram[13498]), .B2(n3499), 
        .ZN(n17739) );
  MOAI22 U26645 ( .A1(n28512), .A2(n3498), .B1(ram[13499]), .B2(n3499), 
        .ZN(n17740) );
  MOAI22 U26646 ( .A1(n28277), .A2(n3498), .B1(ram[13500]), .B2(n3499), 
        .ZN(n17741) );
  MOAI22 U26647 ( .A1(n28042), .A2(n3498), .B1(ram[13501]), .B2(n3499), 
        .ZN(n17742) );
  MOAI22 U26648 ( .A1(n27807), .A2(n3498), .B1(ram[13502]), .B2(n3499), 
        .ZN(n17743) );
  MOAI22 U26649 ( .A1(n27572), .A2(n3498), .B1(ram[13503]), .B2(n3499), 
        .ZN(n17744) );
  MOAI22 U26650 ( .A1(n29217), .A2(n3500), .B1(ram[13504]), .B2(n3501), 
        .ZN(n17745) );
  MOAI22 U26651 ( .A1(n28982), .A2(n3500), .B1(ram[13505]), .B2(n3501), 
        .ZN(n17746) );
  MOAI22 U26652 ( .A1(n28747), .A2(n3500), .B1(ram[13506]), .B2(n3501), 
        .ZN(n17747) );
  MOAI22 U26653 ( .A1(n28512), .A2(n3500), .B1(ram[13507]), .B2(n3501), 
        .ZN(n17748) );
  MOAI22 U26654 ( .A1(n28277), .A2(n3500), .B1(ram[13508]), .B2(n3501), 
        .ZN(n17749) );
  MOAI22 U26655 ( .A1(n28042), .A2(n3500), .B1(ram[13509]), .B2(n3501), 
        .ZN(n17750) );
  MOAI22 U26656 ( .A1(n27807), .A2(n3500), .B1(ram[13510]), .B2(n3501), 
        .ZN(n17751) );
  MOAI22 U26657 ( .A1(n27572), .A2(n3500), .B1(ram[13511]), .B2(n3501), 
        .ZN(n17752) );
  MOAI22 U26658 ( .A1(n29217), .A2(n3502), .B1(ram[13512]), .B2(n3503), 
        .ZN(n17753) );
  MOAI22 U26659 ( .A1(n28982), .A2(n3502), .B1(ram[13513]), .B2(n3503), 
        .ZN(n17754) );
  MOAI22 U26660 ( .A1(n28747), .A2(n3502), .B1(ram[13514]), .B2(n3503), 
        .ZN(n17755) );
  MOAI22 U26661 ( .A1(n28512), .A2(n3502), .B1(ram[13515]), .B2(n3503), 
        .ZN(n17756) );
  MOAI22 U26662 ( .A1(n28277), .A2(n3502), .B1(ram[13516]), .B2(n3503), 
        .ZN(n17757) );
  MOAI22 U26663 ( .A1(n28042), .A2(n3502), .B1(ram[13517]), .B2(n3503), 
        .ZN(n17758) );
  MOAI22 U26664 ( .A1(n27807), .A2(n3502), .B1(ram[13518]), .B2(n3503), 
        .ZN(n17759) );
  MOAI22 U26665 ( .A1(n27572), .A2(n3502), .B1(ram[13519]), .B2(n3503), 
        .ZN(n17760) );
  MOAI22 U26666 ( .A1(n29218), .A2(n3504), .B1(ram[13520]), .B2(n3505), 
        .ZN(n17761) );
  MOAI22 U26667 ( .A1(n28983), .A2(n3504), .B1(ram[13521]), .B2(n3505), 
        .ZN(n17762) );
  MOAI22 U26668 ( .A1(n28748), .A2(n3504), .B1(ram[13522]), .B2(n3505), 
        .ZN(n17763) );
  MOAI22 U26669 ( .A1(n28513), .A2(n3504), .B1(ram[13523]), .B2(n3505), 
        .ZN(n17764) );
  MOAI22 U26670 ( .A1(n28278), .A2(n3504), .B1(ram[13524]), .B2(n3505), 
        .ZN(n17765) );
  MOAI22 U26671 ( .A1(n28043), .A2(n3504), .B1(ram[13525]), .B2(n3505), 
        .ZN(n17766) );
  MOAI22 U26672 ( .A1(n27808), .A2(n3504), .B1(ram[13526]), .B2(n3505), 
        .ZN(n17767) );
  MOAI22 U26673 ( .A1(n27573), .A2(n3504), .B1(ram[13527]), .B2(n3505), 
        .ZN(n17768) );
  MOAI22 U26674 ( .A1(n29218), .A2(n3506), .B1(ram[13528]), .B2(n3507), 
        .ZN(n17769) );
  MOAI22 U26675 ( .A1(n28983), .A2(n3506), .B1(ram[13529]), .B2(n3507), 
        .ZN(n17770) );
  MOAI22 U26676 ( .A1(n28748), .A2(n3506), .B1(ram[13530]), .B2(n3507), 
        .ZN(n17771) );
  MOAI22 U26677 ( .A1(n28513), .A2(n3506), .B1(ram[13531]), .B2(n3507), 
        .ZN(n17772) );
  MOAI22 U26678 ( .A1(n28278), .A2(n3506), .B1(ram[13532]), .B2(n3507), 
        .ZN(n17773) );
  MOAI22 U26679 ( .A1(n28043), .A2(n3506), .B1(ram[13533]), .B2(n3507), 
        .ZN(n17774) );
  MOAI22 U26680 ( .A1(n27808), .A2(n3506), .B1(ram[13534]), .B2(n3507), 
        .ZN(n17775) );
  MOAI22 U26681 ( .A1(n27573), .A2(n3506), .B1(ram[13535]), .B2(n3507), 
        .ZN(n17776) );
  MOAI22 U26682 ( .A1(n29218), .A2(n3508), .B1(ram[13536]), .B2(n3509), 
        .ZN(n17777) );
  MOAI22 U26683 ( .A1(n28983), .A2(n3508), .B1(ram[13537]), .B2(n3509), 
        .ZN(n17778) );
  MOAI22 U26684 ( .A1(n28748), .A2(n3508), .B1(ram[13538]), .B2(n3509), 
        .ZN(n17779) );
  MOAI22 U26685 ( .A1(n28513), .A2(n3508), .B1(ram[13539]), .B2(n3509), 
        .ZN(n17780) );
  MOAI22 U26686 ( .A1(n28278), .A2(n3508), .B1(ram[13540]), .B2(n3509), 
        .ZN(n17781) );
  MOAI22 U26687 ( .A1(n28043), .A2(n3508), .B1(ram[13541]), .B2(n3509), 
        .ZN(n17782) );
  MOAI22 U26688 ( .A1(n27808), .A2(n3508), .B1(ram[13542]), .B2(n3509), 
        .ZN(n17783) );
  MOAI22 U26689 ( .A1(n27573), .A2(n3508), .B1(ram[13543]), .B2(n3509), 
        .ZN(n17784) );
  MOAI22 U26690 ( .A1(n29218), .A2(n3510), .B1(ram[13544]), .B2(n3511), 
        .ZN(n17785) );
  MOAI22 U26691 ( .A1(n28983), .A2(n3510), .B1(ram[13545]), .B2(n3511), 
        .ZN(n17786) );
  MOAI22 U26692 ( .A1(n28748), .A2(n3510), .B1(ram[13546]), .B2(n3511), 
        .ZN(n17787) );
  MOAI22 U26693 ( .A1(n28513), .A2(n3510), .B1(ram[13547]), .B2(n3511), 
        .ZN(n17788) );
  MOAI22 U26694 ( .A1(n28278), .A2(n3510), .B1(ram[13548]), .B2(n3511), 
        .ZN(n17789) );
  MOAI22 U26695 ( .A1(n28043), .A2(n3510), .B1(ram[13549]), .B2(n3511), 
        .ZN(n17790) );
  MOAI22 U26696 ( .A1(n27808), .A2(n3510), .B1(ram[13550]), .B2(n3511), 
        .ZN(n17791) );
  MOAI22 U26697 ( .A1(n27573), .A2(n3510), .B1(ram[13551]), .B2(n3511), 
        .ZN(n17792) );
  MOAI22 U26698 ( .A1(n29218), .A2(n3512), .B1(ram[13552]), .B2(n3513), 
        .ZN(n17793) );
  MOAI22 U26699 ( .A1(n28983), .A2(n3512), .B1(ram[13553]), .B2(n3513), 
        .ZN(n17794) );
  MOAI22 U26700 ( .A1(n28748), .A2(n3512), .B1(ram[13554]), .B2(n3513), 
        .ZN(n17795) );
  MOAI22 U26701 ( .A1(n28513), .A2(n3512), .B1(ram[13555]), .B2(n3513), 
        .ZN(n17796) );
  MOAI22 U26702 ( .A1(n28278), .A2(n3512), .B1(ram[13556]), .B2(n3513), 
        .ZN(n17797) );
  MOAI22 U26703 ( .A1(n28043), .A2(n3512), .B1(ram[13557]), .B2(n3513), 
        .ZN(n17798) );
  MOAI22 U26704 ( .A1(n27808), .A2(n3512), .B1(ram[13558]), .B2(n3513), 
        .ZN(n17799) );
  MOAI22 U26705 ( .A1(n27573), .A2(n3512), .B1(ram[13559]), .B2(n3513), 
        .ZN(n17800) );
  MOAI22 U26706 ( .A1(n29218), .A2(n3514), .B1(ram[13560]), .B2(n3515), 
        .ZN(n17801) );
  MOAI22 U26707 ( .A1(n28983), .A2(n3514), .B1(ram[13561]), .B2(n3515), 
        .ZN(n17802) );
  MOAI22 U26708 ( .A1(n28748), .A2(n3514), .B1(ram[13562]), .B2(n3515), 
        .ZN(n17803) );
  MOAI22 U26709 ( .A1(n28513), .A2(n3514), .B1(ram[13563]), .B2(n3515), 
        .ZN(n17804) );
  MOAI22 U26710 ( .A1(n28278), .A2(n3514), .B1(ram[13564]), .B2(n3515), 
        .ZN(n17805) );
  MOAI22 U26711 ( .A1(n28043), .A2(n3514), .B1(ram[13565]), .B2(n3515), 
        .ZN(n17806) );
  MOAI22 U26712 ( .A1(n27808), .A2(n3514), .B1(ram[13566]), .B2(n3515), 
        .ZN(n17807) );
  MOAI22 U26713 ( .A1(n27573), .A2(n3514), .B1(ram[13567]), .B2(n3515), 
        .ZN(n17808) );
  MOAI22 U26714 ( .A1(n29218), .A2(n3516), .B1(ram[13568]), .B2(n3517), 
        .ZN(n17809) );
  MOAI22 U26715 ( .A1(n28983), .A2(n3516), .B1(ram[13569]), .B2(n3517), 
        .ZN(n17810) );
  MOAI22 U26716 ( .A1(n28748), .A2(n3516), .B1(ram[13570]), .B2(n3517), 
        .ZN(n17811) );
  MOAI22 U26717 ( .A1(n28513), .A2(n3516), .B1(ram[13571]), .B2(n3517), 
        .ZN(n17812) );
  MOAI22 U26718 ( .A1(n28278), .A2(n3516), .B1(ram[13572]), .B2(n3517), 
        .ZN(n17813) );
  MOAI22 U26719 ( .A1(n28043), .A2(n3516), .B1(ram[13573]), .B2(n3517), 
        .ZN(n17814) );
  MOAI22 U26720 ( .A1(n27808), .A2(n3516), .B1(ram[13574]), .B2(n3517), 
        .ZN(n17815) );
  MOAI22 U26721 ( .A1(n27573), .A2(n3516), .B1(ram[13575]), .B2(n3517), 
        .ZN(n17816) );
  MOAI22 U26722 ( .A1(n29218), .A2(n3518), .B1(ram[13576]), .B2(n3519), 
        .ZN(n17817) );
  MOAI22 U26723 ( .A1(n28983), .A2(n3518), .B1(ram[13577]), .B2(n3519), 
        .ZN(n17818) );
  MOAI22 U26724 ( .A1(n28748), .A2(n3518), .B1(ram[13578]), .B2(n3519), 
        .ZN(n17819) );
  MOAI22 U26725 ( .A1(n28513), .A2(n3518), .B1(ram[13579]), .B2(n3519), 
        .ZN(n17820) );
  MOAI22 U26726 ( .A1(n28278), .A2(n3518), .B1(ram[13580]), .B2(n3519), 
        .ZN(n17821) );
  MOAI22 U26727 ( .A1(n28043), .A2(n3518), .B1(ram[13581]), .B2(n3519), 
        .ZN(n17822) );
  MOAI22 U26728 ( .A1(n27808), .A2(n3518), .B1(ram[13582]), .B2(n3519), 
        .ZN(n17823) );
  MOAI22 U26729 ( .A1(n27573), .A2(n3518), .B1(ram[13583]), .B2(n3519), 
        .ZN(n17824) );
  MOAI22 U26730 ( .A1(n29218), .A2(n3520), .B1(ram[13584]), .B2(n3521), 
        .ZN(n17825) );
  MOAI22 U26731 ( .A1(n28983), .A2(n3520), .B1(ram[13585]), .B2(n3521), 
        .ZN(n17826) );
  MOAI22 U26732 ( .A1(n28748), .A2(n3520), .B1(ram[13586]), .B2(n3521), 
        .ZN(n17827) );
  MOAI22 U26733 ( .A1(n28513), .A2(n3520), .B1(ram[13587]), .B2(n3521), 
        .ZN(n17828) );
  MOAI22 U26734 ( .A1(n28278), .A2(n3520), .B1(ram[13588]), .B2(n3521), 
        .ZN(n17829) );
  MOAI22 U26735 ( .A1(n28043), .A2(n3520), .B1(ram[13589]), .B2(n3521), 
        .ZN(n17830) );
  MOAI22 U26736 ( .A1(n27808), .A2(n3520), .B1(ram[13590]), .B2(n3521), 
        .ZN(n17831) );
  MOAI22 U26737 ( .A1(n27573), .A2(n3520), .B1(ram[13591]), .B2(n3521), 
        .ZN(n17832) );
  MOAI22 U26738 ( .A1(n29218), .A2(n3522), .B1(ram[13592]), .B2(n3523), 
        .ZN(n17833) );
  MOAI22 U26739 ( .A1(n28983), .A2(n3522), .B1(ram[13593]), .B2(n3523), 
        .ZN(n17834) );
  MOAI22 U26740 ( .A1(n28748), .A2(n3522), .B1(ram[13594]), .B2(n3523), 
        .ZN(n17835) );
  MOAI22 U26741 ( .A1(n28513), .A2(n3522), .B1(ram[13595]), .B2(n3523), 
        .ZN(n17836) );
  MOAI22 U26742 ( .A1(n28278), .A2(n3522), .B1(ram[13596]), .B2(n3523), 
        .ZN(n17837) );
  MOAI22 U26743 ( .A1(n28043), .A2(n3522), .B1(ram[13597]), .B2(n3523), 
        .ZN(n17838) );
  MOAI22 U26744 ( .A1(n27808), .A2(n3522), .B1(ram[13598]), .B2(n3523), 
        .ZN(n17839) );
  MOAI22 U26745 ( .A1(n27573), .A2(n3522), .B1(ram[13599]), .B2(n3523), 
        .ZN(n17840) );
  MOAI22 U26746 ( .A1(n29218), .A2(n3524), .B1(ram[13600]), .B2(n3525), 
        .ZN(n17841) );
  MOAI22 U26747 ( .A1(n28983), .A2(n3524), .B1(ram[13601]), .B2(n3525), 
        .ZN(n17842) );
  MOAI22 U26748 ( .A1(n28748), .A2(n3524), .B1(ram[13602]), .B2(n3525), 
        .ZN(n17843) );
  MOAI22 U26749 ( .A1(n28513), .A2(n3524), .B1(ram[13603]), .B2(n3525), 
        .ZN(n17844) );
  MOAI22 U26750 ( .A1(n28278), .A2(n3524), .B1(ram[13604]), .B2(n3525), 
        .ZN(n17845) );
  MOAI22 U26751 ( .A1(n28043), .A2(n3524), .B1(ram[13605]), .B2(n3525), 
        .ZN(n17846) );
  MOAI22 U26752 ( .A1(n27808), .A2(n3524), .B1(ram[13606]), .B2(n3525), 
        .ZN(n17847) );
  MOAI22 U26753 ( .A1(n27573), .A2(n3524), .B1(ram[13607]), .B2(n3525), 
        .ZN(n17848) );
  MOAI22 U26754 ( .A1(n29218), .A2(n3526), .B1(ram[13608]), .B2(n3527), 
        .ZN(n17849) );
  MOAI22 U26755 ( .A1(n28983), .A2(n3526), .B1(ram[13609]), .B2(n3527), 
        .ZN(n17850) );
  MOAI22 U26756 ( .A1(n28748), .A2(n3526), .B1(ram[13610]), .B2(n3527), 
        .ZN(n17851) );
  MOAI22 U26757 ( .A1(n28513), .A2(n3526), .B1(ram[13611]), .B2(n3527), 
        .ZN(n17852) );
  MOAI22 U26758 ( .A1(n28278), .A2(n3526), .B1(ram[13612]), .B2(n3527), 
        .ZN(n17853) );
  MOAI22 U26759 ( .A1(n28043), .A2(n3526), .B1(ram[13613]), .B2(n3527), 
        .ZN(n17854) );
  MOAI22 U26760 ( .A1(n27808), .A2(n3526), .B1(ram[13614]), .B2(n3527), 
        .ZN(n17855) );
  MOAI22 U26761 ( .A1(n27573), .A2(n3526), .B1(ram[13615]), .B2(n3527), 
        .ZN(n17856) );
  MOAI22 U26762 ( .A1(n29218), .A2(n3528), .B1(ram[13616]), .B2(n3529), 
        .ZN(n17857) );
  MOAI22 U26763 ( .A1(n28983), .A2(n3528), .B1(ram[13617]), .B2(n3529), 
        .ZN(n17858) );
  MOAI22 U26764 ( .A1(n28748), .A2(n3528), .B1(ram[13618]), .B2(n3529), 
        .ZN(n17859) );
  MOAI22 U26765 ( .A1(n28513), .A2(n3528), .B1(ram[13619]), .B2(n3529), 
        .ZN(n17860) );
  MOAI22 U26766 ( .A1(n28278), .A2(n3528), .B1(ram[13620]), .B2(n3529), 
        .ZN(n17861) );
  MOAI22 U26767 ( .A1(n28043), .A2(n3528), .B1(ram[13621]), .B2(n3529), 
        .ZN(n17862) );
  MOAI22 U26768 ( .A1(n27808), .A2(n3528), .B1(ram[13622]), .B2(n3529), 
        .ZN(n17863) );
  MOAI22 U26769 ( .A1(n27573), .A2(n3528), .B1(ram[13623]), .B2(n3529), 
        .ZN(n17864) );
  MOAI22 U26770 ( .A1(n29219), .A2(n3530), .B1(ram[13624]), .B2(n3531), 
        .ZN(n17865) );
  MOAI22 U26771 ( .A1(n28984), .A2(n3530), .B1(ram[13625]), .B2(n3531), 
        .ZN(n17866) );
  MOAI22 U26772 ( .A1(n28749), .A2(n3530), .B1(ram[13626]), .B2(n3531), 
        .ZN(n17867) );
  MOAI22 U26773 ( .A1(n28514), .A2(n3530), .B1(ram[13627]), .B2(n3531), 
        .ZN(n17868) );
  MOAI22 U26774 ( .A1(n28279), .A2(n3530), .B1(ram[13628]), .B2(n3531), 
        .ZN(n17869) );
  MOAI22 U26775 ( .A1(n28044), .A2(n3530), .B1(ram[13629]), .B2(n3531), 
        .ZN(n17870) );
  MOAI22 U26776 ( .A1(n27809), .A2(n3530), .B1(ram[13630]), .B2(n3531), 
        .ZN(n17871) );
  MOAI22 U26777 ( .A1(n27574), .A2(n3530), .B1(ram[13631]), .B2(n3531), 
        .ZN(n17872) );
  MOAI22 U26778 ( .A1(n29219), .A2(n3532), .B1(ram[13632]), .B2(n3533), 
        .ZN(n17873) );
  MOAI22 U26779 ( .A1(n28984), .A2(n3532), .B1(ram[13633]), .B2(n3533), 
        .ZN(n17874) );
  MOAI22 U26780 ( .A1(n28749), .A2(n3532), .B1(ram[13634]), .B2(n3533), 
        .ZN(n17875) );
  MOAI22 U26781 ( .A1(n28514), .A2(n3532), .B1(ram[13635]), .B2(n3533), 
        .ZN(n17876) );
  MOAI22 U26782 ( .A1(n28279), .A2(n3532), .B1(ram[13636]), .B2(n3533), 
        .ZN(n17877) );
  MOAI22 U26783 ( .A1(n28044), .A2(n3532), .B1(ram[13637]), .B2(n3533), 
        .ZN(n17878) );
  MOAI22 U26784 ( .A1(n27809), .A2(n3532), .B1(ram[13638]), .B2(n3533), 
        .ZN(n17879) );
  MOAI22 U26785 ( .A1(n27574), .A2(n3532), .B1(ram[13639]), .B2(n3533), 
        .ZN(n17880) );
  MOAI22 U26786 ( .A1(n29219), .A2(n3534), .B1(ram[13640]), .B2(n3535), 
        .ZN(n17881) );
  MOAI22 U26787 ( .A1(n28984), .A2(n3534), .B1(ram[13641]), .B2(n3535), 
        .ZN(n17882) );
  MOAI22 U26788 ( .A1(n28749), .A2(n3534), .B1(ram[13642]), .B2(n3535), 
        .ZN(n17883) );
  MOAI22 U26789 ( .A1(n28514), .A2(n3534), .B1(ram[13643]), .B2(n3535), 
        .ZN(n17884) );
  MOAI22 U26790 ( .A1(n28279), .A2(n3534), .B1(ram[13644]), .B2(n3535), 
        .ZN(n17885) );
  MOAI22 U26791 ( .A1(n28044), .A2(n3534), .B1(ram[13645]), .B2(n3535), 
        .ZN(n17886) );
  MOAI22 U26792 ( .A1(n27809), .A2(n3534), .B1(ram[13646]), .B2(n3535), 
        .ZN(n17887) );
  MOAI22 U26793 ( .A1(n27574), .A2(n3534), .B1(ram[13647]), .B2(n3535), 
        .ZN(n17888) );
  MOAI22 U26794 ( .A1(n29219), .A2(n3536), .B1(ram[13648]), .B2(n3537), 
        .ZN(n17889) );
  MOAI22 U26795 ( .A1(n28984), .A2(n3536), .B1(ram[13649]), .B2(n3537), 
        .ZN(n17890) );
  MOAI22 U26796 ( .A1(n28749), .A2(n3536), .B1(ram[13650]), .B2(n3537), 
        .ZN(n17891) );
  MOAI22 U26797 ( .A1(n28514), .A2(n3536), .B1(ram[13651]), .B2(n3537), 
        .ZN(n17892) );
  MOAI22 U26798 ( .A1(n28279), .A2(n3536), .B1(ram[13652]), .B2(n3537), 
        .ZN(n17893) );
  MOAI22 U26799 ( .A1(n28044), .A2(n3536), .B1(ram[13653]), .B2(n3537), 
        .ZN(n17894) );
  MOAI22 U26800 ( .A1(n27809), .A2(n3536), .B1(ram[13654]), .B2(n3537), 
        .ZN(n17895) );
  MOAI22 U26801 ( .A1(n27574), .A2(n3536), .B1(ram[13655]), .B2(n3537), 
        .ZN(n17896) );
  MOAI22 U26802 ( .A1(n29219), .A2(n3538), .B1(ram[13656]), .B2(n3539), 
        .ZN(n17897) );
  MOAI22 U26803 ( .A1(n28984), .A2(n3538), .B1(ram[13657]), .B2(n3539), 
        .ZN(n17898) );
  MOAI22 U26804 ( .A1(n28749), .A2(n3538), .B1(ram[13658]), .B2(n3539), 
        .ZN(n17899) );
  MOAI22 U26805 ( .A1(n28514), .A2(n3538), .B1(ram[13659]), .B2(n3539), 
        .ZN(n17900) );
  MOAI22 U26806 ( .A1(n28279), .A2(n3538), .B1(ram[13660]), .B2(n3539), 
        .ZN(n17901) );
  MOAI22 U26807 ( .A1(n28044), .A2(n3538), .B1(ram[13661]), .B2(n3539), 
        .ZN(n17902) );
  MOAI22 U26808 ( .A1(n27809), .A2(n3538), .B1(ram[13662]), .B2(n3539), 
        .ZN(n17903) );
  MOAI22 U26809 ( .A1(n27574), .A2(n3538), .B1(ram[13663]), .B2(n3539), 
        .ZN(n17904) );
  MOAI22 U26810 ( .A1(n29219), .A2(n3540), .B1(ram[13664]), .B2(n3541), 
        .ZN(n17905) );
  MOAI22 U26811 ( .A1(n28984), .A2(n3540), .B1(ram[13665]), .B2(n3541), 
        .ZN(n17906) );
  MOAI22 U26812 ( .A1(n28749), .A2(n3540), .B1(ram[13666]), .B2(n3541), 
        .ZN(n17907) );
  MOAI22 U26813 ( .A1(n28514), .A2(n3540), .B1(ram[13667]), .B2(n3541), 
        .ZN(n17908) );
  MOAI22 U26814 ( .A1(n28279), .A2(n3540), .B1(ram[13668]), .B2(n3541), 
        .ZN(n17909) );
  MOAI22 U26815 ( .A1(n28044), .A2(n3540), .B1(ram[13669]), .B2(n3541), 
        .ZN(n17910) );
  MOAI22 U26816 ( .A1(n27809), .A2(n3540), .B1(ram[13670]), .B2(n3541), 
        .ZN(n17911) );
  MOAI22 U26817 ( .A1(n27574), .A2(n3540), .B1(ram[13671]), .B2(n3541), 
        .ZN(n17912) );
  MOAI22 U26818 ( .A1(n29219), .A2(n3542), .B1(ram[13672]), .B2(n3543), 
        .ZN(n17913) );
  MOAI22 U26819 ( .A1(n28984), .A2(n3542), .B1(ram[13673]), .B2(n3543), 
        .ZN(n17914) );
  MOAI22 U26820 ( .A1(n28749), .A2(n3542), .B1(ram[13674]), .B2(n3543), 
        .ZN(n17915) );
  MOAI22 U26821 ( .A1(n28514), .A2(n3542), .B1(ram[13675]), .B2(n3543), 
        .ZN(n17916) );
  MOAI22 U26822 ( .A1(n28279), .A2(n3542), .B1(ram[13676]), .B2(n3543), 
        .ZN(n17917) );
  MOAI22 U26823 ( .A1(n28044), .A2(n3542), .B1(ram[13677]), .B2(n3543), 
        .ZN(n17918) );
  MOAI22 U26824 ( .A1(n27809), .A2(n3542), .B1(ram[13678]), .B2(n3543), 
        .ZN(n17919) );
  MOAI22 U26825 ( .A1(n27574), .A2(n3542), .B1(ram[13679]), .B2(n3543), 
        .ZN(n17920) );
  MOAI22 U26826 ( .A1(n29219), .A2(n3544), .B1(ram[13680]), .B2(n3545), 
        .ZN(n17921) );
  MOAI22 U26827 ( .A1(n28984), .A2(n3544), .B1(ram[13681]), .B2(n3545), 
        .ZN(n17922) );
  MOAI22 U26828 ( .A1(n28749), .A2(n3544), .B1(ram[13682]), .B2(n3545), 
        .ZN(n17923) );
  MOAI22 U26829 ( .A1(n28514), .A2(n3544), .B1(ram[13683]), .B2(n3545), 
        .ZN(n17924) );
  MOAI22 U26830 ( .A1(n28279), .A2(n3544), .B1(ram[13684]), .B2(n3545), 
        .ZN(n17925) );
  MOAI22 U26831 ( .A1(n28044), .A2(n3544), .B1(ram[13685]), .B2(n3545), 
        .ZN(n17926) );
  MOAI22 U26832 ( .A1(n27809), .A2(n3544), .B1(ram[13686]), .B2(n3545), 
        .ZN(n17927) );
  MOAI22 U26833 ( .A1(n27574), .A2(n3544), .B1(ram[13687]), .B2(n3545), 
        .ZN(n17928) );
  MOAI22 U26834 ( .A1(n29219), .A2(n3546), .B1(ram[13688]), .B2(n3547), 
        .ZN(n17929) );
  MOAI22 U26835 ( .A1(n28984), .A2(n3546), .B1(ram[13689]), .B2(n3547), 
        .ZN(n17930) );
  MOAI22 U26836 ( .A1(n28749), .A2(n3546), .B1(ram[13690]), .B2(n3547), 
        .ZN(n17931) );
  MOAI22 U26837 ( .A1(n28514), .A2(n3546), .B1(ram[13691]), .B2(n3547), 
        .ZN(n17932) );
  MOAI22 U26838 ( .A1(n28279), .A2(n3546), .B1(ram[13692]), .B2(n3547), 
        .ZN(n17933) );
  MOAI22 U26839 ( .A1(n28044), .A2(n3546), .B1(ram[13693]), .B2(n3547), 
        .ZN(n17934) );
  MOAI22 U26840 ( .A1(n27809), .A2(n3546), .B1(ram[13694]), .B2(n3547), 
        .ZN(n17935) );
  MOAI22 U26841 ( .A1(n27574), .A2(n3546), .B1(ram[13695]), .B2(n3547), 
        .ZN(n17936) );
  MOAI22 U26842 ( .A1(n29219), .A2(n3548), .B1(ram[13696]), .B2(n3549), 
        .ZN(n17937) );
  MOAI22 U26843 ( .A1(n28984), .A2(n3548), .B1(ram[13697]), .B2(n3549), 
        .ZN(n17938) );
  MOAI22 U26844 ( .A1(n28749), .A2(n3548), .B1(ram[13698]), .B2(n3549), 
        .ZN(n17939) );
  MOAI22 U26845 ( .A1(n28514), .A2(n3548), .B1(ram[13699]), .B2(n3549), 
        .ZN(n17940) );
  MOAI22 U26846 ( .A1(n28279), .A2(n3548), .B1(ram[13700]), .B2(n3549), 
        .ZN(n17941) );
  MOAI22 U26847 ( .A1(n28044), .A2(n3548), .B1(ram[13701]), .B2(n3549), 
        .ZN(n17942) );
  MOAI22 U26848 ( .A1(n27809), .A2(n3548), .B1(ram[13702]), .B2(n3549), 
        .ZN(n17943) );
  MOAI22 U26849 ( .A1(n27574), .A2(n3548), .B1(ram[13703]), .B2(n3549), 
        .ZN(n17944) );
  MOAI22 U26850 ( .A1(n29219), .A2(n3550), .B1(ram[13704]), .B2(n3551), 
        .ZN(n17945) );
  MOAI22 U26851 ( .A1(n28984), .A2(n3550), .B1(ram[13705]), .B2(n3551), 
        .ZN(n17946) );
  MOAI22 U26852 ( .A1(n28749), .A2(n3550), .B1(ram[13706]), .B2(n3551), 
        .ZN(n17947) );
  MOAI22 U26853 ( .A1(n28514), .A2(n3550), .B1(ram[13707]), .B2(n3551), 
        .ZN(n17948) );
  MOAI22 U26854 ( .A1(n28279), .A2(n3550), .B1(ram[13708]), .B2(n3551), 
        .ZN(n17949) );
  MOAI22 U26855 ( .A1(n28044), .A2(n3550), .B1(ram[13709]), .B2(n3551), 
        .ZN(n17950) );
  MOAI22 U26856 ( .A1(n27809), .A2(n3550), .B1(ram[13710]), .B2(n3551), 
        .ZN(n17951) );
  MOAI22 U26857 ( .A1(n27574), .A2(n3550), .B1(ram[13711]), .B2(n3551), 
        .ZN(n17952) );
  MOAI22 U26858 ( .A1(n29219), .A2(n3552), .B1(ram[13712]), .B2(n3553), 
        .ZN(n17953) );
  MOAI22 U26859 ( .A1(n28984), .A2(n3552), .B1(ram[13713]), .B2(n3553), 
        .ZN(n17954) );
  MOAI22 U26860 ( .A1(n28749), .A2(n3552), .B1(ram[13714]), .B2(n3553), 
        .ZN(n17955) );
  MOAI22 U26861 ( .A1(n28514), .A2(n3552), .B1(ram[13715]), .B2(n3553), 
        .ZN(n17956) );
  MOAI22 U26862 ( .A1(n28279), .A2(n3552), .B1(ram[13716]), .B2(n3553), 
        .ZN(n17957) );
  MOAI22 U26863 ( .A1(n28044), .A2(n3552), .B1(ram[13717]), .B2(n3553), 
        .ZN(n17958) );
  MOAI22 U26864 ( .A1(n27809), .A2(n3552), .B1(ram[13718]), .B2(n3553), 
        .ZN(n17959) );
  MOAI22 U26865 ( .A1(n27574), .A2(n3552), .B1(ram[13719]), .B2(n3553), 
        .ZN(n17960) );
  MOAI22 U26866 ( .A1(n29219), .A2(n3554), .B1(ram[13720]), .B2(n3555), 
        .ZN(n17961) );
  MOAI22 U26867 ( .A1(n28984), .A2(n3554), .B1(ram[13721]), .B2(n3555), 
        .ZN(n17962) );
  MOAI22 U26868 ( .A1(n28749), .A2(n3554), .B1(ram[13722]), .B2(n3555), 
        .ZN(n17963) );
  MOAI22 U26869 ( .A1(n28514), .A2(n3554), .B1(ram[13723]), .B2(n3555), 
        .ZN(n17964) );
  MOAI22 U26870 ( .A1(n28279), .A2(n3554), .B1(ram[13724]), .B2(n3555), 
        .ZN(n17965) );
  MOAI22 U26871 ( .A1(n28044), .A2(n3554), .B1(ram[13725]), .B2(n3555), 
        .ZN(n17966) );
  MOAI22 U26872 ( .A1(n27809), .A2(n3554), .B1(ram[13726]), .B2(n3555), 
        .ZN(n17967) );
  MOAI22 U26873 ( .A1(n27574), .A2(n3554), .B1(ram[13727]), .B2(n3555), 
        .ZN(n17968) );
  MOAI22 U26874 ( .A1(n29220), .A2(n3556), .B1(ram[13728]), .B2(n3557), 
        .ZN(n17969) );
  MOAI22 U26875 ( .A1(n28985), .A2(n3556), .B1(ram[13729]), .B2(n3557), 
        .ZN(n17970) );
  MOAI22 U26876 ( .A1(n28750), .A2(n3556), .B1(ram[13730]), .B2(n3557), 
        .ZN(n17971) );
  MOAI22 U26877 ( .A1(n28515), .A2(n3556), .B1(ram[13731]), .B2(n3557), 
        .ZN(n17972) );
  MOAI22 U26878 ( .A1(n28280), .A2(n3556), .B1(ram[13732]), .B2(n3557), 
        .ZN(n17973) );
  MOAI22 U26879 ( .A1(n28045), .A2(n3556), .B1(ram[13733]), .B2(n3557), 
        .ZN(n17974) );
  MOAI22 U26880 ( .A1(n27810), .A2(n3556), .B1(ram[13734]), .B2(n3557), 
        .ZN(n17975) );
  MOAI22 U26881 ( .A1(n27575), .A2(n3556), .B1(ram[13735]), .B2(n3557), 
        .ZN(n17976) );
  MOAI22 U26882 ( .A1(n29220), .A2(n3558), .B1(ram[13736]), .B2(n3559), 
        .ZN(n17977) );
  MOAI22 U26883 ( .A1(n28985), .A2(n3558), .B1(ram[13737]), .B2(n3559), 
        .ZN(n17978) );
  MOAI22 U26884 ( .A1(n28750), .A2(n3558), .B1(ram[13738]), .B2(n3559), 
        .ZN(n17979) );
  MOAI22 U26885 ( .A1(n28515), .A2(n3558), .B1(ram[13739]), .B2(n3559), 
        .ZN(n17980) );
  MOAI22 U26886 ( .A1(n28280), .A2(n3558), .B1(ram[13740]), .B2(n3559), 
        .ZN(n17981) );
  MOAI22 U26887 ( .A1(n28045), .A2(n3558), .B1(ram[13741]), .B2(n3559), 
        .ZN(n17982) );
  MOAI22 U26888 ( .A1(n27810), .A2(n3558), .B1(ram[13742]), .B2(n3559), 
        .ZN(n17983) );
  MOAI22 U26889 ( .A1(n27575), .A2(n3558), .B1(ram[13743]), .B2(n3559), 
        .ZN(n17984) );
  MOAI22 U26890 ( .A1(n29220), .A2(n3560), .B1(ram[13744]), .B2(n3561), 
        .ZN(n17985) );
  MOAI22 U26891 ( .A1(n28985), .A2(n3560), .B1(ram[13745]), .B2(n3561), 
        .ZN(n17986) );
  MOAI22 U26892 ( .A1(n28750), .A2(n3560), .B1(ram[13746]), .B2(n3561), 
        .ZN(n17987) );
  MOAI22 U26893 ( .A1(n28515), .A2(n3560), .B1(ram[13747]), .B2(n3561), 
        .ZN(n17988) );
  MOAI22 U26894 ( .A1(n28280), .A2(n3560), .B1(ram[13748]), .B2(n3561), 
        .ZN(n17989) );
  MOAI22 U26895 ( .A1(n28045), .A2(n3560), .B1(ram[13749]), .B2(n3561), 
        .ZN(n17990) );
  MOAI22 U26896 ( .A1(n27810), .A2(n3560), .B1(ram[13750]), .B2(n3561), 
        .ZN(n17991) );
  MOAI22 U26897 ( .A1(n27575), .A2(n3560), .B1(ram[13751]), .B2(n3561), 
        .ZN(n17992) );
  MOAI22 U26898 ( .A1(n29220), .A2(n3562), .B1(ram[13752]), .B2(n3563), 
        .ZN(n17993) );
  MOAI22 U26899 ( .A1(n28985), .A2(n3562), .B1(ram[13753]), .B2(n3563), 
        .ZN(n17994) );
  MOAI22 U26900 ( .A1(n28750), .A2(n3562), .B1(ram[13754]), .B2(n3563), 
        .ZN(n17995) );
  MOAI22 U26901 ( .A1(n28515), .A2(n3562), .B1(ram[13755]), .B2(n3563), 
        .ZN(n17996) );
  MOAI22 U26902 ( .A1(n28280), .A2(n3562), .B1(ram[13756]), .B2(n3563), 
        .ZN(n17997) );
  MOAI22 U26903 ( .A1(n28045), .A2(n3562), .B1(ram[13757]), .B2(n3563), 
        .ZN(n17998) );
  MOAI22 U26904 ( .A1(n27810), .A2(n3562), .B1(ram[13758]), .B2(n3563), 
        .ZN(n17999) );
  MOAI22 U26905 ( .A1(n27575), .A2(n3562), .B1(ram[13759]), .B2(n3563), 
        .ZN(n18000) );
  MOAI22 U26906 ( .A1(n29220), .A2(n3564), .B1(ram[13760]), .B2(n3565), 
        .ZN(n18001) );
  MOAI22 U26907 ( .A1(n28985), .A2(n3564), .B1(ram[13761]), .B2(n3565), 
        .ZN(n18002) );
  MOAI22 U26908 ( .A1(n28750), .A2(n3564), .B1(ram[13762]), .B2(n3565), 
        .ZN(n18003) );
  MOAI22 U26909 ( .A1(n28515), .A2(n3564), .B1(ram[13763]), .B2(n3565), 
        .ZN(n18004) );
  MOAI22 U26910 ( .A1(n28280), .A2(n3564), .B1(ram[13764]), .B2(n3565), 
        .ZN(n18005) );
  MOAI22 U26911 ( .A1(n28045), .A2(n3564), .B1(ram[13765]), .B2(n3565), 
        .ZN(n18006) );
  MOAI22 U26912 ( .A1(n27810), .A2(n3564), .B1(ram[13766]), .B2(n3565), 
        .ZN(n18007) );
  MOAI22 U26913 ( .A1(n27575), .A2(n3564), .B1(ram[13767]), .B2(n3565), 
        .ZN(n18008) );
  MOAI22 U26914 ( .A1(n29220), .A2(n3566), .B1(ram[13768]), .B2(n3567), 
        .ZN(n18009) );
  MOAI22 U26915 ( .A1(n28985), .A2(n3566), .B1(ram[13769]), .B2(n3567), 
        .ZN(n18010) );
  MOAI22 U26916 ( .A1(n28750), .A2(n3566), .B1(ram[13770]), .B2(n3567), 
        .ZN(n18011) );
  MOAI22 U26917 ( .A1(n28515), .A2(n3566), .B1(ram[13771]), .B2(n3567), 
        .ZN(n18012) );
  MOAI22 U26918 ( .A1(n28280), .A2(n3566), .B1(ram[13772]), .B2(n3567), 
        .ZN(n18013) );
  MOAI22 U26919 ( .A1(n28045), .A2(n3566), .B1(ram[13773]), .B2(n3567), 
        .ZN(n18014) );
  MOAI22 U26920 ( .A1(n27810), .A2(n3566), .B1(ram[13774]), .B2(n3567), 
        .ZN(n18015) );
  MOAI22 U26921 ( .A1(n27575), .A2(n3566), .B1(ram[13775]), .B2(n3567), 
        .ZN(n18016) );
  MOAI22 U26922 ( .A1(n29220), .A2(n3568), .B1(ram[13776]), .B2(n3569), 
        .ZN(n18017) );
  MOAI22 U26923 ( .A1(n28985), .A2(n3568), .B1(ram[13777]), .B2(n3569), 
        .ZN(n18018) );
  MOAI22 U26924 ( .A1(n28750), .A2(n3568), .B1(ram[13778]), .B2(n3569), 
        .ZN(n18019) );
  MOAI22 U26925 ( .A1(n28515), .A2(n3568), .B1(ram[13779]), .B2(n3569), 
        .ZN(n18020) );
  MOAI22 U26926 ( .A1(n28280), .A2(n3568), .B1(ram[13780]), .B2(n3569), 
        .ZN(n18021) );
  MOAI22 U26927 ( .A1(n28045), .A2(n3568), .B1(ram[13781]), .B2(n3569), 
        .ZN(n18022) );
  MOAI22 U26928 ( .A1(n27810), .A2(n3568), .B1(ram[13782]), .B2(n3569), 
        .ZN(n18023) );
  MOAI22 U26929 ( .A1(n27575), .A2(n3568), .B1(ram[13783]), .B2(n3569), 
        .ZN(n18024) );
  MOAI22 U26930 ( .A1(n29220), .A2(n3570), .B1(ram[13784]), .B2(n3571), 
        .ZN(n18025) );
  MOAI22 U26931 ( .A1(n28985), .A2(n3570), .B1(ram[13785]), .B2(n3571), 
        .ZN(n18026) );
  MOAI22 U26932 ( .A1(n28750), .A2(n3570), .B1(ram[13786]), .B2(n3571), 
        .ZN(n18027) );
  MOAI22 U26933 ( .A1(n28515), .A2(n3570), .B1(ram[13787]), .B2(n3571), 
        .ZN(n18028) );
  MOAI22 U26934 ( .A1(n28280), .A2(n3570), .B1(ram[13788]), .B2(n3571), 
        .ZN(n18029) );
  MOAI22 U26935 ( .A1(n28045), .A2(n3570), .B1(ram[13789]), .B2(n3571), 
        .ZN(n18030) );
  MOAI22 U26936 ( .A1(n27810), .A2(n3570), .B1(ram[13790]), .B2(n3571), 
        .ZN(n18031) );
  MOAI22 U26937 ( .A1(n27575), .A2(n3570), .B1(ram[13791]), .B2(n3571), 
        .ZN(n18032) );
  MOAI22 U26938 ( .A1(n29220), .A2(n3572), .B1(ram[13792]), .B2(n3573), 
        .ZN(n18033) );
  MOAI22 U26939 ( .A1(n28985), .A2(n3572), .B1(ram[13793]), .B2(n3573), 
        .ZN(n18034) );
  MOAI22 U26940 ( .A1(n28750), .A2(n3572), .B1(ram[13794]), .B2(n3573), 
        .ZN(n18035) );
  MOAI22 U26941 ( .A1(n28515), .A2(n3572), .B1(ram[13795]), .B2(n3573), 
        .ZN(n18036) );
  MOAI22 U26942 ( .A1(n28280), .A2(n3572), .B1(ram[13796]), .B2(n3573), 
        .ZN(n18037) );
  MOAI22 U26943 ( .A1(n28045), .A2(n3572), .B1(ram[13797]), .B2(n3573), 
        .ZN(n18038) );
  MOAI22 U26944 ( .A1(n27810), .A2(n3572), .B1(ram[13798]), .B2(n3573), 
        .ZN(n18039) );
  MOAI22 U26945 ( .A1(n27575), .A2(n3572), .B1(ram[13799]), .B2(n3573), 
        .ZN(n18040) );
  MOAI22 U26946 ( .A1(n29220), .A2(n3574), .B1(ram[13800]), .B2(n3575), 
        .ZN(n18041) );
  MOAI22 U26947 ( .A1(n28985), .A2(n3574), .B1(ram[13801]), .B2(n3575), 
        .ZN(n18042) );
  MOAI22 U26948 ( .A1(n28750), .A2(n3574), .B1(ram[13802]), .B2(n3575), 
        .ZN(n18043) );
  MOAI22 U26949 ( .A1(n28515), .A2(n3574), .B1(ram[13803]), .B2(n3575), 
        .ZN(n18044) );
  MOAI22 U26950 ( .A1(n28280), .A2(n3574), .B1(ram[13804]), .B2(n3575), 
        .ZN(n18045) );
  MOAI22 U26951 ( .A1(n28045), .A2(n3574), .B1(ram[13805]), .B2(n3575), 
        .ZN(n18046) );
  MOAI22 U26952 ( .A1(n27810), .A2(n3574), .B1(ram[13806]), .B2(n3575), 
        .ZN(n18047) );
  MOAI22 U26953 ( .A1(n27575), .A2(n3574), .B1(ram[13807]), .B2(n3575), 
        .ZN(n18048) );
  MOAI22 U26954 ( .A1(n29220), .A2(n3576), .B1(ram[13808]), .B2(n3577), 
        .ZN(n18049) );
  MOAI22 U26955 ( .A1(n28985), .A2(n3576), .B1(ram[13809]), .B2(n3577), 
        .ZN(n18050) );
  MOAI22 U26956 ( .A1(n28750), .A2(n3576), .B1(ram[13810]), .B2(n3577), 
        .ZN(n18051) );
  MOAI22 U26957 ( .A1(n28515), .A2(n3576), .B1(ram[13811]), .B2(n3577), 
        .ZN(n18052) );
  MOAI22 U26958 ( .A1(n28280), .A2(n3576), .B1(ram[13812]), .B2(n3577), 
        .ZN(n18053) );
  MOAI22 U26959 ( .A1(n28045), .A2(n3576), .B1(ram[13813]), .B2(n3577), 
        .ZN(n18054) );
  MOAI22 U26960 ( .A1(n27810), .A2(n3576), .B1(ram[13814]), .B2(n3577), 
        .ZN(n18055) );
  MOAI22 U26961 ( .A1(n27575), .A2(n3576), .B1(ram[13815]), .B2(n3577), 
        .ZN(n18056) );
  MOAI22 U26962 ( .A1(n29220), .A2(n3578), .B1(ram[13816]), .B2(n3579), 
        .ZN(n18057) );
  MOAI22 U26963 ( .A1(n28985), .A2(n3578), .B1(ram[13817]), .B2(n3579), 
        .ZN(n18058) );
  MOAI22 U26964 ( .A1(n28750), .A2(n3578), .B1(ram[13818]), .B2(n3579), 
        .ZN(n18059) );
  MOAI22 U26965 ( .A1(n28515), .A2(n3578), .B1(ram[13819]), .B2(n3579), 
        .ZN(n18060) );
  MOAI22 U26966 ( .A1(n28280), .A2(n3578), .B1(ram[13820]), .B2(n3579), 
        .ZN(n18061) );
  MOAI22 U26967 ( .A1(n28045), .A2(n3578), .B1(ram[13821]), .B2(n3579), 
        .ZN(n18062) );
  MOAI22 U26968 ( .A1(n27810), .A2(n3578), .B1(ram[13822]), .B2(n3579), 
        .ZN(n18063) );
  MOAI22 U26969 ( .A1(n27575), .A2(n3578), .B1(ram[13823]), .B2(n3579), 
        .ZN(n18064) );
  MOAI22 U26970 ( .A1(n29220), .A2(n3580), .B1(ram[13824]), .B2(n3581), 
        .ZN(n18065) );
  MOAI22 U26971 ( .A1(n28985), .A2(n3580), .B1(ram[13825]), .B2(n3581), 
        .ZN(n18066) );
  MOAI22 U26972 ( .A1(n28750), .A2(n3580), .B1(ram[13826]), .B2(n3581), 
        .ZN(n18067) );
  MOAI22 U26973 ( .A1(n28515), .A2(n3580), .B1(ram[13827]), .B2(n3581), 
        .ZN(n18068) );
  MOAI22 U26974 ( .A1(n28280), .A2(n3580), .B1(ram[13828]), .B2(n3581), 
        .ZN(n18069) );
  MOAI22 U26975 ( .A1(n28045), .A2(n3580), .B1(ram[13829]), .B2(n3581), 
        .ZN(n18070) );
  MOAI22 U26976 ( .A1(n27810), .A2(n3580), .B1(ram[13830]), .B2(n3581), 
        .ZN(n18071) );
  MOAI22 U26977 ( .A1(n27575), .A2(n3580), .B1(ram[13831]), .B2(n3581), 
        .ZN(n18072) );
  MOAI22 U26978 ( .A1(n29221), .A2(n3583), .B1(ram[13832]), .B2(n3584), 
        .ZN(n18073) );
  MOAI22 U26979 ( .A1(n28986), .A2(n3583), .B1(ram[13833]), .B2(n3584), 
        .ZN(n18074) );
  MOAI22 U26980 ( .A1(n28751), .A2(n3583), .B1(ram[13834]), .B2(n3584), 
        .ZN(n18075) );
  MOAI22 U26981 ( .A1(n28516), .A2(n3583), .B1(ram[13835]), .B2(n3584), 
        .ZN(n18076) );
  MOAI22 U26982 ( .A1(n28281), .A2(n3583), .B1(ram[13836]), .B2(n3584), 
        .ZN(n18077) );
  MOAI22 U26983 ( .A1(n28046), .A2(n3583), .B1(ram[13837]), .B2(n3584), 
        .ZN(n18078) );
  MOAI22 U26984 ( .A1(n27811), .A2(n3583), .B1(ram[13838]), .B2(n3584), 
        .ZN(n18079) );
  MOAI22 U26985 ( .A1(n27576), .A2(n3583), .B1(ram[13839]), .B2(n3584), 
        .ZN(n18080) );
  MOAI22 U26986 ( .A1(n29221), .A2(n3585), .B1(ram[13840]), .B2(n3586), 
        .ZN(n18081) );
  MOAI22 U26987 ( .A1(n28986), .A2(n3585), .B1(ram[13841]), .B2(n3586), 
        .ZN(n18082) );
  MOAI22 U26988 ( .A1(n28751), .A2(n3585), .B1(ram[13842]), .B2(n3586), 
        .ZN(n18083) );
  MOAI22 U26989 ( .A1(n28516), .A2(n3585), .B1(ram[13843]), .B2(n3586), 
        .ZN(n18084) );
  MOAI22 U26990 ( .A1(n28281), .A2(n3585), .B1(ram[13844]), .B2(n3586), 
        .ZN(n18085) );
  MOAI22 U26991 ( .A1(n28046), .A2(n3585), .B1(ram[13845]), .B2(n3586), 
        .ZN(n18086) );
  MOAI22 U26992 ( .A1(n27811), .A2(n3585), .B1(ram[13846]), .B2(n3586), 
        .ZN(n18087) );
  MOAI22 U26993 ( .A1(n27576), .A2(n3585), .B1(ram[13847]), .B2(n3586), 
        .ZN(n18088) );
  MOAI22 U26994 ( .A1(n29221), .A2(n3587), .B1(ram[13848]), .B2(n3588), 
        .ZN(n18089) );
  MOAI22 U26995 ( .A1(n28986), .A2(n3587), .B1(ram[13849]), .B2(n3588), 
        .ZN(n18090) );
  MOAI22 U26996 ( .A1(n28751), .A2(n3587), .B1(ram[13850]), .B2(n3588), 
        .ZN(n18091) );
  MOAI22 U26997 ( .A1(n28516), .A2(n3587), .B1(ram[13851]), .B2(n3588), 
        .ZN(n18092) );
  MOAI22 U26998 ( .A1(n28281), .A2(n3587), .B1(ram[13852]), .B2(n3588), 
        .ZN(n18093) );
  MOAI22 U26999 ( .A1(n28046), .A2(n3587), .B1(ram[13853]), .B2(n3588), 
        .ZN(n18094) );
  MOAI22 U27000 ( .A1(n27811), .A2(n3587), .B1(ram[13854]), .B2(n3588), 
        .ZN(n18095) );
  MOAI22 U27001 ( .A1(n27576), .A2(n3587), .B1(ram[13855]), .B2(n3588), 
        .ZN(n18096) );
  MOAI22 U27002 ( .A1(n29221), .A2(n3589), .B1(ram[13856]), .B2(n3590), 
        .ZN(n18097) );
  MOAI22 U27003 ( .A1(n28986), .A2(n3589), .B1(ram[13857]), .B2(n3590), 
        .ZN(n18098) );
  MOAI22 U27004 ( .A1(n28751), .A2(n3589), .B1(ram[13858]), .B2(n3590), 
        .ZN(n18099) );
  MOAI22 U27005 ( .A1(n28516), .A2(n3589), .B1(ram[13859]), .B2(n3590), 
        .ZN(n18100) );
  MOAI22 U27006 ( .A1(n28281), .A2(n3589), .B1(ram[13860]), .B2(n3590), 
        .ZN(n18101) );
  MOAI22 U27007 ( .A1(n28046), .A2(n3589), .B1(ram[13861]), .B2(n3590), 
        .ZN(n18102) );
  MOAI22 U27008 ( .A1(n27811), .A2(n3589), .B1(ram[13862]), .B2(n3590), 
        .ZN(n18103) );
  MOAI22 U27009 ( .A1(n27576), .A2(n3589), .B1(ram[13863]), .B2(n3590), 
        .ZN(n18104) );
  MOAI22 U27010 ( .A1(n29221), .A2(n3591), .B1(ram[13864]), .B2(n3592), 
        .ZN(n18105) );
  MOAI22 U27011 ( .A1(n28986), .A2(n3591), .B1(ram[13865]), .B2(n3592), 
        .ZN(n18106) );
  MOAI22 U27012 ( .A1(n28751), .A2(n3591), .B1(ram[13866]), .B2(n3592), 
        .ZN(n18107) );
  MOAI22 U27013 ( .A1(n28516), .A2(n3591), .B1(ram[13867]), .B2(n3592), 
        .ZN(n18108) );
  MOAI22 U27014 ( .A1(n28281), .A2(n3591), .B1(ram[13868]), .B2(n3592), 
        .ZN(n18109) );
  MOAI22 U27015 ( .A1(n28046), .A2(n3591), .B1(ram[13869]), .B2(n3592), 
        .ZN(n18110) );
  MOAI22 U27016 ( .A1(n27811), .A2(n3591), .B1(ram[13870]), .B2(n3592), 
        .ZN(n18111) );
  MOAI22 U27017 ( .A1(n27576), .A2(n3591), .B1(ram[13871]), .B2(n3592), 
        .ZN(n18112) );
  MOAI22 U27018 ( .A1(n29221), .A2(n3593), .B1(ram[13872]), .B2(n3594), 
        .ZN(n18113) );
  MOAI22 U27019 ( .A1(n28986), .A2(n3593), .B1(ram[13873]), .B2(n3594), 
        .ZN(n18114) );
  MOAI22 U27020 ( .A1(n28751), .A2(n3593), .B1(ram[13874]), .B2(n3594), 
        .ZN(n18115) );
  MOAI22 U27021 ( .A1(n28516), .A2(n3593), .B1(ram[13875]), .B2(n3594), 
        .ZN(n18116) );
  MOAI22 U27022 ( .A1(n28281), .A2(n3593), .B1(ram[13876]), .B2(n3594), 
        .ZN(n18117) );
  MOAI22 U27023 ( .A1(n28046), .A2(n3593), .B1(ram[13877]), .B2(n3594), 
        .ZN(n18118) );
  MOAI22 U27024 ( .A1(n27811), .A2(n3593), .B1(ram[13878]), .B2(n3594), 
        .ZN(n18119) );
  MOAI22 U27025 ( .A1(n27576), .A2(n3593), .B1(ram[13879]), .B2(n3594), 
        .ZN(n18120) );
  MOAI22 U27026 ( .A1(n29221), .A2(n3595), .B1(ram[13880]), .B2(n3596), 
        .ZN(n18121) );
  MOAI22 U27027 ( .A1(n28986), .A2(n3595), .B1(ram[13881]), .B2(n3596), 
        .ZN(n18122) );
  MOAI22 U27028 ( .A1(n28751), .A2(n3595), .B1(ram[13882]), .B2(n3596), 
        .ZN(n18123) );
  MOAI22 U27029 ( .A1(n28516), .A2(n3595), .B1(ram[13883]), .B2(n3596), 
        .ZN(n18124) );
  MOAI22 U27030 ( .A1(n28281), .A2(n3595), .B1(ram[13884]), .B2(n3596), 
        .ZN(n18125) );
  MOAI22 U27031 ( .A1(n28046), .A2(n3595), .B1(ram[13885]), .B2(n3596), 
        .ZN(n18126) );
  MOAI22 U27032 ( .A1(n27811), .A2(n3595), .B1(ram[13886]), .B2(n3596), 
        .ZN(n18127) );
  MOAI22 U27033 ( .A1(n27576), .A2(n3595), .B1(ram[13887]), .B2(n3596), 
        .ZN(n18128) );
  MOAI22 U27034 ( .A1(n29221), .A2(n3597), .B1(ram[13888]), .B2(n3598), 
        .ZN(n18129) );
  MOAI22 U27035 ( .A1(n28986), .A2(n3597), .B1(ram[13889]), .B2(n3598), 
        .ZN(n18130) );
  MOAI22 U27036 ( .A1(n28751), .A2(n3597), .B1(ram[13890]), .B2(n3598), 
        .ZN(n18131) );
  MOAI22 U27037 ( .A1(n28516), .A2(n3597), .B1(ram[13891]), .B2(n3598), 
        .ZN(n18132) );
  MOAI22 U27038 ( .A1(n28281), .A2(n3597), .B1(ram[13892]), .B2(n3598), 
        .ZN(n18133) );
  MOAI22 U27039 ( .A1(n28046), .A2(n3597), .B1(ram[13893]), .B2(n3598), 
        .ZN(n18134) );
  MOAI22 U27040 ( .A1(n27811), .A2(n3597), .B1(ram[13894]), .B2(n3598), 
        .ZN(n18135) );
  MOAI22 U27041 ( .A1(n27576), .A2(n3597), .B1(ram[13895]), .B2(n3598), 
        .ZN(n18136) );
  MOAI22 U27042 ( .A1(n29221), .A2(n3599), .B1(ram[13896]), .B2(n3600), 
        .ZN(n18137) );
  MOAI22 U27043 ( .A1(n28986), .A2(n3599), .B1(ram[13897]), .B2(n3600), 
        .ZN(n18138) );
  MOAI22 U27044 ( .A1(n28751), .A2(n3599), .B1(ram[13898]), .B2(n3600), 
        .ZN(n18139) );
  MOAI22 U27045 ( .A1(n28516), .A2(n3599), .B1(ram[13899]), .B2(n3600), 
        .ZN(n18140) );
  MOAI22 U27046 ( .A1(n28281), .A2(n3599), .B1(ram[13900]), .B2(n3600), 
        .ZN(n18141) );
  MOAI22 U27047 ( .A1(n28046), .A2(n3599), .B1(ram[13901]), .B2(n3600), 
        .ZN(n18142) );
  MOAI22 U27048 ( .A1(n27811), .A2(n3599), .B1(ram[13902]), .B2(n3600), 
        .ZN(n18143) );
  MOAI22 U27049 ( .A1(n27576), .A2(n3599), .B1(ram[13903]), .B2(n3600), 
        .ZN(n18144) );
  MOAI22 U27050 ( .A1(n29221), .A2(n3601), .B1(ram[13904]), .B2(n3602), 
        .ZN(n18145) );
  MOAI22 U27051 ( .A1(n28986), .A2(n3601), .B1(ram[13905]), .B2(n3602), 
        .ZN(n18146) );
  MOAI22 U27052 ( .A1(n28751), .A2(n3601), .B1(ram[13906]), .B2(n3602), 
        .ZN(n18147) );
  MOAI22 U27053 ( .A1(n28516), .A2(n3601), .B1(ram[13907]), .B2(n3602), 
        .ZN(n18148) );
  MOAI22 U27054 ( .A1(n28281), .A2(n3601), .B1(ram[13908]), .B2(n3602), 
        .ZN(n18149) );
  MOAI22 U27055 ( .A1(n28046), .A2(n3601), .B1(ram[13909]), .B2(n3602), 
        .ZN(n18150) );
  MOAI22 U27056 ( .A1(n27811), .A2(n3601), .B1(ram[13910]), .B2(n3602), 
        .ZN(n18151) );
  MOAI22 U27057 ( .A1(n27576), .A2(n3601), .B1(ram[13911]), .B2(n3602), 
        .ZN(n18152) );
  MOAI22 U27058 ( .A1(n29221), .A2(n3603), .B1(ram[13912]), .B2(n3604), 
        .ZN(n18153) );
  MOAI22 U27059 ( .A1(n28986), .A2(n3603), .B1(ram[13913]), .B2(n3604), 
        .ZN(n18154) );
  MOAI22 U27060 ( .A1(n28751), .A2(n3603), .B1(ram[13914]), .B2(n3604), 
        .ZN(n18155) );
  MOAI22 U27061 ( .A1(n28516), .A2(n3603), .B1(ram[13915]), .B2(n3604), 
        .ZN(n18156) );
  MOAI22 U27062 ( .A1(n28281), .A2(n3603), .B1(ram[13916]), .B2(n3604), 
        .ZN(n18157) );
  MOAI22 U27063 ( .A1(n28046), .A2(n3603), .B1(ram[13917]), .B2(n3604), 
        .ZN(n18158) );
  MOAI22 U27064 ( .A1(n27811), .A2(n3603), .B1(ram[13918]), .B2(n3604), 
        .ZN(n18159) );
  MOAI22 U27065 ( .A1(n27576), .A2(n3603), .B1(ram[13919]), .B2(n3604), 
        .ZN(n18160) );
  MOAI22 U27066 ( .A1(n29221), .A2(n3605), .B1(ram[13920]), .B2(n3606), 
        .ZN(n18161) );
  MOAI22 U27067 ( .A1(n28986), .A2(n3605), .B1(ram[13921]), .B2(n3606), 
        .ZN(n18162) );
  MOAI22 U27068 ( .A1(n28751), .A2(n3605), .B1(ram[13922]), .B2(n3606), 
        .ZN(n18163) );
  MOAI22 U27069 ( .A1(n28516), .A2(n3605), .B1(ram[13923]), .B2(n3606), 
        .ZN(n18164) );
  MOAI22 U27070 ( .A1(n28281), .A2(n3605), .B1(ram[13924]), .B2(n3606), 
        .ZN(n18165) );
  MOAI22 U27071 ( .A1(n28046), .A2(n3605), .B1(ram[13925]), .B2(n3606), 
        .ZN(n18166) );
  MOAI22 U27072 ( .A1(n27811), .A2(n3605), .B1(ram[13926]), .B2(n3606), 
        .ZN(n18167) );
  MOAI22 U27073 ( .A1(n27576), .A2(n3605), .B1(ram[13927]), .B2(n3606), 
        .ZN(n18168) );
  MOAI22 U27074 ( .A1(n29221), .A2(n3607), .B1(ram[13928]), .B2(n3608), 
        .ZN(n18169) );
  MOAI22 U27075 ( .A1(n28986), .A2(n3607), .B1(ram[13929]), .B2(n3608), 
        .ZN(n18170) );
  MOAI22 U27076 ( .A1(n28751), .A2(n3607), .B1(ram[13930]), .B2(n3608), 
        .ZN(n18171) );
  MOAI22 U27077 ( .A1(n28516), .A2(n3607), .B1(ram[13931]), .B2(n3608), 
        .ZN(n18172) );
  MOAI22 U27078 ( .A1(n28281), .A2(n3607), .B1(ram[13932]), .B2(n3608), 
        .ZN(n18173) );
  MOAI22 U27079 ( .A1(n28046), .A2(n3607), .B1(ram[13933]), .B2(n3608), 
        .ZN(n18174) );
  MOAI22 U27080 ( .A1(n27811), .A2(n3607), .B1(ram[13934]), .B2(n3608), 
        .ZN(n18175) );
  MOAI22 U27081 ( .A1(n27576), .A2(n3607), .B1(ram[13935]), .B2(n3608), 
        .ZN(n18176) );
  MOAI22 U27082 ( .A1(n29222), .A2(n3609), .B1(ram[13936]), .B2(n3610), 
        .ZN(n18177) );
  MOAI22 U27083 ( .A1(n28987), .A2(n3609), .B1(ram[13937]), .B2(n3610), 
        .ZN(n18178) );
  MOAI22 U27084 ( .A1(n28752), .A2(n3609), .B1(ram[13938]), .B2(n3610), 
        .ZN(n18179) );
  MOAI22 U27085 ( .A1(n28517), .A2(n3609), .B1(ram[13939]), .B2(n3610), 
        .ZN(n18180) );
  MOAI22 U27086 ( .A1(n28282), .A2(n3609), .B1(ram[13940]), .B2(n3610), 
        .ZN(n18181) );
  MOAI22 U27087 ( .A1(n28047), .A2(n3609), .B1(ram[13941]), .B2(n3610), 
        .ZN(n18182) );
  MOAI22 U27088 ( .A1(n27812), .A2(n3609), .B1(ram[13942]), .B2(n3610), 
        .ZN(n18183) );
  MOAI22 U27089 ( .A1(n27577), .A2(n3609), .B1(ram[13943]), .B2(n3610), 
        .ZN(n18184) );
  MOAI22 U27090 ( .A1(n29222), .A2(n3611), .B1(ram[13944]), .B2(n3612), 
        .ZN(n18185) );
  MOAI22 U27091 ( .A1(n28987), .A2(n3611), .B1(ram[13945]), .B2(n3612), 
        .ZN(n18186) );
  MOAI22 U27092 ( .A1(n28752), .A2(n3611), .B1(ram[13946]), .B2(n3612), 
        .ZN(n18187) );
  MOAI22 U27093 ( .A1(n28517), .A2(n3611), .B1(ram[13947]), .B2(n3612), 
        .ZN(n18188) );
  MOAI22 U27094 ( .A1(n28282), .A2(n3611), .B1(ram[13948]), .B2(n3612), 
        .ZN(n18189) );
  MOAI22 U27095 ( .A1(n28047), .A2(n3611), .B1(ram[13949]), .B2(n3612), 
        .ZN(n18190) );
  MOAI22 U27096 ( .A1(n27812), .A2(n3611), .B1(ram[13950]), .B2(n3612), 
        .ZN(n18191) );
  MOAI22 U27097 ( .A1(n27577), .A2(n3611), .B1(ram[13951]), .B2(n3612), 
        .ZN(n18192) );
  MOAI22 U27098 ( .A1(n29222), .A2(n3613), .B1(ram[13952]), .B2(n3614), 
        .ZN(n18193) );
  MOAI22 U27099 ( .A1(n28987), .A2(n3613), .B1(ram[13953]), .B2(n3614), 
        .ZN(n18194) );
  MOAI22 U27100 ( .A1(n28752), .A2(n3613), .B1(ram[13954]), .B2(n3614), 
        .ZN(n18195) );
  MOAI22 U27101 ( .A1(n28517), .A2(n3613), .B1(ram[13955]), .B2(n3614), 
        .ZN(n18196) );
  MOAI22 U27102 ( .A1(n28282), .A2(n3613), .B1(ram[13956]), .B2(n3614), 
        .ZN(n18197) );
  MOAI22 U27103 ( .A1(n28047), .A2(n3613), .B1(ram[13957]), .B2(n3614), 
        .ZN(n18198) );
  MOAI22 U27104 ( .A1(n27812), .A2(n3613), .B1(ram[13958]), .B2(n3614), 
        .ZN(n18199) );
  MOAI22 U27105 ( .A1(n27577), .A2(n3613), .B1(ram[13959]), .B2(n3614), 
        .ZN(n18200) );
  MOAI22 U27106 ( .A1(n29222), .A2(n3615), .B1(ram[13960]), .B2(n3616), 
        .ZN(n18201) );
  MOAI22 U27107 ( .A1(n28987), .A2(n3615), .B1(ram[13961]), .B2(n3616), 
        .ZN(n18202) );
  MOAI22 U27108 ( .A1(n28752), .A2(n3615), .B1(ram[13962]), .B2(n3616), 
        .ZN(n18203) );
  MOAI22 U27109 ( .A1(n28517), .A2(n3615), .B1(ram[13963]), .B2(n3616), 
        .ZN(n18204) );
  MOAI22 U27110 ( .A1(n28282), .A2(n3615), .B1(ram[13964]), .B2(n3616), 
        .ZN(n18205) );
  MOAI22 U27111 ( .A1(n28047), .A2(n3615), .B1(ram[13965]), .B2(n3616), 
        .ZN(n18206) );
  MOAI22 U27112 ( .A1(n27812), .A2(n3615), .B1(ram[13966]), .B2(n3616), 
        .ZN(n18207) );
  MOAI22 U27113 ( .A1(n27577), .A2(n3615), .B1(ram[13967]), .B2(n3616), 
        .ZN(n18208) );
  MOAI22 U27114 ( .A1(n29222), .A2(n3617), .B1(ram[13968]), .B2(n3618), 
        .ZN(n18209) );
  MOAI22 U27115 ( .A1(n28987), .A2(n3617), .B1(ram[13969]), .B2(n3618), 
        .ZN(n18210) );
  MOAI22 U27116 ( .A1(n28752), .A2(n3617), .B1(ram[13970]), .B2(n3618), 
        .ZN(n18211) );
  MOAI22 U27117 ( .A1(n28517), .A2(n3617), .B1(ram[13971]), .B2(n3618), 
        .ZN(n18212) );
  MOAI22 U27118 ( .A1(n28282), .A2(n3617), .B1(ram[13972]), .B2(n3618), 
        .ZN(n18213) );
  MOAI22 U27119 ( .A1(n28047), .A2(n3617), .B1(ram[13973]), .B2(n3618), 
        .ZN(n18214) );
  MOAI22 U27120 ( .A1(n27812), .A2(n3617), .B1(ram[13974]), .B2(n3618), 
        .ZN(n18215) );
  MOAI22 U27121 ( .A1(n27577), .A2(n3617), .B1(ram[13975]), .B2(n3618), 
        .ZN(n18216) );
  MOAI22 U27122 ( .A1(n29222), .A2(n3619), .B1(ram[13976]), .B2(n3620), 
        .ZN(n18217) );
  MOAI22 U27123 ( .A1(n28987), .A2(n3619), .B1(ram[13977]), .B2(n3620), 
        .ZN(n18218) );
  MOAI22 U27124 ( .A1(n28752), .A2(n3619), .B1(ram[13978]), .B2(n3620), 
        .ZN(n18219) );
  MOAI22 U27125 ( .A1(n28517), .A2(n3619), .B1(ram[13979]), .B2(n3620), 
        .ZN(n18220) );
  MOAI22 U27126 ( .A1(n28282), .A2(n3619), .B1(ram[13980]), .B2(n3620), 
        .ZN(n18221) );
  MOAI22 U27127 ( .A1(n28047), .A2(n3619), .B1(ram[13981]), .B2(n3620), 
        .ZN(n18222) );
  MOAI22 U27128 ( .A1(n27812), .A2(n3619), .B1(ram[13982]), .B2(n3620), 
        .ZN(n18223) );
  MOAI22 U27129 ( .A1(n27577), .A2(n3619), .B1(ram[13983]), .B2(n3620), 
        .ZN(n18224) );
  MOAI22 U27130 ( .A1(n29222), .A2(n3621), .B1(ram[13984]), .B2(n3622), 
        .ZN(n18225) );
  MOAI22 U27131 ( .A1(n28987), .A2(n3621), .B1(ram[13985]), .B2(n3622), 
        .ZN(n18226) );
  MOAI22 U27132 ( .A1(n28752), .A2(n3621), .B1(ram[13986]), .B2(n3622), 
        .ZN(n18227) );
  MOAI22 U27133 ( .A1(n28517), .A2(n3621), .B1(ram[13987]), .B2(n3622), 
        .ZN(n18228) );
  MOAI22 U27134 ( .A1(n28282), .A2(n3621), .B1(ram[13988]), .B2(n3622), 
        .ZN(n18229) );
  MOAI22 U27135 ( .A1(n28047), .A2(n3621), .B1(ram[13989]), .B2(n3622), 
        .ZN(n18230) );
  MOAI22 U27136 ( .A1(n27812), .A2(n3621), .B1(ram[13990]), .B2(n3622), 
        .ZN(n18231) );
  MOAI22 U27137 ( .A1(n27577), .A2(n3621), .B1(ram[13991]), .B2(n3622), 
        .ZN(n18232) );
  MOAI22 U27138 ( .A1(n29222), .A2(n3623), .B1(ram[13992]), .B2(n3624), 
        .ZN(n18233) );
  MOAI22 U27139 ( .A1(n28987), .A2(n3623), .B1(ram[13993]), .B2(n3624), 
        .ZN(n18234) );
  MOAI22 U27140 ( .A1(n28752), .A2(n3623), .B1(ram[13994]), .B2(n3624), 
        .ZN(n18235) );
  MOAI22 U27141 ( .A1(n28517), .A2(n3623), .B1(ram[13995]), .B2(n3624), 
        .ZN(n18236) );
  MOAI22 U27142 ( .A1(n28282), .A2(n3623), .B1(ram[13996]), .B2(n3624), 
        .ZN(n18237) );
  MOAI22 U27143 ( .A1(n28047), .A2(n3623), .B1(ram[13997]), .B2(n3624), 
        .ZN(n18238) );
  MOAI22 U27144 ( .A1(n27812), .A2(n3623), .B1(ram[13998]), .B2(n3624), 
        .ZN(n18239) );
  MOAI22 U27145 ( .A1(n27577), .A2(n3623), .B1(ram[13999]), .B2(n3624), 
        .ZN(n18240) );
  MOAI22 U27146 ( .A1(n29222), .A2(n3625), .B1(ram[14000]), .B2(n3626), 
        .ZN(n18241) );
  MOAI22 U27147 ( .A1(n28987), .A2(n3625), .B1(ram[14001]), .B2(n3626), 
        .ZN(n18242) );
  MOAI22 U27148 ( .A1(n28752), .A2(n3625), .B1(ram[14002]), .B2(n3626), 
        .ZN(n18243) );
  MOAI22 U27149 ( .A1(n28517), .A2(n3625), .B1(ram[14003]), .B2(n3626), 
        .ZN(n18244) );
  MOAI22 U27150 ( .A1(n28282), .A2(n3625), .B1(ram[14004]), .B2(n3626), 
        .ZN(n18245) );
  MOAI22 U27151 ( .A1(n28047), .A2(n3625), .B1(ram[14005]), .B2(n3626), 
        .ZN(n18246) );
  MOAI22 U27152 ( .A1(n27812), .A2(n3625), .B1(ram[14006]), .B2(n3626), 
        .ZN(n18247) );
  MOAI22 U27153 ( .A1(n27577), .A2(n3625), .B1(ram[14007]), .B2(n3626), 
        .ZN(n18248) );
  MOAI22 U27154 ( .A1(n29222), .A2(n3627), .B1(ram[14008]), .B2(n3628), 
        .ZN(n18249) );
  MOAI22 U27155 ( .A1(n28987), .A2(n3627), .B1(ram[14009]), .B2(n3628), 
        .ZN(n18250) );
  MOAI22 U27156 ( .A1(n28752), .A2(n3627), .B1(ram[14010]), .B2(n3628), 
        .ZN(n18251) );
  MOAI22 U27157 ( .A1(n28517), .A2(n3627), .B1(ram[14011]), .B2(n3628), 
        .ZN(n18252) );
  MOAI22 U27158 ( .A1(n28282), .A2(n3627), .B1(ram[14012]), .B2(n3628), 
        .ZN(n18253) );
  MOAI22 U27159 ( .A1(n28047), .A2(n3627), .B1(ram[14013]), .B2(n3628), 
        .ZN(n18254) );
  MOAI22 U27160 ( .A1(n27812), .A2(n3627), .B1(ram[14014]), .B2(n3628), 
        .ZN(n18255) );
  MOAI22 U27161 ( .A1(n27577), .A2(n3627), .B1(ram[14015]), .B2(n3628), 
        .ZN(n18256) );
  MOAI22 U27162 ( .A1(n29222), .A2(n3629), .B1(ram[14016]), .B2(n3630), 
        .ZN(n18257) );
  MOAI22 U27163 ( .A1(n28987), .A2(n3629), .B1(ram[14017]), .B2(n3630), 
        .ZN(n18258) );
  MOAI22 U27164 ( .A1(n28752), .A2(n3629), .B1(ram[14018]), .B2(n3630), 
        .ZN(n18259) );
  MOAI22 U27165 ( .A1(n28517), .A2(n3629), .B1(ram[14019]), .B2(n3630), 
        .ZN(n18260) );
  MOAI22 U27166 ( .A1(n28282), .A2(n3629), .B1(ram[14020]), .B2(n3630), 
        .ZN(n18261) );
  MOAI22 U27167 ( .A1(n28047), .A2(n3629), .B1(ram[14021]), .B2(n3630), 
        .ZN(n18262) );
  MOAI22 U27168 ( .A1(n27812), .A2(n3629), .B1(ram[14022]), .B2(n3630), 
        .ZN(n18263) );
  MOAI22 U27169 ( .A1(n27577), .A2(n3629), .B1(ram[14023]), .B2(n3630), 
        .ZN(n18264) );
  MOAI22 U27170 ( .A1(n29222), .A2(n3631), .B1(ram[14024]), .B2(n3632), 
        .ZN(n18265) );
  MOAI22 U27171 ( .A1(n28987), .A2(n3631), .B1(ram[14025]), .B2(n3632), 
        .ZN(n18266) );
  MOAI22 U27172 ( .A1(n28752), .A2(n3631), .B1(ram[14026]), .B2(n3632), 
        .ZN(n18267) );
  MOAI22 U27173 ( .A1(n28517), .A2(n3631), .B1(ram[14027]), .B2(n3632), 
        .ZN(n18268) );
  MOAI22 U27174 ( .A1(n28282), .A2(n3631), .B1(ram[14028]), .B2(n3632), 
        .ZN(n18269) );
  MOAI22 U27175 ( .A1(n28047), .A2(n3631), .B1(ram[14029]), .B2(n3632), 
        .ZN(n18270) );
  MOAI22 U27176 ( .A1(n27812), .A2(n3631), .B1(ram[14030]), .B2(n3632), 
        .ZN(n18271) );
  MOAI22 U27177 ( .A1(n27577), .A2(n3631), .B1(ram[14031]), .B2(n3632), 
        .ZN(n18272) );
  MOAI22 U27178 ( .A1(n29222), .A2(n3633), .B1(ram[14032]), .B2(n3634), 
        .ZN(n18273) );
  MOAI22 U27179 ( .A1(n28987), .A2(n3633), .B1(ram[14033]), .B2(n3634), 
        .ZN(n18274) );
  MOAI22 U27180 ( .A1(n28752), .A2(n3633), .B1(ram[14034]), .B2(n3634), 
        .ZN(n18275) );
  MOAI22 U27181 ( .A1(n28517), .A2(n3633), .B1(ram[14035]), .B2(n3634), 
        .ZN(n18276) );
  MOAI22 U27182 ( .A1(n28282), .A2(n3633), .B1(ram[14036]), .B2(n3634), 
        .ZN(n18277) );
  MOAI22 U27183 ( .A1(n28047), .A2(n3633), .B1(ram[14037]), .B2(n3634), 
        .ZN(n18278) );
  MOAI22 U27184 ( .A1(n27812), .A2(n3633), .B1(ram[14038]), .B2(n3634), 
        .ZN(n18279) );
  MOAI22 U27185 ( .A1(n27577), .A2(n3633), .B1(ram[14039]), .B2(n3634), 
        .ZN(n18280) );
  MOAI22 U27186 ( .A1(n29223), .A2(n3635), .B1(ram[14040]), .B2(n3636), 
        .ZN(n18281) );
  MOAI22 U27187 ( .A1(n28988), .A2(n3635), .B1(ram[14041]), .B2(n3636), 
        .ZN(n18282) );
  MOAI22 U27188 ( .A1(n28753), .A2(n3635), .B1(ram[14042]), .B2(n3636), 
        .ZN(n18283) );
  MOAI22 U27189 ( .A1(n28518), .A2(n3635), .B1(ram[14043]), .B2(n3636), 
        .ZN(n18284) );
  MOAI22 U27190 ( .A1(n28283), .A2(n3635), .B1(ram[14044]), .B2(n3636), 
        .ZN(n18285) );
  MOAI22 U27191 ( .A1(n28048), .A2(n3635), .B1(ram[14045]), .B2(n3636), 
        .ZN(n18286) );
  MOAI22 U27192 ( .A1(n27813), .A2(n3635), .B1(ram[14046]), .B2(n3636), 
        .ZN(n18287) );
  MOAI22 U27193 ( .A1(n27578), .A2(n3635), .B1(ram[14047]), .B2(n3636), 
        .ZN(n18288) );
  MOAI22 U27194 ( .A1(n29223), .A2(n3637), .B1(ram[14048]), .B2(n3638), 
        .ZN(n18289) );
  MOAI22 U27195 ( .A1(n28988), .A2(n3637), .B1(ram[14049]), .B2(n3638), 
        .ZN(n18290) );
  MOAI22 U27196 ( .A1(n28753), .A2(n3637), .B1(ram[14050]), .B2(n3638), 
        .ZN(n18291) );
  MOAI22 U27197 ( .A1(n28518), .A2(n3637), .B1(ram[14051]), .B2(n3638), 
        .ZN(n18292) );
  MOAI22 U27198 ( .A1(n28283), .A2(n3637), .B1(ram[14052]), .B2(n3638), 
        .ZN(n18293) );
  MOAI22 U27199 ( .A1(n28048), .A2(n3637), .B1(ram[14053]), .B2(n3638), 
        .ZN(n18294) );
  MOAI22 U27200 ( .A1(n27813), .A2(n3637), .B1(ram[14054]), .B2(n3638), 
        .ZN(n18295) );
  MOAI22 U27201 ( .A1(n27578), .A2(n3637), .B1(ram[14055]), .B2(n3638), 
        .ZN(n18296) );
  MOAI22 U27202 ( .A1(n29223), .A2(n3639), .B1(ram[14056]), .B2(n3640), 
        .ZN(n18297) );
  MOAI22 U27203 ( .A1(n28988), .A2(n3639), .B1(ram[14057]), .B2(n3640), 
        .ZN(n18298) );
  MOAI22 U27204 ( .A1(n28753), .A2(n3639), .B1(ram[14058]), .B2(n3640), 
        .ZN(n18299) );
  MOAI22 U27205 ( .A1(n28518), .A2(n3639), .B1(ram[14059]), .B2(n3640), 
        .ZN(n18300) );
  MOAI22 U27206 ( .A1(n28283), .A2(n3639), .B1(ram[14060]), .B2(n3640), 
        .ZN(n18301) );
  MOAI22 U27207 ( .A1(n28048), .A2(n3639), .B1(ram[14061]), .B2(n3640), 
        .ZN(n18302) );
  MOAI22 U27208 ( .A1(n27813), .A2(n3639), .B1(ram[14062]), .B2(n3640), 
        .ZN(n18303) );
  MOAI22 U27209 ( .A1(n27578), .A2(n3639), .B1(ram[14063]), .B2(n3640), 
        .ZN(n18304) );
  MOAI22 U27210 ( .A1(n29223), .A2(n3641), .B1(ram[14064]), .B2(n3642), 
        .ZN(n18305) );
  MOAI22 U27211 ( .A1(n28988), .A2(n3641), .B1(ram[14065]), .B2(n3642), 
        .ZN(n18306) );
  MOAI22 U27212 ( .A1(n28753), .A2(n3641), .B1(ram[14066]), .B2(n3642), 
        .ZN(n18307) );
  MOAI22 U27213 ( .A1(n28518), .A2(n3641), .B1(ram[14067]), .B2(n3642), 
        .ZN(n18308) );
  MOAI22 U27214 ( .A1(n28283), .A2(n3641), .B1(ram[14068]), .B2(n3642), 
        .ZN(n18309) );
  MOAI22 U27215 ( .A1(n28048), .A2(n3641), .B1(ram[14069]), .B2(n3642), 
        .ZN(n18310) );
  MOAI22 U27216 ( .A1(n27813), .A2(n3641), .B1(ram[14070]), .B2(n3642), 
        .ZN(n18311) );
  MOAI22 U27217 ( .A1(n27578), .A2(n3641), .B1(ram[14071]), .B2(n3642), 
        .ZN(n18312) );
  MOAI22 U27218 ( .A1(n29223), .A2(n3643), .B1(ram[14072]), .B2(n3644), 
        .ZN(n18313) );
  MOAI22 U27219 ( .A1(n28988), .A2(n3643), .B1(ram[14073]), .B2(n3644), 
        .ZN(n18314) );
  MOAI22 U27220 ( .A1(n28753), .A2(n3643), .B1(ram[14074]), .B2(n3644), 
        .ZN(n18315) );
  MOAI22 U27221 ( .A1(n28518), .A2(n3643), .B1(ram[14075]), .B2(n3644), 
        .ZN(n18316) );
  MOAI22 U27222 ( .A1(n28283), .A2(n3643), .B1(ram[14076]), .B2(n3644), 
        .ZN(n18317) );
  MOAI22 U27223 ( .A1(n28048), .A2(n3643), .B1(ram[14077]), .B2(n3644), 
        .ZN(n18318) );
  MOAI22 U27224 ( .A1(n27813), .A2(n3643), .B1(ram[14078]), .B2(n3644), 
        .ZN(n18319) );
  MOAI22 U27225 ( .A1(n27578), .A2(n3643), .B1(ram[14079]), .B2(n3644), 
        .ZN(n18320) );
  MOAI22 U27226 ( .A1(n29223), .A2(n3645), .B1(ram[14080]), .B2(n3646), 
        .ZN(n18321) );
  MOAI22 U27227 ( .A1(n28988), .A2(n3645), .B1(ram[14081]), .B2(n3646), 
        .ZN(n18322) );
  MOAI22 U27228 ( .A1(n28753), .A2(n3645), .B1(ram[14082]), .B2(n3646), 
        .ZN(n18323) );
  MOAI22 U27229 ( .A1(n28518), .A2(n3645), .B1(ram[14083]), .B2(n3646), 
        .ZN(n18324) );
  MOAI22 U27230 ( .A1(n28283), .A2(n3645), .B1(ram[14084]), .B2(n3646), 
        .ZN(n18325) );
  MOAI22 U27231 ( .A1(n28048), .A2(n3645), .B1(ram[14085]), .B2(n3646), 
        .ZN(n18326) );
  MOAI22 U27232 ( .A1(n27813), .A2(n3645), .B1(ram[14086]), .B2(n3646), 
        .ZN(n18327) );
  MOAI22 U27233 ( .A1(n27578), .A2(n3645), .B1(ram[14087]), .B2(n3646), 
        .ZN(n18328) );
  MOAI22 U27234 ( .A1(n29223), .A2(n3647), .B1(ram[14088]), .B2(n3648), 
        .ZN(n18329) );
  MOAI22 U27235 ( .A1(n28988), .A2(n3647), .B1(ram[14089]), .B2(n3648), 
        .ZN(n18330) );
  MOAI22 U27236 ( .A1(n28753), .A2(n3647), .B1(ram[14090]), .B2(n3648), 
        .ZN(n18331) );
  MOAI22 U27237 ( .A1(n28518), .A2(n3647), .B1(ram[14091]), .B2(n3648), 
        .ZN(n18332) );
  MOAI22 U27238 ( .A1(n28283), .A2(n3647), .B1(ram[14092]), .B2(n3648), 
        .ZN(n18333) );
  MOAI22 U27239 ( .A1(n28048), .A2(n3647), .B1(ram[14093]), .B2(n3648), 
        .ZN(n18334) );
  MOAI22 U27240 ( .A1(n27813), .A2(n3647), .B1(ram[14094]), .B2(n3648), 
        .ZN(n18335) );
  MOAI22 U27241 ( .A1(n27578), .A2(n3647), .B1(ram[14095]), .B2(n3648), 
        .ZN(n18336) );
  MOAI22 U27242 ( .A1(n29223), .A2(n3649), .B1(ram[14096]), .B2(n3650), 
        .ZN(n18337) );
  MOAI22 U27243 ( .A1(n28988), .A2(n3649), .B1(ram[14097]), .B2(n3650), 
        .ZN(n18338) );
  MOAI22 U27244 ( .A1(n28753), .A2(n3649), .B1(ram[14098]), .B2(n3650), 
        .ZN(n18339) );
  MOAI22 U27245 ( .A1(n28518), .A2(n3649), .B1(ram[14099]), .B2(n3650), 
        .ZN(n18340) );
  MOAI22 U27246 ( .A1(n28283), .A2(n3649), .B1(ram[14100]), .B2(n3650), 
        .ZN(n18341) );
  MOAI22 U27247 ( .A1(n28048), .A2(n3649), .B1(ram[14101]), .B2(n3650), 
        .ZN(n18342) );
  MOAI22 U27248 ( .A1(n27813), .A2(n3649), .B1(ram[14102]), .B2(n3650), 
        .ZN(n18343) );
  MOAI22 U27249 ( .A1(n27578), .A2(n3649), .B1(ram[14103]), .B2(n3650), 
        .ZN(n18344) );
  MOAI22 U27250 ( .A1(n29223), .A2(n3651), .B1(ram[14104]), .B2(n3652), 
        .ZN(n18345) );
  MOAI22 U27251 ( .A1(n28988), .A2(n3651), .B1(ram[14105]), .B2(n3652), 
        .ZN(n18346) );
  MOAI22 U27252 ( .A1(n28753), .A2(n3651), .B1(ram[14106]), .B2(n3652), 
        .ZN(n18347) );
  MOAI22 U27253 ( .A1(n28518), .A2(n3651), .B1(ram[14107]), .B2(n3652), 
        .ZN(n18348) );
  MOAI22 U27254 ( .A1(n28283), .A2(n3651), .B1(ram[14108]), .B2(n3652), 
        .ZN(n18349) );
  MOAI22 U27255 ( .A1(n28048), .A2(n3651), .B1(ram[14109]), .B2(n3652), 
        .ZN(n18350) );
  MOAI22 U27256 ( .A1(n27813), .A2(n3651), .B1(ram[14110]), .B2(n3652), 
        .ZN(n18351) );
  MOAI22 U27257 ( .A1(n27578), .A2(n3651), .B1(ram[14111]), .B2(n3652), 
        .ZN(n18352) );
  MOAI22 U27258 ( .A1(n29223), .A2(n3653), .B1(ram[14112]), .B2(n3654), 
        .ZN(n18353) );
  MOAI22 U27259 ( .A1(n28988), .A2(n3653), .B1(ram[14113]), .B2(n3654), 
        .ZN(n18354) );
  MOAI22 U27260 ( .A1(n28753), .A2(n3653), .B1(ram[14114]), .B2(n3654), 
        .ZN(n18355) );
  MOAI22 U27261 ( .A1(n28518), .A2(n3653), .B1(ram[14115]), .B2(n3654), 
        .ZN(n18356) );
  MOAI22 U27262 ( .A1(n28283), .A2(n3653), .B1(ram[14116]), .B2(n3654), 
        .ZN(n18357) );
  MOAI22 U27263 ( .A1(n28048), .A2(n3653), .B1(ram[14117]), .B2(n3654), 
        .ZN(n18358) );
  MOAI22 U27264 ( .A1(n27813), .A2(n3653), .B1(ram[14118]), .B2(n3654), 
        .ZN(n18359) );
  MOAI22 U27265 ( .A1(n27578), .A2(n3653), .B1(ram[14119]), .B2(n3654), 
        .ZN(n18360) );
  MOAI22 U27266 ( .A1(n29223), .A2(n3655), .B1(ram[14120]), .B2(n3656), 
        .ZN(n18361) );
  MOAI22 U27267 ( .A1(n28988), .A2(n3655), .B1(ram[14121]), .B2(n3656), 
        .ZN(n18362) );
  MOAI22 U27268 ( .A1(n28753), .A2(n3655), .B1(ram[14122]), .B2(n3656), 
        .ZN(n18363) );
  MOAI22 U27269 ( .A1(n28518), .A2(n3655), .B1(ram[14123]), .B2(n3656), 
        .ZN(n18364) );
  MOAI22 U27270 ( .A1(n28283), .A2(n3655), .B1(ram[14124]), .B2(n3656), 
        .ZN(n18365) );
  MOAI22 U27271 ( .A1(n28048), .A2(n3655), .B1(ram[14125]), .B2(n3656), 
        .ZN(n18366) );
  MOAI22 U27272 ( .A1(n27813), .A2(n3655), .B1(ram[14126]), .B2(n3656), 
        .ZN(n18367) );
  MOAI22 U27273 ( .A1(n27578), .A2(n3655), .B1(ram[14127]), .B2(n3656), 
        .ZN(n18368) );
  MOAI22 U27274 ( .A1(n29223), .A2(n3657), .B1(ram[14128]), .B2(n3658), 
        .ZN(n18369) );
  MOAI22 U27275 ( .A1(n28988), .A2(n3657), .B1(ram[14129]), .B2(n3658), 
        .ZN(n18370) );
  MOAI22 U27276 ( .A1(n28753), .A2(n3657), .B1(ram[14130]), .B2(n3658), 
        .ZN(n18371) );
  MOAI22 U27277 ( .A1(n28518), .A2(n3657), .B1(ram[14131]), .B2(n3658), 
        .ZN(n18372) );
  MOAI22 U27278 ( .A1(n28283), .A2(n3657), .B1(ram[14132]), .B2(n3658), 
        .ZN(n18373) );
  MOAI22 U27279 ( .A1(n28048), .A2(n3657), .B1(ram[14133]), .B2(n3658), 
        .ZN(n18374) );
  MOAI22 U27280 ( .A1(n27813), .A2(n3657), .B1(ram[14134]), .B2(n3658), 
        .ZN(n18375) );
  MOAI22 U27281 ( .A1(n27578), .A2(n3657), .B1(ram[14135]), .B2(n3658), 
        .ZN(n18376) );
  MOAI22 U27282 ( .A1(n29223), .A2(n3659), .B1(ram[14136]), .B2(n3660), 
        .ZN(n18377) );
  MOAI22 U27283 ( .A1(n28988), .A2(n3659), .B1(ram[14137]), .B2(n3660), 
        .ZN(n18378) );
  MOAI22 U27284 ( .A1(n28753), .A2(n3659), .B1(ram[14138]), .B2(n3660), 
        .ZN(n18379) );
  MOAI22 U27285 ( .A1(n28518), .A2(n3659), .B1(ram[14139]), .B2(n3660), 
        .ZN(n18380) );
  MOAI22 U27286 ( .A1(n28283), .A2(n3659), .B1(ram[14140]), .B2(n3660), 
        .ZN(n18381) );
  MOAI22 U27287 ( .A1(n28048), .A2(n3659), .B1(ram[14141]), .B2(n3660), 
        .ZN(n18382) );
  MOAI22 U27288 ( .A1(n27813), .A2(n3659), .B1(ram[14142]), .B2(n3660), 
        .ZN(n18383) );
  MOAI22 U27289 ( .A1(n27578), .A2(n3659), .B1(ram[14143]), .B2(n3660), 
        .ZN(n18384) );
  MOAI22 U27290 ( .A1(n29224), .A2(n3661), .B1(ram[14144]), .B2(n3662), 
        .ZN(n18385) );
  MOAI22 U27291 ( .A1(n28989), .A2(n3661), .B1(ram[14145]), .B2(n3662), 
        .ZN(n18386) );
  MOAI22 U27292 ( .A1(n28754), .A2(n3661), .B1(ram[14146]), .B2(n3662), 
        .ZN(n18387) );
  MOAI22 U27293 ( .A1(n28519), .A2(n3661), .B1(ram[14147]), .B2(n3662), 
        .ZN(n18388) );
  MOAI22 U27294 ( .A1(n28284), .A2(n3661), .B1(ram[14148]), .B2(n3662), 
        .ZN(n18389) );
  MOAI22 U27295 ( .A1(n28049), .A2(n3661), .B1(ram[14149]), .B2(n3662), 
        .ZN(n18390) );
  MOAI22 U27296 ( .A1(n27814), .A2(n3661), .B1(ram[14150]), .B2(n3662), 
        .ZN(n18391) );
  MOAI22 U27297 ( .A1(n27579), .A2(n3661), .B1(ram[14151]), .B2(n3662), 
        .ZN(n18392) );
  MOAI22 U27298 ( .A1(n29224), .A2(n3663), .B1(ram[14152]), .B2(n3664), 
        .ZN(n18393) );
  MOAI22 U27299 ( .A1(n28989), .A2(n3663), .B1(ram[14153]), .B2(n3664), 
        .ZN(n18394) );
  MOAI22 U27300 ( .A1(n28754), .A2(n3663), .B1(ram[14154]), .B2(n3664), 
        .ZN(n18395) );
  MOAI22 U27301 ( .A1(n28519), .A2(n3663), .B1(ram[14155]), .B2(n3664), 
        .ZN(n18396) );
  MOAI22 U27302 ( .A1(n28284), .A2(n3663), .B1(ram[14156]), .B2(n3664), 
        .ZN(n18397) );
  MOAI22 U27303 ( .A1(n28049), .A2(n3663), .B1(ram[14157]), .B2(n3664), 
        .ZN(n18398) );
  MOAI22 U27304 ( .A1(n27814), .A2(n3663), .B1(ram[14158]), .B2(n3664), 
        .ZN(n18399) );
  MOAI22 U27305 ( .A1(n27579), .A2(n3663), .B1(ram[14159]), .B2(n3664), 
        .ZN(n18400) );
  MOAI22 U27306 ( .A1(n29224), .A2(n3665), .B1(ram[14160]), .B2(n3666), 
        .ZN(n18401) );
  MOAI22 U27307 ( .A1(n28989), .A2(n3665), .B1(ram[14161]), .B2(n3666), 
        .ZN(n18402) );
  MOAI22 U27308 ( .A1(n28754), .A2(n3665), .B1(ram[14162]), .B2(n3666), 
        .ZN(n18403) );
  MOAI22 U27309 ( .A1(n28519), .A2(n3665), .B1(ram[14163]), .B2(n3666), 
        .ZN(n18404) );
  MOAI22 U27310 ( .A1(n28284), .A2(n3665), .B1(ram[14164]), .B2(n3666), 
        .ZN(n18405) );
  MOAI22 U27311 ( .A1(n28049), .A2(n3665), .B1(ram[14165]), .B2(n3666), 
        .ZN(n18406) );
  MOAI22 U27312 ( .A1(n27814), .A2(n3665), .B1(ram[14166]), .B2(n3666), 
        .ZN(n18407) );
  MOAI22 U27313 ( .A1(n27579), .A2(n3665), .B1(ram[14167]), .B2(n3666), 
        .ZN(n18408) );
  MOAI22 U27314 ( .A1(n29224), .A2(n3667), .B1(ram[14168]), .B2(n3668), 
        .ZN(n18409) );
  MOAI22 U27315 ( .A1(n28989), .A2(n3667), .B1(ram[14169]), .B2(n3668), 
        .ZN(n18410) );
  MOAI22 U27316 ( .A1(n28754), .A2(n3667), .B1(ram[14170]), .B2(n3668), 
        .ZN(n18411) );
  MOAI22 U27317 ( .A1(n28519), .A2(n3667), .B1(ram[14171]), .B2(n3668), 
        .ZN(n18412) );
  MOAI22 U27318 ( .A1(n28284), .A2(n3667), .B1(ram[14172]), .B2(n3668), 
        .ZN(n18413) );
  MOAI22 U27319 ( .A1(n28049), .A2(n3667), .B1(ram[14173]), .B2(n3668), 
        .ZN(n18414) );
  MOAI22 U27320 ( .A1(n27814), .A2(n3667), .B1(ram[14174]), .B2(n3668), 
        .ZN(n18415) );
  MOAI22 U27321 ( .A1(n27579), .A2(n3667), .B1(ram[14175]), .B2(n3668), 
        .ZN(n18416) );
  MOAI22 U27322 ( .A1(n29224), .A2(n3669), .B1(ram[14176]), .B2(n3670), 
        .ZN(n18417) );
  MOAI22 U27323 ( .A1(n28989), .A2(n3669), .B1(ram[14177]), .B2(n3670), 
        .ZN(n18418) );
  MOAI22 U27324 ( .A1(n28754), .A2(n3669), .B1(ram[14178]), .B2(n3670), 
        .ZN(n18419) );
  MOAI22 U27325 ( .A1(n28519), .A2(n3669), .B1(ram[14179]), .B2(n3670), 
        .ZN(n18420) );
  MOAI22 U27326 ( .A1(n28284), .A2(n3669), .B1(ram[14180]), .B2(n3670), 
        .ZN(n18421) );
  MOAI22 U27327 ( .A1(n28049), .A2(n3669), .B1(ram[14181]), .B2(n3670), 
        .ZN(n18422) );
  MOAI22 U27328 ( .A1(n27814), .A2(n3669), .B1(ram[14182]), .B2(n3670), 
        .ZN(n18423) );
  MOAI22 U27329 ( .A1(n27579), .A2(n3669), .B1(ram[14183]), .B2(n3670), 
        .ZN(n18424) );
  MOAI22 U27330 ( .A1(n29224), .A2(n3671), .B1(ram[14184]), .B2(n3672), 
        .ZN(n18425) );
  MOAI22 U27331 ( .A1(n28989), .A2(n3671), .B1(ram[14185]), .B2(n3672), 
        .ZN(n18426) );
  MOAI22 U27332 ( .A1(n28754), .A2(n3671), .B1(ram[14186]), .B2(n3672), 
        .ZN(n18427) );
  MOAI22 U27333 ( .A1(n28519), .A2(n3671), .B1(ram[14187]), .B2(n3672), 
        .ZN(n18428) );
  MOAI22 U27334 ( .A1(n28284), .A2(n3671), .B1(ram[14188]), .B2(n3672), 
        .ZN(n18429) );
  MOAI22 U27335 ( .A1(n28049), .A2(n3671), .B1(ram[14189]), .B2(n3672), 
        .ZN(n18430) );
  MOAI22 U27336 ( .A1(n27814), .A2(n3671), .B1(ram[14190]), .B2(n3672), 
        .ZN(n18431) );
  MOAI22 U27337 ( .A1(n27579), .A2(n3671), .B1(ram[14191]), .B2(n3672), 
        .ZN(n18432) );
  MOAI22 U27338 ( .A1(n29224), .A2(n3673), .B1(ram[14192]), .B2(n3674), 
        .ZN(n18433) );
  MOAI22 U27339 ( .A1(n28989), .A2(n3673), .B1(ram[14193]), .B2(n3674), 
        .ZN(n18434) );
  MOAI22 U27340 ( .A1(n28754), .A2(n3673), .B1(ram[14194]), .B2(n3674), 
        .ZN(n18435) );
  MOAI22 U27341 ( .A1(n28519), .A2(n3673), .B1(ram[14195]), .B2(n3674), 
        .ZN(n18436) );
  MOAI22 U27342 ( .A1(n28284), .A2(n3673), .B1(ram[14196]), .B2(n3674), 
        .ZN(n18437) );
  MOAI22 U27343 ( .A1(n28049), .A2(n3673), .B1(ram[14197]), .B2(n3674), 
        .ZN(n18438) );
  MOAI22 U27344 ( .A1(n27814), .A2(n3673), .B1(ram[14198]), .B2(n3674), 
        .ZN(n18439) );
  MOAI22 U27345 ( .A1(n27579), .A2(n3673), .B1(ram[14199]), .B2(n3674), 
        .ZN(n18440) );
  MOAI22 U27346 ( .A1(n29224), .A2(n3675), .B1(ram[14200]), .B2(n3676), 
        .ZN(n18441) );
  MOAI22 U27347 ( .A1(n28989), .A2(n3675), .B1(ram[14201]), .B2(n3676), 
        .ZN(n18442) );
  MOAI22 U27348 ( .A1(n28754), .A2(n3675), .B1(ram[14202]), .B2(n3676), 
        .ZN(n18443) );
  MOAI22 U27349 ( .A1(n28519), .A2(n3675), .B1(ram[14203]), .B2(n3676), 
        .ZN(n18444) );
  MOAI22 U27350 ( .A1(n28284), .A2(n3675), .B1(ram[14204]), .B2(n3676), 
        .ZN(n18445) );
  MOAI22 U27351 ( .A1(n28049), .A2(n3675), .B1(ram[14205]), .B2(n3676), 
        .ZN(n18446) );
  MOAI22 U27352 ( .A1(n27814), .A2(n3675), .B1(ram[14206]), .B2(n3676), 
        .ZN(n18447) );
  MOAI22 U27353 ( .A1(n27579), .A2(n3675), .B1(ram[14207]), .B2(n3676), 
        .ZN(n18448) );
  MOAI22 U27354 ( .A1(n29224), .A2(n3677), .B1(ram[14208]), .B2(n3678), 
        .ZN(n18449) );
  MOAI22 U27355 ( .A1(n28989), .A2(n3677), .B1(ram[14209]), .B2(n3678), 
        .ZN(n18450) );
  MOAI22 U27356 ( .A1(n28754), .A2(n3677), .B1(ram[14210]), .B2(n3678), 
        .ZN(n18451) );
  MOAI22 U27357 ( .A1(n28519), .A2(n3677), .B1(ram[14211]), .B2(n3678), 
        .ZN(n18452) );
  MOAI22 U27358 ( .A1(n28284), .A2(n3677), .B1(ram[14212]), .B2(n3678), 
        .ZN(n18453) );
  MOAI22 U27359 ( .A1(n28049), .A2(n3677), .B1(ram[14213]), .B2(n3678), 
        .ZN(n18454) );
  MOAI22 U27360 ( .A1(n27814), .A2(n3677), .B1(ram[14214]), .B2(n3678), 
        .ZN(n18455) );
  MOAI22 U27361 ( .A1(n27579), .A2(n3677), .B1(ram[14215]), .B2(n3678), 
        .ZN(n18456) );
  MOAI22 U27362 ( .A1(n29224), .A2(n3679), .B1(ram[14216]), .B2(n3680), 
        .ZN(n18457) );
  MOAI22 U27363 ( .A1(n28989), .A2(n3679), .B1(ram[14217]), .B2(n3680), 
        .ZN(n18458) );
  MOAI22 U27364 ( .A1(n28754), .A2(n3679), .B1(ram[14218]), .B2(n3680), 
        .ZN(n18459) );
  MOAI22 U27365 ( .A1(n28519), .A2(n3679), .B1(ram[14219]), .B2(n3680), 
        .ZN(n18460) );
  MOAI22 U27366 ( .A1(n28284), .A2(n3679), .B1(ram[14220]), .B2(n3680), 
        .ZN(n18461) );
  MOAI22 U27367 ( .A1(n28049), .A2(n3679), .B1(ram[14221]), .B2(n3680), 
        .ZN(n18462) );
  MOAI22 U27368 ( .A1(n27814), .A2(n3679), .B1(ram[14222]), .B2(n3680), 
        .ZN(n18463) );
  MOAI22 U27369 ( .A1(n27579), .A2(n3679), .B1(ram[14223]), .B2(n3680), 
        .ZN(n18464) );
  MOAI22 U27370 ( .A1(n29224), .A2(n3681), .B1(ram[14224]), .B2(n3682), 
        .ZN(n18465) );
  MOAI22 U27371 ( .A1(n28989), .A2(n3681), .B1(ram[14225]), .B2(n3682), 
        .ZN(n18466) );
  MOAI22 U27372 ( .A1(n28754), .A2(n3681), .B1(ram[14226]), .B2(n3682), 
        .ZN(n18467) );
  MOAI22 U27373 ( .A1(n28519), .A2(n3681), .B1(ram[14227]), .B2(n3682), 
        .ZN(n18468) );
  MOAI22 U27374 ( .A1(n28284), .A2(n3681), .B1(ram[14228]), .B2(n3682), 
        .ZN(n18469) );
  MOAI22 U27375 ( .A1(n28049), .A2(n3681), .B1(ram[14229]), .B2(n3682), 
        .ZN(n18470) );
  MOAI22 U27376 ( .A1(n27814), .A2(n3681), .B1(ram[14230]), .B2(n3682), 
        .ZN(n18471) );
  MOAI22 U27377 ( .A1(n27579), .A2(n3681), .B1(ram[14231]), .B2(n3682), 
        .ZN(n18472) );
  MOAI22 U27378 ( .A1(n29224), .A2(n3683), .B1(ram[14232]), .B2(n3684), 
        .ZN(n18473) );
  MOAI22 U27379 ( .A1(n28989), .A2(n3683), .B1(ram[14233]), .B2(n3684), 
        .ZN(n18474) );
  MOAI22 U27380 ( .A1(n28754), .A2(n3683), .B1(ram[14234]), .B2(n3684), 
        .ZN(n18475) );
  MOAI22 U27381 ( .A1(n28519), .A2(n3683), .B1(ram[14235]), .B2(n3684), 
        .ZN(n18476) );
  MOAI22 U27382 ( .A1(n28284), .A2(n3683), .B1(ram[14236]), .B2(n3684), 
        .ZN(n18477) );
  MOAI22 U27383 ( .A1(n28049), .A2(n3683), .B1(ram[14237]), .B2(n3684), 
        .ZN(n18478) );
  MOAI22 U27384 ( .A1(n27814), .A2(n3683), .B1(ram[14238]), .B2(n3684), 
        .ZN(n18479) );
  MOAI22 U27385 ( .A1(n27579), .A2(n3683), .B1(ram[14239]), .B2(n3684), 
        .ZN(n18480) );
  MOAI22 U27386 ( .A1(n29224), .A2(n3685), .B1(ram[14240]), .B2(n3686), 
        .ZN(n18481) );
  MOAI22 U27387 ( .A1(n28989), .A2(n3685), .B1(ram[14241]), .B2(n3686), 
        .ZN(n18482) );
  MOAI22 U27388 ( .A1(n28754), .A2(n3685), .B1(ram[14242]), .B2(n3686), 
        .ZN(n18483) );
  MOAI22 U27389 ( .A1(n28519), .A2(n3685), .B1(ram[14243]), .B2(n3686), 
        .ZN(n18484) );
  MOAI22 U27390 ( .A1(n28284), .A2(n3685), .B1(ram[14244]), .B2(n3686), 
        .ZN(n18485) );
  MOAI22 U27391 ( .A1(n28049), .A2(n3685), .B1(ram[14245]), .B2(n3686), 
        .ZN(n18486) );
  MOAI22 U27392 ( .A1(n27814), .A2(n3685), .B1(ram[14246]), .B2(n3686), 
        .ZN(n18487) );
  MOAI22 U27393 ( .A1(n27579), .A2(n3685), .B1(ram[14247]), .B2(n3686), 
        .ZN(n18488) );
  MOAI22 U27394 ( .A1(n29225), .A2(n3687), .B1(ram[14248]), .B2(n3688), 
        .ZN(n18489) );
  MOAI22 U27395 ( .A1(n28990), .A2(n3687), .B1(ram[14249]), .B2(n3688), 
        .ZN(n18490) );
  MOAI22 U27396 ( .A1(n28755), .A2(n3687), .B1(ram[14250]), .B2(n3688), 
        .ZN(n18491) );
  MOAI22 U27397 ( .A1(n28520), .A2(n3687), .B1(ram[14251]), .B2(n3688), 
        .ZN(n18492) );
  MOAI22 U27398 ( .A1(n28285), .A2(n3687), .B1(ram[14252]), .B2(n3688), 
        .ZN(n18493) );
  MOAI22 U27399 ( .A1(n28050), .A2(n3687), .B1(ram[14253]), .B2(n3688), 
        .ZN(n18494) );
  MOAI22 U27400 ( .A1(n27815), .A2(n3687), .B1(ram[14254]), .B2(n3688), 
        .ZN(n18495) );
  MOAI22 U27401 ( .A1(n27580), .A2(n3687), .B1(ram[14255]), .B2(n3688), 
        .ZN(n18496) );
  MOAI22 U27402 ( .A1(n29225), .A2(n3689), .B1(ram[14256]), .B2(n3690), 
        .ZN(n18497) );
  MOAI22 U27403 ( .A1(n28990), .A2(n3689), .B1(ram[14257]), .B2(n3690), 
        .ZN(n18498) );
  MOAI22 U27404 ( .A1(n28755), .A2(n3689), .B1(ram[14258]), .B2(n3690), 
        .ZN(n18499) );
  MOAI22 U27405 ( .A1(n28520), .A2(n3689), .B1(ram[14259]), .B2(n3690), 
        .ZN(n18500) );
  MOAI22 U27406 ( .A1(n28285), .A2(n3689), .B1(ram[14260]), .B2(n3690), 
        .ZN(n18501) );
  MOAI22 U27407 ( .A1(n28050), .A2(n3689), .B1(ram[14261]), .B2(n3690), 
        .ZN(n18502) );
  MOAI22 U27408 ( .A1(n27815), .A2(n3689), .B1(ram[14262]), .B2(n3690), 
        .ZN(n18503) );
  MOAI22 U27409 ( .A1(n27580), .A2(n3689), .B1(ram[14263]), .B2(n3690), 
        .ZN(n18504) );
  MOAI22 U27410 ( .A1(n29225), .A2(n3691), .B1(ram[14264]), .B2(n3692), 
        .ZN(n18505) );
  MOAI22 U27411 ( .A1(n28990), .A2(n3691), .B1(ram[14265]), .B2(n3692), 
        .ZN(n18506) );
  MOAI22 U27412 ( .A1(n28755), .A2(n3691), .B1(ram[14266]), .B2(n3692), 
        .ZN(n18507) );
  MOAI22 U27413 ( .A1(n28520), .A2(n3691), .B1(ram[14267]), .B2(n3692), 
        .ZN(n18508) );
  MOAI22 U27414 ( .A1(n28285), .A2(n3691), .B1(ram[14268]), .B2(n3692), 
        .ZN(n18509) );
  MOAI22 U27415 ( .A1(n28050), .A2(n3691), .B1(ram[14269]), .B2(n3692), 
        .ZN(n18510) );
  MOAI22 U27416 ( .A1(n27815), .A2(n3691), .B1(ram[14270]), .B2(n3692), 
        .ZN(n18511) );
  MOAI22 U27417 ( .A1(n27580), .A2(n3691), .B1(ram[14271]), .B2(n3692), 
        .ZN(n18512) );
  MOAI22 U27418 ( .A1(n29225), .A2(n3693), .B1(ram[14272]), .B2(n3694), 
        .ZN(n18513) );
  MOAI22 U27419 ( .A1(n28990), .A2(n3693), .B1(ram[14273]), .B2(n3694), 
        .ZN(n18514) );
  MOAI22 U27420 ( .A1(n28755), .A2(n3693), .B1(ram[14274]), .B2(n3694), 
        .ZN(n18515) );
  MOAI22 U27421 ( .A1(n28520), .A2(n3693), .B1(ram[14275]), .B2(n3694), 
        .ZN(n18516) );
  MOAI22 U27422 ( .A1(n28285), .A2(n3693), .B1(ram[14276]), .B2(n3694), 
        .ZN(n18517) );
  MOAI22 U27423 ( .A1(n28050), .A2(n3693), .B1(ram[14277]), .B2(n3694), 
        .ZN(n18518) );
  MOAI22 U27424 ( .A1(n27815), .A2(n3693), .B1(ram[14278]), .B2(n3694), 
        .ZN(n18519) );
  MOAI22 U27425 ( .A1(n27580), .A2(n3693), .B1(ram[14279]), .B2(n3694), 
        .ZN(n18520) );
  MOAI22 U27426 ( .A1(n29225), .A2(n3695), .B1(ram[14280]), .B2(n3696), 
        .ZN(n18521) );
  MOAI22 U27427 ( .A1(n28990), .A2(n3695), .B1(ram[14281]), .B2(n3696), 
        .ZN(n18522) );
  MOAI22 U27428 ( .A1(n28755), .A2(n3695), .B1(ram[14282]), .B2(n3696), 
        .ZN(n18523) );
  MOAI22 U27429 ( .A1(n28520), .A2(n3695), .B1(ram[14283]), .B2(n3696), 
        .ZN(n18524) );
  MOAI22 U27430 ( .A1(n28285), .A2(n3695), .B1(ram[14284]), .B2(n3696), 
        .ZN(n18525) );
  MOAI22 U27431 ( .A1(n28050), .A2(n3695), .B1(ram[14285]), .B2(n3696), 
        .ZN(n18526) );
  MOAI22 U27432 ( .A1(n27815), .A2(n3695), .B1(ram[14286]), .B2(n3696), 
        .ZN(n18527) );
  MOAI22 U27433 ( .A1(n27580), .A2(n3695), .B1(ram[14287]), .B2(n3696), 
        .ZN(n18528) );
  MOAI22 U27434 ( .A1(n29225), .A2(n3697), .B1(ram[14288]), .B2(n3698), 
        .ZN(n18529) );
  MOAI22 U27435 ( .A1(n28990), .A2(n3697), .B1(ram[14289]), .B2(n3698), 
        .ZN(n18530) );
  MOAI22 U27436 ( .A1(n28755), .A2(n3697), .B1(ram[14290]), .B2(n3698), 
        .ZN(n18531) );
  MOAI22 U27437 ( .A1(n28520), .A2(n3697), .B1(ram[14291]), .B2(n3698), 
        .ZN(n18532) );
  MOAI22 U27438 ( .A1(n28285), .A2(n3697), .B1(ram[14292]), .B2(n3698), 
        .ZN(n18533) );
  MOAI22 U27439 ( .A1(n28050), .A2(n3697), .B1(ram[14293]), .B2(n3698), 
        .ZN(n18534) );
  MOAI22 U27440 ( .A1(n27815), .A2(n3697), .B1(ram[14294]), .B2(n3698), 
        .ZN(n18535) );
  MOAI22 U27441 ( .A1(n27580), .A2(n3697), .B1(ram[14295]), .B2(n3698), 
        .ZN(n18536) );
  MOAI22 U27442 ( .A1(n29225), .A2(n3699), .B1(ram[14296]), .B2(n3700), 
        .ZN(n18537) );
  MOAI22 U27443 ( .A1(n28990), .A2(n3699), .B1(ram[14297]), .B2(n3700), 
        .ZN(n18538) );
  MOAI22 U27444 ( .A1(n28755), .A2(n3699), .B1(ram[14298]), .B2(n3700), 
        .ZN(n18539) );
  MOAI22 U27445 ( .A1(n28520), .A2(n3699), .B1(ram[14299]), .B2(n3700), 
        .ZN(n18540) );
  MOAI22 U27446 ( .A1(n28285), .A2(n3699), .B1(ram[14300]), .B2(n3700), 
        .ZN(n18541) );
  MOAI22 U27447 ( .A1(n28050), .A2(n3699), .B1(ram[14301]), .B2(n3700), 
        .ZN(n18542) );
  MOAI22 U27448 ( .A1(n27815), .A2(n3699), .B1(ram[14302]), .B2(n3700), 
        .ZN(n18543) );
  MOAI22 U27449 ( .A1(n27580), .A2(n3699), .B1(ram[14303]), .B2(n3700), 
        .ZN(n18544) );
  MOAI22 U27450 ( .A1(n29225), .A2(n3701), .B1(ram[14304]), .B2(n3702), 
        .ZN(n18545) );
  MOAI22 U27451 ( .A1(n28990), .A2(n3701), .B1(ram[14305]), .B2(n3702), 
        .ZN(n18546) );
  MOAI22 U27452 ( .A1(n28755), .A2(n3701), .B1(ram[14306]), .B2(n3702), 
        .ZN(n18547) );
  MOAI22 U27453 ( .A1(n28520), .A2(n3701), .B1(ram[14307]), .B2(n3702), 
        .ZN(n18548) );
  MOAI22 U27454 ( .A1(n28285), .A2(n3701), .B1(ram[14308]), .B2(n3702), 
        .ZN(n18549) );
  MOAI22 U27455 ( .A1(n28050), .A2(n3701), .B1(ram[14309]), .B2(n3702), 
        .ZN(n18550) );
  MOAI22 U27456 ( .A1(n27815), .A2(n3701), .B1(ram[14310]), .B2(n3702), 
        .ZN(n18551) );
  MOAI22 U27457 ( .A1(n27580), .A2(n3701), .B1(ram[14311]), .B2(n3702), 
        .ZN(n18552) );
  MOAI22 U27458 ( .A1(n29225), .A2(n3703), .B1(ram[14312]), .B2(n3704), 
        .ZN(n18553) );
  MOAI22 U27459 ( .A1(n28990), .A2(n3703), .B1(ram[14313]), .B2(n3704), 
        .ZN(n18554) );
  MOAI22 U27460 ( .A1(n28755), .A2(n3703), .B1(ram[14314]), .B2(n3704), 
        .ZN(n18555) );
  MOAI22 U27461 ( .A1(n28520), .A2(n3703), .B1(ram[14315]), .B2(n3704), 
        .ZN(n18556) );
  MOAI22 U27462 ( .A1(n28285), .A2(n3703), .B1(ram[14316]), .B2(n3704), 
        .ZN(n18557) );
  MOAI22 U27463 ( .A1(n28050), .A2(n3703), .B1(ram[14317]), .B2(n3704), 
        .ZN(n18558) );
  MOAI22 U27464 ( .A1(n27815), .A2(n3703), .B1(ram[14318]), .B2(n3704), 
        .ZN(n18559) );
  MOAI22 U27465 ( .A1(n27580), .A2(n3703), .B1(ram[14319]), .B2(n3704), 
        .ZN(n18560) );
  MOAI22 U27466 ( .A1(n29225), .A2(n3705), .B1(ram[14320]), .B2(n3706), 
        .ZN(n18561) );
  MOAI22 U27467 ( .A1(n28990), .A2(n3705), .B1(ram[14321]), .B2(n3706), 
        .ZN(n18562) );
  MOAI22 U27468 ( .A1(n28755), .A2(n3705), .B1(ram[14322]), .B2(n3706), 
        .ZN(n18563) );
  MOAI22 U27469 ( .A1(n28520), .A2(n3705), .B1(ram[14323]), .B2(n3706), 
        .ZN(n18564) );
  MOAI22 U27470 ( .A1(n28285), .A2(n3705), .B1(ram[14324]), .B2(n3706), 
        .ZN(n18565) );
  MOAI22 U27471 ( .A1(n28050), .A2(n3705), .B1(ram[14325]), .B2(n3706), 
        .ZN(n18566) );
  MOAI22 U27472 ( .A1(n27815), .A2(n3705), .B1(ram[14326]), .B2(n3706), 
        .ZN(n18567) );
  MOAI22 U27473 ( .A1(n27580), .A2(n3705), .B1(ram[14327]), .B2(n3706), 
        .ZN(n18568) );
  MOAI22 U27474 ( .A1(n29225), .A2(n3707), .B1(ram[14328]), .B2(n3708), 
        .ZN(n18569) );
  MOAI22 U27475 ( .A1(n28990), .A2(n3707), .B1(ram[14329]), .B2(n3708), 
        .ZN(n18570) );
  MOAI22 U27476 ( .A1(n28755), .A2(n3707), .B1(ram[14330]), .B2(n3708), 
        .ZN(n18571) );
  MOAI22 U27477 ( .A1(n28520), .A2(n3707), .B1(ram[14331]), .B2(n3708), 
        .ZN(n18572) );
  MOAI22 U27478 ( .A1(n28285), .A2(n3707), .B1(ram[14332]), .B2(n3708), 
        .ZN(n18573) );
  MOAI22 U27479 ( .A1(n28050), .A2(n3707), .B1(ram[14333]), .B2(n3708), 
        .ZN(n18574) );
  MOAI22 U27480 ( .A1(n27815), .A2(n3707), .B1(ram[14334]), .B2(n3708), 
        .ZN(n18575) );
  MOAI22 U27481 ( .A1(n27580), .A2(n3707), .B1(ram[14335]), .B2(n3708), 
        .ZN(n18576) );
  MOAI22 U27482 ( .A1(n29225), .A2(n3709), .B1(ram[14336]), .B2(n3710), 
        .ZN(n18577) );
  MOAI22 U27483 ( .A1(n28990), .A2(n3709), .B1(ram[14337]), .B2(n3710), 
        .ZN(n18578) );
  MOAI22 U27484 ( .A1(n28755), .A2(n3709), .B1(ram[14338]), .B2(n3710), 
        .ZN(n18579) );
  MOAI22 U27485 ( .A1(n28520), .A2(n3709), .B1(ram[14339]), .B2(n3710), 
        .ZN(n18580) );
  MOAI22 U27486 ( .A1(n28285), .A2(n3709), .B1(ram[14340]), .B2(n3710), 
        .ZN(n18581) );
  MOAI22 U27487 ( .A1(n28050), .A2(n3709), .B1(ram[14341]), .B2(n3710), 
        .ZN(n18582) );
  MOAI22 U27488 ( .A1(n27815), .A2(n3709), .B1(ram[14342]), .B2(n3710), 
        .ZN(n18583) );
  MOAI22 U27489 ( .A1(n27580), .A2(n3709), .B1(ram[14343]), .B2(n3710), 
        .ZN(n18584) );
  MOAI22 U27490 ( .A1(n29225), .A2(n3712), .B1(ram[14344]), .B2(n3713), 
        .ZN(n18585) );
  MOAI22 U27491 ( .A1(n28990), .A2(n3712), .B1(ram[14345]), .B2(n3713), 
        .ZN(n18586) );
  MOAI22 U27492 ( .A1(n28755), .A2(n3712), .B1(ram[14346]), .B2(n3713), 
        .ZN(n18587) );
  MOAI22 U27493 ( .A1(n28520), .A2(n3712), .B1(ram[14347]), .B2(n3713), 
        .ZN(n18588) );
  MOAI22 U27494 ( .A1(n28285), .A2(n3712), .B1(ram[14348]), .B2(n3713), 
        .ZN(n18589) );
  MOAI22 U27495 ( .A1(n28050), .A2(n3712), .B1(ram[14349]), .B2(n3713), 
        .ZN(n18590) );
  MOAI22 U27496 ( .A1(n27815), .A2(n3712), .B1(ram[14350]), .B2(n3713), 
        .ZN(n18591) );
  MOAI22 U27497 ( .A1(n27580), .A2(n3712), .B1(ram[14351]), .B2(n3713), 
        .ZN(n18592) );
  MOAI22 U27498 ( .A1(n29226), .A2(n3714), .B1(ram[14352]), .B2(n3715), 
        .ZN(n18593) );
  MOAI22 U27499 ( .A1(n28991), .A2(n3714), .B1(ram[14353]), .B2(n3715), 
        .ZN(n18594) );
  MOAI22 U27500 ( .A1(n28756), .A2(n3714), .B1(ram[14354]), .B2(n3715), 
        .ZN(n18595) );
  MOAI22 U27501 ( .A1(n28521), .A2(n3714), .B1(ram[14355]), .B2(n3715), 
        .ZN(n18596) );
  MOAI22 U27502 ( .A1(n28286), .A2(n3714), .B1(ram[14356]), .B2(n3715), 
        .ZN(n18597) );
  MOAI22 U27503 ( .A1(n28051), .A2(n3714), .B1(ram[14357]), .B2(n3715), 
        .ZN(n18598) );
  MOAI22 U27504 ( .A1(n27816), .A2(n3714), .B1(ram[14358]), .B2(n3715), 
        .ZN(n18599) );
  MOAI22 U27505 ( .A1(n27581), .A2(n3714), .B1(ram[14359]), .B2(n3715), 
        .ZN(n18600) );
  MOAI22 U27506 ( .A1(n29226), .A2(n3716), .B1(ram[14360]), .B2(n3717), 
        .ZN(n18601) );
  MOAI22 U27507 ( .A1(n28991), .A2(n3716), .B1(ram[14361]), .B2(n3717), 
        .ZN(n18602) );
  MOAI22 U27508 ( .A1(n28756), .A2(n3716), .B1(ram[14362]), .B2(n3717), 
        .ZN(n18603) );
  MOAI22 U27509 ( .A1(n28521), .A2(n3716), .B1(ram[14363]), .B2(n3717), 
        .ZN(n18604) );
  MOAI22 U27510 ( .A1(n28286), .A2(n3716), .B1(ram[14364]), .B2(n3717), 
        .ZN(n18605) );
  MOAI22 U27511 ( .A1(n28051), .A2(n3716), .B1(ram[14365]), .B2(n3717), 
        .ZN(n18606) );
  MOAI22 U27512 ( .A1(n27816), .A2(n3716), .B1(ram[14366]), .B2(n3717), 
        .ZN(n18607) );
  MOAI22 U27513 ( .A1(n27581), .A2(n3716), .B1(ram[14367]), .B2(n3717), 
        .ZN(n18608) );
  MOAI22 U27514 ( .A1(n29226), .A2(n3718), .B1(ram[14368]), .B2(n3719), 
        .ZN(n18609) );
  MOAI22 U27515 ( .A1(n28991), .A2(n3718), .B1(ram[14369]), .B2(n3719), 
        .ZN(n18610) );
  MOAI22 U27516 ( .A1(n28756), .A2(n3718), .B1(ram[14370]), .B2(n3719), 
        .ZN(n18611) );
  MOAI22 U27517 ( .A1(n28521), .A2(n3718), .B1(ram[14371]), .B2(n3719), 
        .ZN(n18612) );
  MOAI22 U27518 ( .A1(n28286), .A2(n3718), .B1(ram[14372]), .B2(n3719), 
        .ZN(n18613) );
  MOAI22 U27519 ( .A1(n28051), .A2(n3718), .B1(ram[14373]), .B2(n3719), 
        .ZN(n18614) );
  MOAI22 U27520 ( .A1(n27816), .A2(n3718), .B1(ram[14374]), .B2(n3719), 
        .ZN(n18615) );
  MOAI22 U27521 ( .A1(n27581), .A2(n3718), .B1(ram[14375]), .B2(n3719), 
        .ZN(n18616) );
  MOAI22 U27522 ( .A1(n29226), .A2(n3720), .B1(ram[14376]), .B2(n3721), 
        .ZN(n18617) );
  MOAI22 U27523 ( .A1(n28991), .A2(n3720), .B1(ram[14377]), .B2(n3721), 
        .ZN(n18618) );
  MOAI22 U27524 ( .A1(n28756), .A2(n3720), .B1(ram[14378]), .B2(n3721), 
        .ZN(n18619) );
  MOAI22 U27525 ( .A1(n28521), .A2(n3720), .B1(ram[14379]), .B2(n3721), 
        .ZN(n18620) );
  MOAI22 U27526 ( .A1(n28286), .A2(n3720), .B1(ram[14380]), .B2(n3721), 
        .ZN(n18621) );
  MOAI22 U27527 ( .A1(n28051), .A2(n3720), .B1(ram[14381]), .B2(n3721), 
        .ZN(n18622) );
  MOAI22 U27528 ( .A1(n27816), .A2(n3720), .B1(ram[14382]), .B2(n3721), 
        .ZN(n18623) );
  MOAI22 U27529 ( .A1(n27581), .A2(n3720), .B1(ram[14383]), .B2(n3721), 
        .ZN(n18624) );
  MOAI22 U27530 ( .A1(n29226), .A2(n3722), .B1(ram[14384]), .B2(n3723), 
        .ZN(n18625) );
  MOAI22 U27531 ( .A1(n28991), .A2(n3722), .B1(ram[14385]), .B2(n3723), 
        .ZN(n18626) );
  MOAI22 U27532 ( .A1(n28756), .A2(n3722), .B1(ram[14386]), .B2(n3723), 
        .ZN(n18627) );
  MOAI22 U27533 ( .A1(n28521), .A2(n3722), .B1(ram[14387]), .B2(n3723), 
        .ZN(n18628) );
  MOAI22 U27534 ( .A1(n28286), .A2(n3722), .B1(ram[14388]), .B2(n3723), 
        .ZN(n18629) );
  MOAI22 U27535 ( .A1(n28051), .A2(n3722), .B1(ram[14389]), .B2(n3723), 
        .ZN(n18630) );
  MOAI22 U27536 ( .A1(n27816), .A2(n3722), .B1(ram[14390]), .B2(n3723), 
        .ZN(n18631) );
  MOAI22 U27537 ( .A1(n27581), .A2(n3722), .B1(ram[14391]), .B2(n3723), 
        .ZN(n18632) );
  MOAI22 U27538 ( .A1(n29226), .A2(n3724), .B1(ram[14392]), .B2(n3725), 
        .ZN(n18633) );
  MOAI22 U27539 ( .A1(n28991), .A2(n3724), .B1(ram[14393]), .B2(n3725), 
        .ZN(n18634) );
  MOAI22 U27540 ( .A1(n28756), .A2(n3724), .B1(ram[14394]), .B2(n3725), 
        .ZN(n18635) );
  MOAI22 U27541 ( .A1(n28521), .A2(n3724), .B1(ram[14395]), .B2(n3725), 
        .ZN(n18636) );
  MOAI22 U27542 ( .A1(n28286), .A2(n3724), .B1(ram[14396]), .B2(n3725), 
        .ZN(n18637) );
  MOAI22 U27543 ( .A1(n28051), .A2(n3724), .B1(ram[14397]), .B2(n3725), 
        .ZN(n18638) );
  MOAI22 U27544 ( .A1(n27816), .A2(n3724), .B1(ram[14398]), .B2(n3725), 
        .ZN(n18639) );
  MOAI22 U27545 ( .A1(n27581), .A2(n3724), .B1(ram[14399]), .B2(n3725), 
        .ZN(n18640) );
  MOAI22 U27546 ( .A1(n29226), .A2(n3726), .B1(ram[14400]), .B2(n3727), 
        .ZN(n18641) );
  MOAI22 U27547 ( .A1(n28991), .A2(n3726), .B1(ram[14401]), .B2(n3727), 
        .ZN(n18642) );
  MOAI22 U27548 ( .A1(n28756), .A2(n3726), .B1(ram[14402]), .B2(n3727), 
        .ZN(n18643) );
  MOAI22 U27549 ( .A1(n28521), .A2(n3726), .B1(ram[14403]), .B2(n3727), 
        .ZN(n18644) );
  MOAI22 U27550 ( .A1(n28286), .A2(n3726), .B1(ram[14404]), .B2(n3727), 
        .ZN(n18645) );
  MOAI22 U27551 ( .A1(n28051), .A2(n3726), .B1(ram[14405]), .B2(n3727), 
        .ZN(n18646) );
  MOAI22 U27552 ( .A1(n27816), .A2(n3726), .B1(ram[14406]), .B2(n3727), 
        .ZN(n18647) );
  MOAI22 U27553 ( .A1(n27581), .A2(n3726), .B1(ram[14407]), .B2(n3727), 
        .ZN(n18648) );
  MOAI22 U27554 ( .A1(n29226), .A2(n3728), .B1(ram[14408]), .B2(n3729), 
        .ZN(n18649) );
  MOAI22 U27555 ( .A1(n28991), .A2(n3728), .B1(ram[14409]), .B2(n3729), 
        .ZN(n18650) );
  MOAI22 U27556 ( .A1(n28756), .A2(n3728), .B1(ram[14410]), .B2(n3729), 
        .ZN(n18651) );
  MOAI22 U27557 ( .A1(n28521), .A2(n3728), .B1(ram[14411]), .B2(n3729), 
        .ZN(n18652) );
  MOAI22 U27558 ( .A1(n28286), .A2(n3728), .B1(ram[14412]), .B2(n3729), 
        .ZN(n18653) );
  MOAI22 U27559 ( .A1(n28051), .A2(n3728), .B1(ram[14413]), .B2(n3729), 
        .ZN(n18654) );
  MOAI22 U27560 ( .A1(n27816), .A2(n3728), .B1(ram[14414]), .B2(n3729), 
        .ZN(n18655) );
  MOAI22 U27561 ( .A1(n27581), .A2(n3728), .B1(ram[14415]), .B2(n3729), 
        .ZN(n18656) );
  MOAI22 U27562 ( .A1(n29226), .A2(n3730), .B1(ram[14416]), .B2(n3731), 
        .ZN(n18657) );
  MOAI22 U27563 ( .A1(n28991), .A2(n3730), .B1(ram[14417]), .B2(n3731), 
        .ZN(n18658) );
  MOAI22 U27564 ( .A1(n28756), .A2(n3730), .B1(ram[14418]), .B2(n3731), 
        .ZN(n18659) );
  MOAI22 U27565 ( .A1(n28521), .A2(n3730), .B1(ram[14419]), .B2(n3731), 
        .ZN(n18660) );
  MOAI22 U27566 ( .A1(n28286), .A2(n3730), .B1(ram[14420]), .B2(n3731), 
        .ZN(n18661) );
  MOAI22 U27567 ( .A1(n28051), .A2(n3730), .B1(ram[14421]), .B2(n3731), 
        .ZN(n18662) );
  MOAI22 U27568 ( .A1(n27816), .A2(n3730), .B1(ram[14422]), .B2(n3731), 
        .ZN(n18663) );
  MOAI22 U27569 ( .A1(n27581), .A2(n3730), .B1(ram[14423]), .B2(n3731), 
        .ZN(n18664) );
  MOAI22 U27570 ( .A1(n29226), .A2(n3732), .B1(ram[14424]), .B2(n3733), 
        .ZN(n18665) );
  MOAI22 U27571 ( .A1(n28991), .A2(n3732), .B1(ram[14425]), .B2(n3733), 
        .ZN(n18666) );
  MOAI22 U27572 ( .A1(n28756), .A2(n3732), .B1(ram[14426]), .B2(n3733), 
        .ZN(n18667) );
  MOAI22 U27573 ( .A1(n28521), .A2(n3732), .B1(ram[14427]), .B2(n3733), 
        .ZN(n18668) );
  MOAI22 U27574 ( .A1(n28286), .A2(n3732), .B1(ram[14428]), .B2(n3733), 
        .ZN(n18669) );
  MOAI22 U27575 ( .A1(n28051), .A2(n3732), .B1(ram[14429]), .B2(n3733), 
        .ZN(n18670) );
  MOAI22 U27576 ( .A1(n27816), .A2(n3732), .B1(ram[14430]), .B2(n3733), 
        .ZN(n18671) );
  MOAI22 U27577 ( .A1(n27581), .A2(n3732), .B1(ram[14431]), .B2(n3733), 
        .ZN(n18672) );
  MOAI22 U27578 ( .A1(n29226), .A2(n3734), .B1(ram[14432]), .B2(n3735), 
        .ZN(n18673) );
  MOAI22 U27579 ( .A1(n28991), .A2(n3734), .B1(ram[14433]), .B2(n3735), 
        .ZN(n18674) );
  MOAI22 U27580 ( .A1(n28756), .A2(n3734), .B1(ram[14434]), .B2(n3735), 
        .ZN(n18675) );
  MOAI22 U27581 ( .A1(n28521), .A2(n3734), .B1(ram[14435]), .B2(n3735), 
        .ZN(n18676) );
  MOAI22 U27582 ( .A1(n28286), .A2(n3734), .B1(ram[14436]), .B2(n3735), 
        .ZN(n18677) );
  MOAI22 U27583 ( .A1(n28051), .A2(n3734), .B1(ram[14437]), .B2(n3735), 
        .ZN(n18678) );
  MOAI22 U27584 ( .A1(n27816), .A2(n3734), .B1(ram[14438]), .B2(n3735), 
        .ZN(n18679) );
  MOAI22 U27585 ( .A1(n27581), .A2(n3734), .B1(ram[14439]), .B2(n3735), 
        .ZN(n18680) );
  MOAI22 U27586 ( .A1(n29226), .A2(n3736), .B1(ram[14440]), .B2(n3737), 
        .ZN(n18681) );
  MOAI22 U27587 ( .A1(n28991), .A2(n3736), .B1(ram[14441]), .B2(n3737), 
        .ZN(n18682) );
  MOAI22 U27588 ( .A1(n28756), .A2(n3736), .B1(ram[14442]), .B2(n3737), 
        .ZN(n18683) );
  MOAI22 U27589 ( .A1(n28521), .A2(n3736), .B1(ram[14443]), .B2(n3737), 
        .ZN(n18684) );
  MOAI22 U27590 ( .A1(n28286), .A2(n3736), .B1(ram[14444]), .B2(n3737), 
        .ZN(n18685) );
  MOAI22 U27591 ( .A1(n28051), .A2(n3736), .B1(ram[14445]), .B2(n3737), 
        .ZN(n18686) );
  MOAI22 U27592 ( .A1(n27816), .A2(n3736), .B1(ram[14446]), .B2(n3737), 
        .ZN(n18687) );
  MOAI22 U27593 ( .A1(n27581), .A2(n3736), .B1(ram[14447]), .B2(n3737), 
        .ZN(n18688) );
  MOAI22 U27594 ( .A1(n29226), .A2(n3738), .B1(ram[14448]), .B2(n3739), 
        .ZN(n18689) );
  MOAI22 U27595 ( .A1(n28991), .A2(n3738), .B1(ram[14449]), .B2(n3739), 
        .ZN(n18690) );
  MOAI22 U27596 ( .A1(n28756), .A2(n3738), .B1(ram[14450]), .B2(n3739), 
        .ZN(n18691) );
  MOAI22 U27597 ( .A1(n28521), .A2(n3738), .B1(ram[14451]), .B2(n3739), 
        .ZN(n18692) );
  MOAI22 U27598 ( .A1(n28286), .A2(n3738), .B1(ram[14452]), .B2(n3739), 
        .ZN(n18693) );
  MOAI22 U27599 ( .A1(n28051), .A2(n3738), .B1(ram[14453]), .B2(n3739), 
        .ZN(n18694) );
  MOAI22 U27600 ( .A1(n27816), .A2(n3738), .B1(ram[14454]), .B2(n3739), 
        .ZN(n18695) );
  MOAI22 U27601 ( .A1(n27581), .A2(n3738), .B1(ram[14455]), .B2(n3739), 
        .ZN(n18696) );
  MOAI22 U27602 ( .A1(n29227), .A2(n3740), .B1(ram[14456]), .B2(n3741), 
        .ZN(n18697) );
  MOAI22 U27603 ( .A1(n28992), .A2(n3740), .B1(ram[14457]), .B2(n3741), 
        .ZN(n18698) );
  MOAI22 U27604 ( .A1(n28757), .A2(n3740), .B1(ram[14458]), .B2(n3741), 
        .ZN(n18699) );
  MOAI22 U27605 ( .A1(n28522), .A2(n3740), .B1(ram[14459]), .B2(n3741), 
        .ZN(n18700) );
  MOAI22 U27606 ( .A1(n28287), .A2(n3740), .B1(ram[14460]), .B2(n3741), 
        .ZN(n18701) );
  MOAI22 U27607 ( .A1(n28052), .A2(n3740), .B1(ram[14461]), .B2(n3741), 
        .ZN(n18702) );
  MOAI22 U27608 ( .A1(n27817), .A2(n3740), .B1(ram[14462]), .B2(n3741), 
        .ZN(n18703) );
  MOAI22 U27609 ( .A1(n27582), .A2(n3740), .B1(ram[14463]), .B2(n3741), 
        .ZN(n18704) );
  MOAI22 U27610 ( .A1(n29227), .A2(n3742), .B1(ram[14464]), .B2(n3743), 
        .ZN(n18705) );
  MOAI22 U27611 ( .A1(n28992), .A2(n3742), .B1(ram[14465]), .B2(n3743), 
        .ZN(n18706) );
  MOAI22 U27612 ( .A1(n28757), .A2(n3742), .B1(ram[14466]), .B2(n3743), 
        .ZN(n18707) );
  MOAI22 U27613 ( .A1(n28522), .A2(n3742), .B1(ram[14467]), .B2(n3743), 
        .ZN(n18708) );
  MOAI22 U27614 ( .A1(n28287), .A2(n3742), .B1(ram[14468]), .B2(n3743), 
        .ZN(n18709) );
  MOAI22 U27615 ( .A1(n28052), .A2(n3742), .B1(ram[14469]), .B2(n3743), 
        .ZN(n18710) );
  MOAI22 U27616 ( .A1(n27817), .A2(n3742), .B1(ram[14470]), .B2(n3743), 
        .ZN(n18711) );
  MOAI22 U27617 ( .A1(n27582), .A2(n3742), .B1(ram[14471]), .B2(n3743), 
        .ZN(n18712) );
  MOAI22 U27618 ( .A1(n29227), .A2(n3744), .B1(ram[14472]), .B2(n3745), 
        .ZN(n18713) );
  MOAI22 U27619 ( .A1(n28992), .A2(n3744), .B1(ram[14473]), .B2(n3745), 
        .ZN(n18714) );
  MOAI22 U27620 ( .A1(n28757), .A2(n3744), .B1(ram[14474]), .B2(n3745), 
        .ZN(n18715) );
  MOAI22 U27621 ( .A1(n28522), .A2(n3744), .B1(ram[14475]), .B2(n3745), 
        .ZN(n18716) );
  MOAI22 U27622 ( .A1(n28287), .A2(n3744), .B1(ram[14476]), .B2(n3745), 
        .ZN(n18717) );
  MOAI22 U27623 ( .A1(n28052), .A2(n3744), .B1(ram[14477]), .B2(n3745), 
        .ZN(n18718) );
  MOAI22 U27624 ( .A1(n27817), .A2(n3744), .B1(ram[14478]), .B2(n3745), 
        .ZN(n18719) );
  MOAI22 U27625 ( .A1(n27582), .A2(n3744), .B1(ram[14479]), .B2(n3745), 
        .ZN(n18720) );
  MOAI22 U27626 ( .A1(n29227), .A2(n3746), .B1(ram[14480]), .B2(n3747), 
        .ZN(n18721) );
  MOAI22 U27627 ( .A1(n28992), .A2(n3746), .B1(ram[14481]), .B2(n3747), 
        .ZN(n18722) );
  MOAI22 U27628 ( .A1(n28757), .A2(n3746), .B1(ram[14482]), .B2(n3747), 
        .ZN(n18723) );
  MOAI22 U27629 ( .A1(n28522), .A2(n3746), .B1(ram[14483]), .B2(n3747), 
        .ZN(n18724) );
  MOAI22 U27630 ( .A1(n28287), .A2(n3746), .B1(ram[14484]), .B2(n3747), 
        .ZN(n18725) );
  MOAI22 U27631 ( .A1(n28052), .A2(n3746), .B1(ram[14485]), .B2(n3747), 
        .ZN(n18726) );
  MOAI22 U27632 ( .A1(n27817), .A2(n3746), .B1(ram[14486]), .B2(n3747), 
        .ZN(n18727) );
  MOAI22 U27633 ( .A1(n27582), .A2(n3746), .B1(ram[14487]), .B2(n3747), 
        .ZN(n18728) );
  MOAI22 U27634 ( .A1(n29227), .A2(n3748), .B1(ram[14488]), .B2(n3749), 
        .ZN(n18729) );
  MOAI22 U27635 ( .A1(n28992), .A2(n3748), .B1(ram[14489]), .B2(n3749), 
        .ZN(n18730) );
  MOAI22 U27636 ( .A1(n28757), .A2(n3748), .B1(ram[14490]), .B2(n3749), 
        .ZN(n18731) );
  MOAI22 U27637 ( .A1(n28522), .A2(n3748), .B1(ram[14491]), .B2(n3749), 
        .ZN(n18732) );
  MOAI22 U27638 ( .A1(n28287), .A2(n3748), .B1(ram[14492]), .B2(n3749), 
        .ZN(n18733) );
  MOAI22 U27639 ( .A1(n28052), .A2(n3748), .B1(ram[14493]), .B2(n3749), 
        .ZN(n18734) );
  MOAI22 U27640 ( .A1(n27817), .A2(n3748), .B1(ram[14494]), .B2(n3749), 
        .ZN(n18735) );
  MOAI22 U27641 ( .A1(n27582), .A2(n3748), .B1(ram[14495]), .B2(n3749), 
        .ZN(n18736) );
  MOAI22 U27642 ( .A1(n29227), .A2(n3750), .B1(ram[14496]), .B2(n3751), 
        .ZN(n18737) );
  MOAI22 U27643 ( .A1(n28992), .A2(n3750), .B1(ram[14497]), .B2(n3751), 
        .ZN(n18738) );
  MOAI22 U27644 ( .A1(n28757), .A2(n3750), .B1(ram[14498]), .B2(n3751), 
        .ZN(n18739) );
  MOAI22 U27645 ( .A1(n28522), .A2(n3750), .B1(ram[14499]), .B2(n3751), 
        .ZN(n18740) );
  MOAI22 U27646 ( .A1(n28287), .A2(n3750), .B1(ram[14500]), .B2(n3751), 
        .ZN(n18741) );
  MOAI22 U27647 ( .A1(n28052), .A2(n3750), .B1(ram[14501]), .B2(n3751), 
        .ZN(n18742) );
  MOAI22 U27648 ( .A1(n27817), .A2(n3750), .B1(ram[14502]), .B2(n3751), 
        .ZN(n18743) );
  MOAI22 U27649 ( .A1(n27582), .A2(n3750), .B1(ram[14503]), .B2(n3751), 
        .ZN(n18744) );
  MOAI22 U27650 ( .A1(n29227), .A2(n3752), .B1(ram[14504]), .B2(n3753), 
        .ZN(n18745) );
  MOAI22 U27651 ( .A1(n28992), .A2(n3752), .B1(ram[14505]), .B2(n3753), 
        .ZN(n18746) );
  MOAI22 U27652 ( .A1(n28757), .A2(n3752), .B1(ram[14506]), .B2(n3753), 
        .ZN(n18747) );
  MOAI22 U27653 ( .A1(n28522), .A2(n3752), .B1(ram[14507]), .B2(n3753), 
        .ZN(n18748) );
  MOAI22 U27654 ( .A1(n28287), .A2(n3752), .B1(ram[14508]), .B2(n3753), 
        .ZN(n18749) );
  MOAI22 U27655 ( .A1(n28052), .A2(n3752), .B1(ram[14509]), .B2(n3753), 
        .ZN(n18750) );
  MOAI22 U27656 ( .A1(n27817), .A2(n3752), .B1(ram[14510]), .B2(n3753), 
        .ZN(n18751) );
  MOAI22 U27657 ( .A1(n27582), .A2(n3752), .B1(ram[14511]), .B2(n3753), 
        .ZN(n18752) );
  MOAI22 U27658 ( .A1(n29227), .A2(n3754), .B1(ram[14512]), .B2(n3755), 
        .ZN(n18753) );
  MOAI22 U27659 ( .A1(n28992), .A2(n3754), .B1(ram[14513]), .B2(n3755), 
        .ZN(n18754) );
  MOAI22 U27660 ( .A1(n28757), .A2(n3754), .B1(ram[14514]), .B2(n3755), 
        .ZN(n18755) );
  MOAI22 U27661 ( .A1(n28522), .A2(n3754), .B1(ram[14515]), .B2(n3755), 
        .ZN(n18756) );
  MOAI22 U27662 ( .A1(n28287), .A2(n3754), .B1(ram[14516]), .B2(n3755), 
        .ZN(n18757) );
  MOAI22 U27663 ( .A1(n28052), .A2(n3754), .B1(ram[14517]), .B2(n3755), 
        .ZN(n18758) );
  MOAI22 U27664 ( .A1(n27817), .A2(n3754), .B1(ram[14518]), .B2(n3755), 
        .ZN(n18759) );
  MOAI22 U27665 ( .A1(n27582), .A2(n3754), .B1(ram[14519]), .B2(n3755), 
        .ZN(n18760) );
  MOAI22 U27666 ( .A1(n29227), .A2(n3756), .B1(ram[14520]), .B2(n3757), 
        .ZN(n18761) );
  MOAI22 U27667 ( .A1(n28992), .A2(n3756), .B1(ram[14521]), .B2(n3757), 
        .ZN(n18762) );
  MOAI22 U27668 ( .A1(n28757), .A2(n3756), .B1(ram[14522]), .B2(n3757), 
        .ZN(n18763) );
  MOAI22 U27669 ( .A1(n28522), .A2(n3756), .B1(ram[14523]), .B2(n3757), 
        .ZN(n18764) );
  MOAI22 U27670 ( .A1(n28287), .A2(n3756), .B1(ram[14524]), .B2(n3757), 
        .ZN(n18765) );
  MOAI22 U27671 ( .A1(n28052), .A2(n3756), .B1(ram[14525]), .B2(n3757), 
        .ZN(n18766) );
  MOAI22 U27672 ( .A1(n27817), .A2(n3756), .B1(ram[14526]), .B2(n3757), 
        .ZN(n18767) );
  MOAI22 U27673 ( .A1(n27582), .A2(n3756), .B1(ram[14527]), .B2(n3757), 
        .ZN(n18768) );
  MOAI22 U27674 ( .A1(n29227), .A2(n3758), .B1(ram[14528]), .B2(n3759), 
        .ZN(n18769) );
  MOAI22 U27675 ( .A1(n28992), .A2(n3758), .B1(ram[14529]), .B2(n3759), 
        .ZN(n18770) );
  MOAI22 U27676 ( .A1(n28757), .A2(n3758), .B1(ram[14530]), .B2(n3759), 
        .ZN(n18771) );
  MOAI22 U27677 ( .A1(n28522), .A2(n3758), .B1(ram[14531]), .B2(n3759), 
        .ZN(n18772) );
  MOAI22 U27678 ( .A1(n28287), .A2(n3758), .B1(ram[14532]), .B2(n3759), 
        .ZN(n18773) );
  MOAI22 U27679 ( .A1(n28052), .A2(n3758), .B1(ram[14533]), .B2(n3759), 
        .ZN(n18774) );
  MOAI22 U27680 ( .A1(n27817), .A2(n3758), .B1(ram[14534]), .B2(n3759), 
        .ZN(n18775) );
  MOAI22 U27681 ( .A1(n27582), .A2(n3758), .B1(ram[14535]), .B2(n3759), 
        .ZN(n18776) );
  MOAI22 U27682 ( .A1(n29227), .A2(n3760), .B1(ram[14536]), .B2(n3761), 
        .ZN(n18777) );
  MOAI22 U27683 ( .A1(n28992), .A2(n3760), .B1(ram[14537]), .B2(n3761), 
        .ZN(n18778) );
  MOAI22 U27684 ( .A1(n28757), .A2(n3760), .B1(ram[14538]), .B2(n3761), 
        .ZN(n18779) );
  MOAI22 U27685 ( .A1(n28522), .A2(n3760), .B1(ram[14539]), .B2(n3761), 
        .ZN(n18780) );
  MOAI22 U27686 ( .A1(n28287), .A2(n3760), .B1(ram[14540]), .B2(n3761), 
        .ZN(n18781) );
  MOAI22 U27687 ( .A1(n28052), .A2(n3760), .B1(ram[14541]), .B2(n3761), 
        .ZN(n18782) );
  MOAI22 U27688 ( .A1(n27817), .A2(n3760), .B1(ram[14542]), .B2(n3761), 
        .ZN(n18783) );
  MOAI22 U27689 ( .A1(n27582), .A2(n3760), .B1(ram[14543]), .B2(n3761), 
        .ZN(n18784) );
  MOAI22 U27690 ( .A1(n29227), .A2(n3762), .B1(ram[14544]), .B2(n3763), 
        .ZN(n18785) );
  MOAI22 U27691 ( .A1(n28992), .A2(n3762), .B1(ram[14545]), .B2(n3763), 
        .ZN(n18786) );
  MOAI22 U27692 ( .A1(n28757), .A2(n3762), .B1(ram[14546]), .B2(n3763), 
        .ZN(n18787) );
  MOAI22 U27693 ( .A1(n28522), .A2(n3762), .B1(ram[14547]), .B2(n3763), 
        .ZN(n18788) );
  MOAI22 U27694 ( .A1(n28287), .A2(n3762), .B1(ram[14548]), .B2(n3763), 
        .ZN(n18789) );
  MOAI22 U27695 ( .A1(n28052), .A2(n3762), .B1(ram[14549]), .B2(n3763), 
        .ZN(n18790) );
  MOAI22 U27696 ( .A1(n27817), .A2(n3762), .B1(ram[14550]), .B2(n3763), 
        .ZN(n18791) );
  MOAI22 U27697 ( .A1(n27582), .A2(n3762), .B1(ram[14551]), .B2(n3763), 
        .ZN(n18792) );
  MOAI22 U27698 ( .A1(n29227), .A2(n3764), .B1(ram[14552]), .B2(n3765), 
        .ZN(n18793) );
  MOAI22 U27699 ( .A1(n28992), .A2(n3764), .B1(ram[14553]), .B2(n3765), 
        .ZN(n18794) );
  MOAI22 U27700 ( .A1(n28757), .A2(n3764), .B1(ram[14554]), .B2(n3765), 
        .ZN(n18795) );
  MOAI22 U27701 ( .A1(n28522), .A2(n3764), .B1(ram[14555]), .B2(n3765), 
        .ZN(n18796) );
  MOAI22 U27702 ( .A1(n28287), .A2(n3764), .B1(ram[14556]), .B2(n3765), 
        .ZN(n18797) );
  MOAI22 U27703 ( .A1(n28052), .A2(n3764), .B1(ram[14557]), .B2(n3765), 
        .ZN(n18798) );
  MOAI22 U27704 ( .A1(n27817), .A2(n3764), .B1(ram[14558]), .B2(n3765), 
        .ZN(n18799) );
  MOAI22 U27705 ( .A1(n27582), .A2(n3764), .B1(ram[14559]), .B2(n3765), 
        .ZN(n18800) );
  MOAI22 U27706 ( .A1(n29228), .A2(n3766), .B1(ram[14560]), .B2(n3767), 
        .ZN(n18801) );
  MOAI22 U27707 ( .A1(n28993), .A2(n3766), .B1(ram[14561]), .B2(n3767), 
        .ZN(n18802) );
  MOAI22 U27708 ( .A1(n28758), .A2(n3766), .B1(ram[14562]), .B2(n3767), 
        .ZN(n18803) );
  MOAI22 U27709 ( .A1(n28523), .A2(n3766), .B1(ram[14563]), .B2(n3767), 
        .ZN(n18804) );
  MOAI22 U27710 ( .A1(n28288), .A2(n3766), .B1(ram[14564]), .B2(n3767), 
        .ZN(n18805) );
  MOAI22 U27711 ( .A1(n28053), .A2(n3766), .B1(ram[14565]), .B2(n3767), 
        .ZN(n18806) );
  MOAI22 U27712 ( .A1(n27818), .A2(n3766), .B1(ram[14566]), .B2(n3767), 
        .ZN(n18807) );
  MOAI22 U27713 ( .A1(n27583), .A2(n3766), .B1(ram[14567]), .B2(n3767), 
        .ZN(n18808) );
  MOAI22 U27714 ( .A1(n29228), .A2(n3768), .B1(ram[14568]), .B2(n3769), 
        .ZN(n18809) );
  MOAI22 U27715 ( .A1(n28993), .A2(n3768), .B1(ram[14569]), .B2(n3769), 
        .ZN(n18810) );
  MOAI22 U27716 ( .A1(n28758), .A2(n3768), .B1(ram[14570]), .B2(n3769), 
        .ZN(n18811) );
  MOAI22 U27717 ( .A1(n28523), .A2(n3768), .B1(ram[14571]), .B2(n3769), 
        .ZN(n18812) );
  MOAI22 U27718 ( .A1(n28288), .A2(n3768), .B1(ram[14572]), .B2(n3769), 
        .ZN(n18813) );
  MOAI22 U27719 ( .A1(n28053), .A2(n3768), .B1(ram[14573]), .B2(n3769), 
        .ZN(n18814) );
  MOAI22 U27720 ( .A1(n27818), .A2(n3768), .B1(ram[14574]), .B2(n3769), 
        .ZN(n18815) );
  MOAI22 U27721 ( .A1(n27583), .A2(n3768), .B1(ram[14575]), .B2(n3769), 
        .ZN(n18816) );
  MOAI22 U27722 ( .A1(n29228), .A2(n3770), .B1(ram[14576]), .B2(n3771), 
        .ZN(n18817) );
  MOAI22 U27723 ( .A1(n28993), .A2(n3770), .B1(ram[14577]), .B2(n3771), 
        .ZN(n18818) );
  MOAI22 U27724 ( .A1(n28758), .A2(n3770), .B1(ram[14578]), .B2(n3771), 
        .ZN(n18819) );
  MOAI22 U27725 ( .A1(n28523), .A2(n3770), .B1(ram[14579]), .B2(n3771), 
        .ZN(n18820) );
  MOAI22 U27726 ( .A1(n28288), .A2(n3770), .B1(ram[14580]), .B2(n3771), 
        .ZN(n18821) );
  MOAI22 U27727 ( .A1(n28053), .A2(n3770), .B1(ram[14581]), .B2(n3771), 
        .ZN(n18822) );
  MOAI22 U27728 ( .A1(n27818), .A2(n3770), .B1(ram[14582]), .B2(n3771), 
        .ZN(n18823) );
  MOAI22 U27729 ( .A1(n27583), .A2(n3770), .B1(ram[14583]), .B2(n3771), 
        .ZN(n18824) );
  MOAI22 U27730 ( .A1(n29228), .A2(n3772), .B1(ram[14584]), .B2(n3773), 
        .ZN(n18825) );
  MOAI22 U27731 ( .A1(n28993), .A2(n3772), .B1(ram[14585]), .B2(n3773), 
        .ZN(n18826) );
  MOAI22 U27732 ( .A1(n28758), .A2(n3772), .B1(ram[14586]), .B2(n3773), 
        .ZN(n18827) );
  MOAI22 U27733 ( .A1(n28523), .A2(n3772), .B1(ram[14587]), .B2(n3773), 
        .ZN(n18828) );
  MOAI22 U27734 ( .A1(n28288), .A2(n3772), .B1(ram[14588]), .B2(n3773), 
        .ZN(n18829) );
  MOAI22 U27735 ( .A1(n28053), .A2(n3772), .B1(ram[14589]), .B2(n3773), 
        .ZN(n18830) );
  MOAI22 U27736 ( .A1(n27818), .A2(n3772), .B1(ram[14590]), .B2(n3773), 
        .ZN(n18831) );
  MOAI22 U27737 ( .A1(n27583), .A2(n3772), .B1(ram[14591]), .B2(n3773), 
        .ZN(n18832) );
  MOAI22 U27738 ( .A1(n29228), .A2(n3774), .B1(ram[14592]), .B2(n3775), 
        .ZN(n18833) );
  MOAI22 U27739 ( .A1(n28993), .A2(n3774), .B1(ram[14593]), .B2(n3775), 
        .ZN(n18834) );
  MOAI22 U27740 ( .A1(n28758), .A2(n3774), .B1(ram[14594]), .B2(n3775), 
        .ZN(n18835) );
  MOAI22 U27741 ( .A1(n28523), .A2(n3774), .B1(ram[14595]), .B2(n3775), 
        .ZN(n18836) );
  MOAI22 U27742 ( .A1(n28288), .A2(n3774), .B1(ram[14596]), .B2(n3775), 
        .ZN(n18837) );
  MOAI22 U27743 ( .A1(n28053), .A2(n3774), .B1(ram[14597]), .B2(n3775), 
        .ZN(n18838) );
  MOAI22 U27744 ( .A1(n27818), .A2(n3774), .B1(ram[14598]), .B2(n3775), 
        .ZN(n18839) );
  MOAI22 U27745 ( .A1(n27583), .A2(n3774), .B1(ram[14599]), .B2(n3775), 
        .ZN(n18840) );
  MOAI22 U27746 ( .A1(n29228), .A2(n3776), .B1(ram[14600]), .B2(n3777), 
        .ZN(n18841) );
  MOAI22 U27747 ( .A1(n28993), .A2(n3776), .B1(ram[14601]), .B2(n3777), 
        .ZN(n18842) );
  MOAI22 U27748 ( .A1(n28758), .A2(n3776), .B1(ram[14602]), .B2(n3777), 
        .ZN(n18843) );
  MOAI22 U27749 ( .A1(n28523), .A2(n3776), .B1(ram[14603]), .B2(n3777), 
        .ZN(n18844) );
  MOAI22 U27750 ( .A1(n28288), .A2(n3776), .B1(ram[14604]), .B2(n3777), 
        .ZN(n18845) );
  MOAI22 U27751 ( .A1(n28053), .A2(n3776), .B1(ram[14605]), .B2(n3777), 
        .ZN(n18846) );
  MOAI22 U27752 ( .A1(n27818), .A2(n3776), .B1(ram[14606]), .B2(n3777), 
        .ZN(n18847) );
  MOAI22 U27753 ( .A1(n27583), .A2(n3776), .B1(ram[14607]), .B2(n3777), 
        .ZN(n18848) );
  MOAI22 U27754 ( .A1(n29228), .A2(n3778), .B1(ram[14608]), .B2(n3779), 
        .ZN(n18849) );
  MOAI22 U27755 ( .A1(n28993), .A2(n3778), .B1(ram[14609]), .B2(n3779), 
        .ZN(n18850) );
  MOAI22 U27756 ( .A1(n28758), .A2(n3778), .B1(ram[14610]), .B2(n3779), 
        .ZN(n18851) );
  MOAI22 U27757 ( .A1(n28523), .A2(n3778), .B1(ram[14611]), .B2(n3779), 
        .ZN(n18852) );
  MOAI22 U27758 ( .A1(n28288), .A2(n3778), .B1(ram[14612]), .B2(n3779), 
        .ZN(n18853) );
  MOAI22 U27759 ( .A1(n28053), .A2(n3778), .B1(ram[14613]), .B2(n3779), 
        .ZN(n18854) );
  MOAI22 U27760 ( .A1(n27818), .A2(n3778), .B1(ram[14614]), .B2(n3779), 
        .ZN(n18855) );
  MOAI22 U27761 ( .A1(n27583), .A2(n3778), .B1(ram[14615]), .B2(n3779), 
        .ZN(n18856) );
  MOAI22 U27762 ( .A1(n29228), .A2(n3780), .B1(ram[14616]), .B2(n3781), 
        .ZN(n18857) );
  MOAI22 U27763 ( .A1(n28993), .A2(n3780), .B1(ram[14617]), .B2(n3781), 
        .ZN(n18858) );
  MOAI22 U27764 ( .A1(n28758), .A2(n3780), .B1(ram[14618]), .B2(n3781), 
        .ZN(n18859) );
  MOAI22 U27765 ( .A1(n28523), .A2(n3780), .B1(ram[14619]), .B2(n3781), 
        .ZN(n18860) );
  MOAI22 U27766 ( .A1(n28288), .A2(n3780), .B1(ram[14620]), .B2(n3781), 
        .ZN(n18861) );
  MOAI22 U27767 ( .A1(n28053), .A2(n3780), .B1(ram[14621]), .B2(n3781), 
        .ZN(n18862) );
  MOAI22 U27768 ( .A1(n27818), .A2(n3780), .B1(ram[14622]), .B2(n3781), 
        .ZN(n18863) );
  MOAI22 U27769 ( .A1(n27583), .A2(n3780), .B1(ram[14623]), .B2(n3781), 
        .ZN(n18864) );
  MOAI22 U27770 ( .A1(n29228), .A2(n3782), .B1(ram[14624]), .B2(n3783), 
        .ZN(n18865) );
  MOAI22 U27771 ( .A1(n28993), .A2(n3782), .B1(ram[14625]), .B2(n3783), 
        .ZN(n18866) );
  MOAI22 U27772 ( .A1(n28758), .A2(n3782), .B1(ram[14626]), .B2(n3783), 
        .ZN(n18867) );
  MOAI22 U27773 ( .A1(n28523), .A2(n3782), .B1(ram[14627]), .B2(n3783), 
        .ZN(n18868) );
  MOAI22 U27774 ( .A1(n28288), .A2(n3782), .B1(ram[14628]), .B2(n3783), 
        .ZN(n18869) );
  MOAI22 U27775 ( .A1(n28053), .A2(n3782), .B1(ram[14629]), .B2(n3783), 
        .ZN(n18870) );
  MOAI22 U27776 ( .A1(n27818), .A2(n3782), .B1(ram[14630]), .B2(n3783), 
        .ZN(n18871) );
  MOAI22 U27777 ( .A1(n27583), .A2(n3782), .B1(ram[14631]), .B2(n3783), 
        .ZN(n18872) );
  MOAI22 U27778 ( .A1(n29228), .A2(n3784), .B1(ram[14632]), .B2(n3785), 
        .ZN(n18873) );
  MOAI22 U27779 ( .A1(n28993), .A2(n3784), .B1(ram[14633]), .B2(n3785), 
        .ZN(n18874) );
  MOAI22 U27780 ( .A1(n28758), .A2(n3784), .B1(ram[14634]), .B2(n3785), 
        .ZN(n18875) );
  MOAI22 U27781 ( .A1(n28523), .A2(n3784), .B1(ram[14635]), .B2(n3785), 
        .ZN(n18876) );
  MOAI22 U27782 ( .A1(n28288), .A2(n3784), .B1(ram[14636]), .B2(n3785), 
        .ZN(n18877) );
  MOAI22 U27783 ( .A1(n28053), .A2(n3784), .B1(ram[14637]), .B2(n3785), 
        .ZN(n18878) );
  MOAI22 U27784 ( .A1(n27818), .A2(n3784), .B1(ram[14638]), .B2(n3785), 
        .ZN(n18879) );
  MOAI22 U27785 ( .A1(n27583), .A2(n3784), .B1(ram[14639]), .B2(n3785), 
        .ZN(n18880) );
  MOAI22 U27786 ( .A1(n29228), .A2(n3786), .B1(ram[14640]), .B2(n3787), 
        .ZN(n18881) );
  MOAI22 U27787 ( .A1(n28993), .A2(n3786), .B1(ram[14641]), .B2(n3787), 
        .ZN(n18882) );
  MOAI22 U27788 ( .A1(n28758), .A2(n3786), .B1(ram[14642]), .B2(n3787), 
        .ZN(n18883) );
  MOAI22 U27789 ( .A1(n28523), .A2(n3786), .B1(ram[14643]), .B2(n3787), 
        .ZN(n18884) );
  MOAI22 U27790 ( .A1(n28288), .A2(n3786), .B1(ram[14644]), .B2(n3787), 
        .ZN(n18885) );
  MOAI22 U27791 ( .A1(n28053), .A2(n3786), .B1(ram[14645]), .B2(n3787), 
        .ZN(n18886) );
  MOAI22 U27792 ( .A1(n27818), .A2(n3786), .B1(ram[14646]), .B2(n3787), 
        .ZN(n18887) );
  MOAI22 U27793 ( .A1(n27583), .A2(n3786), .B1(ram[14647]), .B2(n3787), 
        .ZN(n18888) );
  MOAI22 U27794 ( .A1(n29228), .A2(n3788), .B1(ram[14648]), .B2(n3789), 
        .ZN(n18889) );
  MOAI22 U27795 ( .A1(n28993), .A2(n3788), .B1(ram[14649]), .B2(n3789), 
        .ZN(n18890) );
  MOAI22 U27796 ( .A1(n28758), .A2(n3788), .B1(ram[14650]), .B2(n3789), 
        .ZN(n18891) );
  MOAI22 U27797 ( .A1(n28523), .A2(n3788), .B1(ram[14651]), .B2(n3789), 
        .ZN(n18892) );
  MOAI22 U27798 ( .A1(n28288), .A2(n3788), .B1(ram[14652]), .B2(n3789), 
        .ZN(n18893) );
  MOAI22 U27799 ( .A1(n28053), .A2(n3788), .B1(ram[14653]), .B2(n3789), 
        .ZN(n18894) );
  MOAI22 U27800 ( .A1(n27818), .A2(n3788), .B1(ram[14654]), .B2(n3789), 
        .ZN(n18895) );
  MOAI22 U27801 ( .A1(n27583), .A2(n3788), .B1(ram[14655]), .B2(n3789), 
        .ZN(n18896) );
  MOAI22 U27802 ( .A1(n29228), .A2(n3790), .B1(ram[14656]), .B2(n3791), 
        .ZN(n18897) );
  MOAI22 U27803 ( .A1(n28993), .A2(n3790), .B1(ram[14657]), .B2(n3791), 
        .ZN(n18898) );
  MOAI22 U27804 ( .A1(n28758), .A2(n3790), .B1(ram[14658]), .B2(n3791), 
        .ZN(n18899) );
  MOAI22 U27805 ( .A1(n28523), .A2(n3790), .B1(ram[14659]), .B2(n3791), 
        .ZN(n18900) );
  MOAI22 U27806 ( .A1(n28288), .A2(n3790), .B1(ram[14660]), .B2(n3791), 
        .ZN(n18901) );
  MOAI22 U27807 ( .A1(n28053), .A2(n3790), .B1(ram[14661]), .B2(n3791), 
        .ZN(n18902) );
  MOAI22 U27808 ( .A1(n27818), .A2(n3790), .B1(ram[14662]), .B2(n3791), 
        .ZN(n18903) );
  MOAI22 U27809 ( .A1(n27583), .A2(n3790), .B1(ram[14663]), .B2(n3791), 
        .ZN(n18904) );
  MOAI22 U27810 ( .A1(n29229), .A2(n3792), .B1(ram[14664]), .B2(n3793), 
        .ZN(n18905) );
  MOAI22 U27811 ( .A1(n28994), .A2(n3792), .B1(ram[14665]), .B2(n3793), 
        .ZN(n18906) );
  MOAI22 U27812 ( .A1(n28759), .A2(n3792), .B1(ram[14666]), .B2(n3793), 
        .ZN(n18907) );
  MOAI22 U27813 ( .A1(n28524), .A2(n3792), .B1(ram[14667]), .B2(n3793), 
        .ZN(n18908) );
  MOAI22 U27814 ( .A1(n28289), .A2(n3792), .B1(ram[14668]), .B2(n3793), 
        .ZN(n18909) );
  MOAI22 U27815 ( .A1(n28054), .A2(n3792), .B1(ram[14669]), .B2(n3793), 
        .ZN(n18910) );
  MOAI22 U27816 ( .A1(n27819), .A2(n3792), .B1(ram[14670]), .B2(n3793), 
        .ZN(n18911) );
  MOAI22 U27817 ( .A1(n27584), .A2(n3792), .B1(ram[14671]), .B2(n3793), 
        .ZN(n18912) );
  MOAI22 U27818 ( .A1(n29229), .A2(n3794), .B1(ram[14672]), .B2(n3795), 
        .ZN(n18913) );
  MOAI22 U27819 ( .A1(n28994), .A2(n3794), .B1(ram[14673]), .B2(n3795), 
        .ZN(n18914) );
  MOAI22 U27820 ( .A1(n28759), .A2(n3794), .B1(ram[14674]), .B2(n3795), 
        .ZN(n18915) );
  MOAI22 U27821 ( .A1(n28524), .A2(n3794), .B1(ram[14675]), .B2(n3795), 
        .ZN(n18916) );
  MOAI22 U27822 ( .A1(n28289), .A2(n3794), .B1(ram[14676]), .B2(n3795), 
        .ZN(n18917) );
  MOAI22 U27823 ( .A1(n28054), .A2(n3794), .B1(ram[14677]), .B2(n3795), 
        .ZN(n18918) );
  MOAI22 U27824 ( .A1(n27819), .A2(n3794), .B1(ram[14678]), .B2(n3795), 
        .ZN(n18919) );
  MOAI22 U27825 ( .A1(n27584), .A2(n3794), .B1(ram[14679]), .B2(n3795), 
        .ZN(n18920) );
  MOAI22 U27826 ( .A1(n29229), .A2(n3796), .B1(ram[14680]), .B2(n3797), 
        .ZN(n18921) );
  MOAI22 U27827 ( .A1(n28994), .A2(n3796), .B1(ram[14681]), .B2(n3797), 
        .ZN(n18922) );
  MOAI22 U27828 ( .A1(n28759), .A2(n3796), .B1(ram[14682]), .B2(n3797), 
        .ZN(n18923) );
  MOAI22 U27829 ( .A1(n28524), .A2(n3796), .B1(ram[14683]), .B2(n3797), 
        .ZN(n18924) );
  MOAI22 U27830 ( .A1(n28289), .A2(n3796), .B1(ram[14684]), .B2(n3797), 
        .ZN(n18925) );
  MOAI22 U27831 ( .A1(n28054), .A2(n3796), .B1(ram[14685]), .B2(n3797), 
        .ZN(n18926) );
  MOAI22 U27832 ( .A1(n27819), .A2(n3796), .B1(ram[14686]), .B2(n3797), 
        .ZN(n18927) );
  MOAI22 U27833 ( .A1(n27584), .A2(n3796), .B1(ram[14687]), .B2(n3797), 
        .ZN(n18928) );
  MOAI22 U27834 ( .A1(n29229), .A2(n3798), .B1(ram[14688]), .B2(n3799), 
        .ZN(n18929) );
  MOAI22 U27835 ( .A1(n28994), .A2(n3798), .B1(ram[14689]), .B2(n3799), 
        .ZN(n18930) );
  MOAI22 U27836 ( .A1(n28759), .A2(n3798), .B1(ram[14690]), .B2(n3799), 
        .ZN(n18931) );
  MOAI22 U27837 ( .A1(n28524), .A2(n3798), .B1(ram[14691]), .B2(n3799), 
        .ZN(n18932) );
  MOAI22 U27838 ( .A1(n28289), .A2(n3798), .B1(ram[14692]), .B2(n3799), 
        .ZN(n18933) );
  MOAI22 U27839 ( .A1(n28054), .A2(n3798), .B1(ram[14693]), .B2(n3799), 
        .ZN(n18934) );
  MOAI22 U27840 ( .A1(n27819), .A2(n3798), .B1(ram[14694]), .B2(n3799), 
        .ZN(n18935) );
  MOAI22 U27841 ( .A1(n27584), .A2(n3798), .B1(ram[14695]), .B2(n3799), 
        .ZN(n18936) );
  MOAI22 U27842 ( .A1(n29229), .A2(n3800), .B1(ram[14696]), .B2(n3801), 
        .ZN(n18937) );
  MOAI22 U27843 ( .A1(n28994), .A2(n3800), .B1(ram[14697]), .B2(n3801), 
        .ZN(n18938) );
  MOAI22 U27844 ( .A1(n28759), .A2(n3800), .B1(ram[14698]), .B2(n3801), 
        .ZN(n18939) );
  MOAI22 U27845 ( .A1(n28524), .A2(n3800), .B1(ram[14699]), .B2(n3801), 
        .ZN(n18940) );
  MOAI22 U27846 ( .A1(n28289), .A2(n3800), .B1(ram[14700]), .B2(n3801), 
        .ZN(n18941) );
  MOAI22 U27847 ( .A1(n28054), .A2(n3800), .B1(ram[14701]), .B2(n3801), 
        .ZN(n18942) );
  MOAI22 U27848 ( .A1(n27819), .A2(n3800), .B1(ram[14702]), .B2(n3801), 
        .ZN(n18943) );
  MOAI22 U27849 ( .A1(n27584), .A2(n3800), .B1(ram[14703]), .B2(n3801), 
        .ZN(n18944) );
  MOAI22 U27850 ( .A1(n29229), .A2(n3802), .B1(ram[14704]), .B2(n3803), 
        .ZN(n18945) );
  MOAI22 U27851 ( .A1(n28994), .A2(n3802), .B1(ram[14705]), .B2(n3803), 
        .ZN(n18946) );
  MOAI22 U27852 ( .A1(n28759), .A2(n3802), .B1(ram[14706]), .B2(n3803), 
        .ZN(n18947) );
  MOAI22 U27853 ( .A1(n28524), .A2(n3802), .B1(ram[14707]), .B2(n3803), 
        .ZN(n18948) );
  MOAI22 U27854 ( .A1(n28289), .A2(n3802), .B1(ram[14708]), .B2(n3803), 
        .ZN(n18949) );
  MOAI22 U27855 ( .A1(n28054), .A2(n3802), .B1(ram[14709]), .B2(n3803), 
        .ZN(n18950) );
  MOAI22 U27856 ( .A1(n27819), .A2(n3802), .B1(ram[14710]), .B2(n3803), 
        .ZN(n18951) );
  MOAI22 U27857 ( .A1(n27584), .A2(n3802), .B1(ram[14711]), .B2(n3803), 
        .ZN(n18952) );
  MOAI22 U27858 ( .A1(n29229), .A2(n3804), .B1(ram[14712]), .B2(n3805), 
        .ZN(n18953) );
  MOAI22 U27859 ( .A1(n28994), .A2(n3804), .B1(ram[14713]), .B2(n3805), 
        .ZN(n18954) );
  MOAI22 U27860 ( .A1(n28759), .A2(n3804), .B1(ram[14714]), .B2(n3805), 
        .ZN(n18955) );
  MOAI22 U27861 ( .A1(n28524), .A2(n3804), .B1(ram[14715]), .B2(n3805), 
        .ZN(n18956) );
  MOAI22 U27862 ( .A1(n28289), .A2(n3804), .B1(ram[14716]), .B2(n3805), 
        .ZN(n18957) );
  MOAI22 U27863 ( .A1(n28054), .A2(n3804), .B1(ram[14717]), .B2(n3805), 
        .ZN(n18958) );
  MOAI22 U27864 ( .A1(n27819), .A2(n3804), .B1(ram[14718]), .B2(n3805), 
        .ZN(n18959) );
  MOAI22 U27865 ( .A1(n27584), .A2(n3804), .B1(ram[14719]), .B2(n3805), 
        .ZN(n18960) );
  MOAI22 U27866 ( .A1(n29229), .A2(n3806), .B1(ram[14720]), .B2(n3807), 
        .ZN(n18961) );
  MOAI22 U27867 ( .A1(n28994), .A2(n3806), .B1(ram[14721]), .B2(n3807), 
        .ZN(n18962) );
  MOAI22 U27868 ( .A1(n28759), .A2(n3806), .B1(ram[14722]), .B2(n3807), 
        .ZN(n18963) );
  MOAI22 U27869 ( .A1(n28524), .A2(n3806), .B1(ram[14723]), .B2(n3807), 
        .ZN(n18964) );
  MOAI22 U27870 ( .A1(n28289), .A2(n3806), .B1(ram[14724]), .B2(n3807), 
        .ZN(n18965) );
  MOAI22 U27871 ( .A1(n28054), .A2(n3806), .B1(ram[14725]), .B2(n3807), 
        .ZN(n18966) );
  MOAI22 U27872 ( .A1(n27819), .A2(n3806), .B1(ram[14726]), .B2(n3807), 
        .ZN(n18967) );
  MOAI22 U27873 ( .A1(n27584), .A2(n3806), .B1(ram[14727]), .B2(n3807), 
        .ZN(n18968) );
  MOAI22 U27874 ( .A1(n29229), .A2(n3808), .B1(ram[14728]), .B2(n3809), 
        .ZN(n18969) );
  MOAI22 U27875 ( .A1(n28994), .A2(n3808), .B1(ram[14729]), .B2(n3809), 
        .ZN(n18970) );
  MOAI22 U27876 ( .A1(n28759), .A2(n3808), .B1(ram[14730]), .B2(n3809), 
        .ZN(n18971) );
  MOAI22 U27877 ( .A1(n28524), .A2(n3808), .B1(ram[14731]), .B2(n3809), 
        .ZN(n18972) );
  MOAI22 U27878 ( .A1(n28289), .A2(n3808), .B1(ram[14732]), .B2(n3809), 
        .ZN(n18973) );
  MOAI22 U27879 ( .A1(n28054), .A2(n3808), .B1(ram[14733]), .B2(n3809), 
        .ZN(n18974) );
  MOAI22 U27880 ( .A1(n27819), .A2(n3808), .B1(ram[14734]), .B2(n3809), 
        .ZN(n18975) );
  MOAI22 U27881 ( .A1(n27584), .A2(n3808), .B1(ram[14735]), .B2(n3809), 
        .ZN(n18976) );
  MOAI22 U27882 ( .A1(n29229), .A2(n3810), .B1(ram[14736]), .B2(n3811), 
        .ZN(n18977) );
  MOAI22 U27883 ( .A1(n28994), .A2(n3810), .B1(ram[14737]), .B2(n3811), 
        .ZN(n18978) );
  MOAI22 U27884 ( .A1(n28759), .A2(n3810), .B1(ram[14738]), .B2(n3811), 
        .ZN(n18979) );
  MOAI22 U27885 ( .A1(n28524), .A2(n3810), .B1(ram[14739]), .B2(n3811), 
        .ZN(n18980) );
  MOAI22 U27886 ( .A1(n28289), .A2(n3810), .B1(ram[14740]), .B2(n3811), 
        .ZN(n18981) );
  MOAI22 U27887 ( .A1(n28054), .A2(n3810), .B1(ram[14741]), .B2(n3811), 
        .ZN(n18982) );
  MOAI22 U27888 ( .A1(n27819), .A2(n3810), .B1(ram[14742]), .B2(n3811), 
        .ZN(n18983) );
  MOAI22 U27889 ( .A1(n27584), .A2(n3810), .B1(ram[14743]), .B2(n3811), 
        .ZN(n18984) );
  MOAI22 U27890 ( .A1(n29229), .A2(n3812), .B1(ram[14744]), .B2(n3813), 
        .ZN(n18985) );
  MOAI22 U27891 ( .A1(n28994), .A2(n3812), .B1(ram[14745]), .B2(n3813), 
        .ZN(n18986) );
  MOAI22 U27892 ( .A1(n28759), .A2(n3812), .B1(ram[14746]), .B2(n3813), 
        .ZN(n18987) );
  MOAI22 U27893 ( .A1(n28524), .A2(n3812), .B1(ram[14747]), .B2(n3813), 
        .ZN(n18988) );
  MOAI22 U27894 ( .A1(n28289), .A2(n3812), .B1(ram[14748]), .B2(n3813), 
        .ZN(n18989) );
  MOAI22 U27895 ( .A1(n28054), .A2(n3812), .B1(ram[14749]), .B2(n3813), 
        .ZN(n18990) );
  MOAI22 U27896 ( .A1(n27819), .A2(n3812), .B1(ram[14750]), .B2(n3813), 
        .ZN(n18991) );
  MOAI22 U27897 ( .A1(n27584), .A2(n3812), .B1(ram[14751]), .B2(n3813), 
        .ZN(n18992) );
  MOAI22 U27898 ( .A1(n29229), .A2(n3814), .B1(ram[14752]), .B2(n3815), 
        .ZN(n18993) );
  MOAI22 U27899 ( .A1(n28994), .A2(n3814), .B1(ram[14753]), .B2(n3815), 
        .ZN(n18994) );
  MOAI22 U27900 ( .A1(n28759), .A2(n3814), .B1(ram[14754]), .B2(n3815), 
        .ZN(n18995) );
  MOAI22 U27901 ( .A1(n28524), .A2(n3814), .B1(ram[14755]), .B2(n3815), 
        .ZN(n18996) );
  MOAI22 U27902 ( .A1(n28289), .A2(n3814), .B1(ram[14756]), .B2(n3815), 
        .ZN(n18997) );
  MOAI22 U27903 ( .A1(n28054), .A2(n3814), .B1(ram[14757]), .B2(n3815), 
        .ZN(n18998) );
  MOAI22 U27904 ( .A1(n27819), .A2(n3814), .B1(ram[14758]), .B2(n3815), 
        .ZN(n18999) );
  MOAI22 U27905 ( .A1(n27584), .A2(n3814), .B1(ram[14759]), .B2(n3815), 
        .ZN(n19000) );
  MOAI22 U27906 ( .A1(n29229), .A2(n3816), .B1(ram[14760]), .B2(n3817), 
        .ZN(n19001) );
  MOAI22 U27907 ( .A1(n28994), .A2(n3816), .B1(ram[14761]), .B2(n3817), 
        .ZN(n19002) );
  MOAI22 U27908 ( .A1(n28759), .A2(n3816), .B1(ram[14762]), .B2(n3817), 
        .ZN(n19003) );
  MOAI22 U27909 ( .A1(n28524), .A2(n3816), .B1(ram[14763]), .B2(n3817), 
        .ZN(n19004) );
  MOAI22 U27910 ( .A1(n28289), .A2(n3816), .B1(ram[14764]), .B2(n3817), 
        .ZN(n19005) );
  MOAI22 U27911 ( .A1(n28054), .A2(n3816), .B1(ram[14765]), .B2(n3817), 
        .ZN(n19006) );
  MOAI22 U27912 ( .A1(n27819), .A2(n3816), .B1(ram[14766]), .B2(n3817), 
        .ZN(n19007) );
  MOAI22 U27913 ( .A1(n27584), .A2(n3816), .B1(ram[14767]), .B2(n3817), 
        .ZN(n19008) );
  MOAI22 U27914 ( .A1(n29230), .A2(n3818), .B1(ram[14768]), .B2(n3819), 
        .ZN(n19009) );
  MOAI22 U27915 ( .A1(n28995), .A2(n3818), .B1(ram[14769]), .B2(n3819), 
        .ZN(n19010) );
  MOAI22 U27916 ( .A1(n28760), .A2(n3818), .B1(ram[14770]), .B2(n3819), 
        .ZN(n19011) );
  MOAI22 U27917 ( .A1(n28525), .A2(n3818), .B1(ram[14771]), .B2(n3819), 
        .ZN(n19012) );
  MOAI22 U27918 ( .A1(n28290), .A2(n3818), .B1(ram[14772]), .B2(n3819), 
        .ZN(n19013) );
  MOAI22 U27919 ( .A1(n28055), .A2(n3818), .B1(ram[14773]), .B2(n3819), 
        .ZN(n19014) );
  MOAI22 U27920 ( .A1(n27820), .A2(n3818), .B1(ram[14774]), .B2(n3819), 
        .ZN(n19015) );
  MOAI22 U27921 ( .A1(n27585), .A2(n3818), .B1(ram[14775]), .B2(n3819), 
        .ZN(n19016) );
  MOAI22 U27922 ( .A1(n29230), .A2(n3820), .B1(ram[14776]), .B2(n3821), 
        .ZN(n19017) );
  MOAI22 U27923 ( .A1(n28995), .A2(n3820), .B1(ram[14777]), .B2(n3821), 
        .ZN(n19018) );
  MOAI22 U27924 ( .A1(n28760), .A2(n3820), .B1(ram[14778]), .B2(n3821), 
        .ZN(n19019) );
  MOAI22 U27925 ( .A1(n28525), .A2(n3820), .B1(ram[14779]), .B2(n3821), 
        .ZN(n19020) );
  MOAI22 U27926 ( .A1(n28290), .A2(n3820), .B1(ram[14780]), .B2(n3821), 
        .ZN(n19021) );
  MOAI22 U27927 ( .A1(n28055), .A2(n3820), .B1(ram[14781]), .B2(n3821), 
        .ZN(n19022) );
  MOAI22 U27928 ( .A1(n27820), .A2(n3820), .B1(ram[14782]), .B2(n3821), 
        .ZN(n19023) );
  MOAI22 U27929 ( .A1(n27585), .A2(n3820), .B1(ram[14783]), .B2(n3821), 
        .ZN(n19024) );
  MOAI22 U27930 ( .A1(n29230), .A2(n3822), .B1(ram[14784]), .B2(n3823), 
        .ZN(n19025) );
  MOAI22 U27931 ( .A1(n28995), .A2(n3822), .B1(ram[14785]), .B2(n3823), 
        .ZN(n19026) );
  MOAI22 U27932 ( .A1(n28760), .A2(n3822), .B1(ram[14786]), .B2(n3823), 
        .ZN(n19027) );
  MOAI22 U27933 ( .A1(n28525), .A2(n3822), .B1(ram[14787]), .B2(n3823), 
        .ZN(n19028) );
  MOAI22 U27934 ( .A1(n28290), .A2(n3822), .B1(ram[14788]), .B2(n3823), 
        .ZN(n19029) );
  MOAI22 U27935 ( .A1(n28055), .A2(n3822), .B1(ram[14789]), .B2(n3823), 
        .ZN(n19030) );
  MOAI22 U27936 ( .A1(n27820), .A2(n3822), .B1(ram[14790]), .B2(n3823), 
        .ZN(n19031) );
  MOAI22 U27937 ( .A1(n27585), .A2(n3822), .B1(ram[14791]), .B2(n3823), 
        .ZN(n19032) );
  MOAI22 U27938 ( .A1(n29230), .A2(n3824), .B1(ram[14792]), .B2(n3825), 
        .ZN(n19033) );
  MOAI22 U27939 ( .A1(n28995), .A2(n3824), .B1(ram[14793]), .B2(n3825), 
        .ZN(n19034) );
  MOAI22 U27940 ( .A1(n28760), .A2(n3824), .B1(ram[14794]), .B2(n3825), 
        .ZN(n19035) );
  MOAI22 U27941 ( .A1(n28525), .A2(n3824), .B1(ram[14795]), .B2(n3825), 
        .ZN(n19036) );
  MOAI22 U27942 ( .A1(n28290), .A2(n3824), .B1(ram[14796]), .B2(n3825), 
        .ZN(n19037) );
  MOAI22 U27943 ( .A1(n28055), .A2(n3824), .B1(ram[14797]), .B2(n3825), 
        .ZN(n19038) );
  MOAI22 U27944 ( .A1(n27820), .A2(n3824), .B1(ram[14798]), .B2(n3825), 
        .ZN(n19039) );
  MOAI22 U27945 ( .A1(n27585), .A2(n3824), .B1(ram[14799]), .B2(n3825), 
        .ZN(n19040) );
  MOAI22 U27946 ( .A1(n29230), .A2(n3826), .B1(ram[14800]), .B2(n3827), 
        .ZN(n19041) );
  MOAI22 U27947 ( .A1(n28995), .A2(n3826), .B1(ram[14801]), .B2(n3827), 
        .ZN(n19042) );
  MOAI22 U27948 ( .A1(n28760), .A2(n3826), .B1(ram[14802]), .B2(n3827), 
        .ZN(n19043) );
  MOAI22 U27949 ( .A1(n28525), .A2(n3826), .B1(ram[14803]), .B2(n3827), 
        .ZN(n19044) );
  MOAI22 U27950 ( .A1(n28290), .A2(n3826), .B1(ram[14804]), .B2(n3827), 
        .ZN(n19045) );
  MOAI22 U27951 ( .A1(n28055), .A2(n3826), .B1(ram[14805]), .B2(n3827), 
        .ZN(n19046) );
  MOAI22 U27952 ( .A1(n27820), .A2(n3826), .B1(ram[14806]), .B2(n3827), 
        .ZN(n19047) );
  MOAI22 U27953 ( .A1(n27585), .A2(n3826), .B1(ram[14807]), .B2(n3827), 
        .ZN(n19048) );
  MOAI22 U27954 ( .A1(n29230), .A2(n3828), .B1(ram[14808]), .B2(n3829), 
        .ZN(n19049) );
  MOAI22 U27955 ( .A1(n28995), .A2(n3828), .B1(ram[14809]), .B2(n3829), 
        .ZN(n19050) );
  MOAI22 U27956 ( .A1(n28760), .A2(n3828), .B1(ram[14810]), .B2(n3829), 
        .ZN(n19051) );
  MOAI22 U27957 ( .A1(n28525), .A2(n3828), .B1(ram[14811]), .B2(n3829), 
        .ZN(n19052) );
  MOAI22 U27958 ( .A1(n28290), .A2(n3828), .B1(ram[14812]), .B2(n3829), 
        .ZN(n19053) );
  MOAI22 U27959 ( .A1(n28055), .A2(n3828), .B1(ram[14813]), .B2(n3829), 
        .ZN(n19054) );
  MOAI22 U27960 ( .A1(n27820), .A2(n3828), .B1(ram[14814]), .B2(n3829), 
        .ZN(n19055) );
  MOAI22 U27961 ( .A1(n27585), .A2(n3828), .B1(ram[14815]), .B2(n3829), 
        .ZN(n19056) );
  MOAI22 U27962 ( .A1(n29230), .A2(n3830), .B1(ram[14816]), .B2(n3831), 
        .ZN(n19057) );
  MOAI22 U27963 ( .A1(n28995), .A2(n3830), .B1(ram[14817]), .B2(n3831), 
        .ZN(n19058) );
  MOAI22 U27964 ( .A1(n28760), .A2(n3830), .B1(ram[14818]), .B2(n3831), 
        .ZN(n19059) );
  MOAI22 U27965 ( .A1(n28525), .A2(n3830), .B1(ram[14819]), .B2(n3831), 
        .ZN(n19060) );
  MOAI22 U27966 ( .A1(n28290), .A2(n3830), .B1(ram[14820]), .B2(n3831), 
        .ZN(n19061) );
  MOAI22 U27967 ( .A1(n28055), .A2(n3830), .B1(ram[14821]), .B2(n3831), 
        .ZN(n19062) );
  MOAI22 U27968 ( .A1(n27820), .A2(n3830), .B1(ram[14822]), .B2(n3831), 
        .ZN(n19063) );
  MOAI22 U27969 ( .A1(n27585), .A2(n3830), .B1(ram[14823]), .B2(n3831), 
        .ZN(n19064) );
  MOAI22 U27970 ( .A1(n29230), .A2(n3832), .B1(ram[14824]), .B2(n3833), 
        .ZN(n19065) );
  MOAI22 U27971 ( .A1(n28995), .A2(n3832), .B1(ram[14825]), .B2(n3833), 
        .ZN(n19066) );
  MOAI22 U27972 ( .A1(n28760), .A2(n3832), .B1(ram[14826]), .B2(n3833), 
        .ZN(n19067) );
  MOAI22 U27973 ( .A1(n28525), .A2(n3832), .B1(ram[14827]), .B2(n3833), 
        .ZN(n19068) );
  MOAI22 U27974 ( .A1(n28290), .A2(n3832), .B1(ram[14828]), .B2(n3833), 
        .ZN(n19069) );
  MOAI22 U27975 ( .A1(n28055), .A2(n3832), .B1(ram[14829]), .B2(n3833), 
        .ZN(n19070) );
  MOAI22 U27976 ( .A1(n27820), .A2(n3832), .B1(ram[14830]), .B2(n3833), 
        .ZN(n19071) );
  MOAI22 U27977 ( .A1(n27585), .A2(n3832), .B1(ram[14831]), .B2(n3833), 
        .ZN(n19072) );
  MOAI22 U27978 ( .A1(n29230), .A2(n3834), .B1(ram[14832]), .B2(n3835), 
        .ZN(n19073) );
  MOAI22 U27979 ( .A1(n28995), .A2(n3834), .B1(ram[14833]), .B2(n3835), 
        .ZN(n19074) );
  MOAI22 U27980 ( .A1(n28760), .A2(n3834), .B1(ram[14834]), .B2(n3835), 
        .ZN(n19075) );
  MOAI22 U27981 ( .A1(n28525), .A2(n3834), .B1(ram[14835]), .B2(n3835), 
        .ZN(n19076) );
  MOAI22 U27982 ( .A1(n28290), .A2(n3834), .B1(ram[14836]), .B2(n3835), 
        .ZN(n19077) );
  MOAI22 U27983 ( .A1(n28055), .A2(n3834), .B1(ram[14837]), .B2(n3835), 
        .ZN(n19078) );
  MOAI22 U27984 ( .A1(n27820), .A2(n3834), .B1(ram[14838]), .B2(n3835), 
        .ZN(n19079) );
  MOAI22 U27985 ( .A1(n27585), .A2(n3834), .B1(ram[14839]), .B2(n3835), 
        .ZN(n19080) );
  MOAI22 U27986 ( .A1(n29230), .A2(n3836), .B1(ram[14840]), .B2(n3837), 
        .ZN(n19081) );
  MOAI22 U27987 ( .A1(n28995), .A2(n3836), .B1(ram[14841]), .B2(n3837), 
        .ZN(n19082) );
  MOAI22 U27988 ( .A1(n28760), .A2(n3836), .B1(ram[14842]), .B2(n3837), 
        .ZN(n19083) );
  MOAI22 U27989 ( .A1(n28525), .A2(n3836), .B1(ram[14843]), .B2(n3837), 
        .ZN(n19084) );
  MOAI22 U27990 ( .A1(n28290), .A2(n3836), .B1(ram[14844]), .B2(n3837), 
        .ZN(n19085) );
  MOAI22 U27991 ( .A1(n28055), .A2(n3836), .B1(ram[14845]), .B2(n3837), 
        .ZN(n19086) );
  MOAI22 U27992 ( .A1(n27820), .A2(n3836), .B1(ram[14846]), .B2(n3837), 
        .ZN(n19087) );
  MOAI22 U27993 ( .A1(n27585), .A2(n3836), .B1(ram[14847]), .B2(n3837), 
        .ZN(n19088) );
  MOAI22 U27994 ( .A1(n29230), .A2(n3838), .B1(ram[14848]), .B2(n3839), 
        .ZN(n19089) );
  MOAI22 U27995 ( .A1(n28995), .A2(n3838), .B1(ram[14849]), .B2(n3839), 
        .ZN(n19090) );
  MOAI22 U27996 ( .A1(n28760), .A2(n3838), .B1(ram[14850]), .B2(n3839), 
        .ZN(n19091) );
  MOAI22 U27997 ( .A1(n28525), .A2(n3838), .B1(ram[14851]), .B2(n3839), 
        .ZN(n19092) );
  MOAI22 U27998 ( .A1(n28290), .A2(n3838), .B1(ram[14852]), .B2(n3839), 
        .ZN(n19093) );
  MOAI22 U27999 ( .A1(n28055), .A2(n3838), .B1(ram[14853]), .B2(n3839), 
        .ZN(n19094) );
  MOAI22 U28000 ( .A1(n27820), .A2(n3838), .B1(ram[14854]), .B2(n3839), 
        .ZN(n19095) );
  MOAI22 U28001 ( .A1(n27585), .A2(n3838), .B1(ram[14855]), .B2(n3839), 
        .ZN(n19096) );
  MOAI22 U28002 ( .A1(n29230), .A2(n3841), .B1(ram[14856]), .B2(n3842), 
        .ZN(n19097) );
  MOAI22 U28003 ( .A1(n28995), .A2(n3841), .B1(ram[14857]), .B2(n3842), 
        .ZN(n19098) );
  MOAI22 U28004 ( .A1(n28760), .A2(n3841), .B1(ram[14858]), .B2(n3842), 
        .ZN(n19099) );
  MOAI22 U28005 ( .A1(n28525), .A2(n3841), .B1(ram[14859]), .B2(n3842), 
        .ZN(n19100) );
  MOAI22 U28006 ( .A1(n28290), .A2(n3841), .B1(ram[14860]), .B2(n3842), 
        .ZN(n19101) );
  MOAI22 U28007 ( .A1(n28055), .A2(n3841), .B1(ram[14861]), .B2(n3842), 
        .ZN(n19102) );
  MOAI22 U28008 ( .A1(n27820), .A2(n3841), .B1(ram[14862]), .B2(n3842), 
        .ZN(n19103) );
  MOAI22 U28009 ( .A1(n27585), .A2(n3841), .B1(ram[14863]), .B2(n3842), 
        .ZN(n19104) );
  MOAI22 U28010 ( .A1(n29230), .A2(n3843), .B1(ram[14864]), .B2(n3844), 
        .ZN(n19105) );
  MOAI22 U28011 ( .A1(n28995), .A2(n3843), .B1(ram[14865]), .B2(n3844), 
        .ZN(n19106) );
  MOAI22 U28012 ( .A1(n28760), .A2(n3843), .B1(ram[14866]), .B2(n3844), 
        .ZN(n19107) );
  MOAI22 U28013 ( .A1(n28525), .A2(n3843), .B1(ram[14867]), .B2(n3844), 
        .ZN(n19108) );
  MOAI22 U28014 ( .A1(n28290), .A2(n3843), .B1(ram[14868]), .B2(n3844), 
        .ZN(n19109) );
  MOAI22 U28015 ( .A1(n28055), .A2(n3843), .B1(ram[14869]), .B2(n3844), 
        .ZN(n19110) );
  MOAI22 U28016 ( .A1(n27820), .A2(n3843), .B1(ram[14870]), .B2(n3844), 
        .ZN(n19111) );
  MOAI22 U28017 ( .A1(n27585), .A2(n3843), .B1(ram[14871]), .B2(n3844), 
        .ZN(n19112) );
  MOAI22 U28018 ( .A1(n29231), .A2(n3845), .B1(ram[14872]), .B2(n3846), 
        .ZN(n19113) );
  MOAI22 U28019 ( .A1(n28996), .A2(n3845), .B1(ram[14873]), .B2(n3846), 
        .ZN(n19114) );
  MOAI22 U28020 ( .A1(n28761), .A2(n3845), .B1(ram[14874]), .B2(n3846), 
        .ZN(n19115) );
  MOAI22 U28021 ( .A1(n28526), .A2(n3845), .B1(ram[14875]), .B2(n3846), 
        .ZN(n19116) );
  MOAI22 U28022 ( .A1(n28291), .A2(n3845), .B1(ram[14876]), .B2(n3846), 
        .ZN(n19117) );
  MOAI22 U28023 ( .A1(n28056), .A2(n3845), .B1(ram[14877]), .B2(n3846), 
        .ZN(n19118) );
  MOAI22 U28024 ( .A1(n27821), .A2(n3845), .B1(ram[14878]), .B2(n3846), 
        .ZN(n19119) );
  MOAI22 U28025 ( .A1(n27586), .A2(n3845), .B1(ram[14879]), .B2(n3846), 
        .ZN(n19120) );
  MOAI22 U28026 ( .A1(n29231), .A2(n3847), .B1(ram[14880]), .B2(n3848), 
        .ZN(n19121) );
  MOAI22 U28027 ( .A1(n28996), .A2(n3847), .B1(ram[14881]), .B2(n3848), 
        .ZN(n19122) );
  MOAI22 U28028 ( .A1(n28761), .A2(n3847), .B1(ram[14882]), .B2(n3848), 
        .ZN(n19123) );
  MOAI22 U28029 ( .A1(n28526), .A2(n3847), .B1(ram[14883]), .B2(n3848), 
        .ZN(n19124) );
  MOAI22 U28030 ( .A1(n28291), .A2(n3847), .B1(ram[14884]), .B2(n3848), 
        .ZN(n19125) );
  MOAI22 U28031 ( .A1(n28056), .A2(n3847), .B1(ram[14885]), .B2(n3848), 
        .ZN(n19126) );
  MOAI22 U28032 ( .A1(n27821), .A2(n3847), .B1(ram[14886]), .B2(n3848), 
        .ZN(n19127) );
  MOAI22 U28033 ( .A1(n27586), .A2(n3847), .B1(ram[14887]), .B2(n3848), 
        .ZN(n19128) );
  MOAI22 U28034 ( .A1(n29231), .A2(n3849), .B1(ram[14888]), .B2(n3850), 
        .ZN(n19129) );
  MOAI22 U28035 ( .A1(n28996), .A2(n3849), .B1(ram[14889]), .B2(n3850), 
        .ZN(n19130) );
  MOAI22 U28036 ( .A1(n28761), .A2(n3849), .B1(ram[14890]), .B2(n3850), 
        .ZN(n19131) );
  MOAI22 U28037 ( .A1(n28526), .A2(n3849), .B1(ram[14891]), .B2(n3850), 
        .ZN(n19132) );
  MOAI22 U28038 ( .A1(n28291), .A2(n3849), .B1(ram[14892]), .B2(n3850), 
        .ZN(n19133) );
  MOAI22 U28039 ( .A1(n28056), .A2(n3849), .B1(ram[14893]), .B2(n3850), 
        .ZN(n19134) );
  MOAI22 U28040 ( .A1(n27821), .A2(n3849), .B1(ram[14894]), .B2(n3850), 
        .ZN(n19135) );
  MOAI22 U28041 ( .A1(n27586), .A2(n3849), .B1(ram[14895]), .B2(n3850), 
        .ZN(n19136) );
  MOAI22 U28042 ( .A1(n29231), .A2(n3851), .B1(ram[14896]), .B2(n3852), 
        .ZN(n19137) );
  MOAI22 U28043 ( .A1(n28996), .A2(n3851), .B1(ram[14897]), .B2(n3852), 
        .ZN(n19138) );
  MOAI22 U28044 ( .A1(n28761), .A2(n3851), .B1(ram[14898]), .B2(n3852), 
        .ZN(n19139) );
  MOAI22 U28045 ( .A1(n28526), .A2(n3851), .B1(ram[14899]), .B2(n3852), 
        .ZN(n19140) );
  MOAI22 U28046 ( .A1(n28291), .A2(n3851), .B1(ram[14900]), .B2(n3852), 
        .ZN(n19141) );
  MOAI22 U28047 ( .A1(n28056), .A2(n3851), .B1(ram[14901]), .B2(n3852), 
        .ZN(n19142) );
  MOAI22 U28048 ( .A1(n27821), .A2(n3851), .B1(ram[14902]), .B2(n3852), 
        .ZN(n19143) );
  MOAI22 U28049 ( .A1(n27586), .A2(n3851), .B1(ram[14903]), .B2(n3852), 
        .ZN(n19144) );
  MOAI22 U28050 ( .A1(n29231), .A2(n3853), .B1(ram[14904]), .B2(n3854), 
        .ZN(n19145) );
  MOAI22 U28051 ( .A1(n28996), .A2(n3853), .B1(ram[14905]), .B2(n3854), 
        .ZN(n19146) );
  MOAI22 U28052 ( .A1(n28761), .A2(n3853), .B1(ram[14906]), .B2(n3854), 
        .ZN(n19147) );
  MOAI22 U28053 ( .A1(n28526), .A2(n3853), .B1(ram[14907]), .B2(n3854), 
        .ZN(n19148) );
  MOAI22 U28054 ( .A1(n28291), .A2(n3853), .B1(ram[14908]), .B2(n3854), 
        .ZN(n19149) );
  MOAI22 U28055 ( .A1(n28056), .A2(n3853), .B1(ram[14909]), .B2(n3854), 
        .ZN(n19150) );
  MOAI22 U28056 ( .A1(n27821), .A2(n3853), .B1(ram[14910]), .B2(n3854), 
        .ZN(n19151) );
  MOAI22 U28057 ( .A1(n27586), .A2(n3853), .B1(ram[14911]), .B2(n3854), 
        .ZN(n19152) );
  MOAI22 U28058 ( .A1(n29231), .A2(n3855), .B1(ram[14912]), .B2(n3856), 
        .ZN(n19153) );
  MOAI22 U28059 ( .A1(n28996), .A2(n3855), .B1(ram[14913]), .B2(n3856), 
        .ZN(n19154) );
  MOAI22 U28060 ( .A1(n28761), .A2(n3855), .B1(ram[14914]), .B2(n3856), 
        .ZN(n19155) );
  MOAI22 U28061 ( .A1(n28526), .A2(n3855), .B1(ram[14915]), .B2(n3856), 
        .ZN(n19156) );
  MOAI22 U28062 ( .A1(n28291), .A2(n3855), .B1(ram[14916]), .B2(n3856), 
        .ZN(n19157) );
  MOAI22 U28063 ( .A1(n28056), .A2(n3855), .B1(ram[14917]), .B2(n3856), 
        .ZN(n19158) );
  MOAI22 U28064 ( .A1(n27821), .A2(n3855), .B1(ram[14918]), .B2(n3856), 
        .ZN(n19159) );
  MOAI22 U28065 ( .A1(n27586), .A2(n3855), .B1(ram[14919]), .B2(n3856), 
        .ZN(n19160) );
  MOAI22 U28066 ( .A1(n29231), .A2(n3857), .B1(ram[14920]), .B2(n3858), 
        .ZN(n19161) );
  MOAI22 U28067 ( .A1(n28996), .A2(n3857), .B1(ram[14921]), .B2(n3858), 
        .ZN(n19162) );
  MOAI22 U28068 ( .A1(n28761), .A2(n3857), .B1(ram[14922]), .B2(n3858), 
        .ZN(n19163) );
  MOAI22 U28069 ( .A1(n28526), .A2(n3857), .B1(ram[14923]), .B2(n3858), 
        .ZN(n19164) );
  MOAI22 U28070 ( .A1(n28291), .A2(n3857), .B1(ram[14924]), .B2(n3858), 
        .ZN(n19165) );
  MOAI22 U28071 ( .A1(n28056), .A2(n3857), .B1(ram[14925]), .B2(n3858), 
        .ZN(n19166) );
  MOAI22 U28072 ( .A1(n27821), .A2(n3857), .B1(ram[14926]), .B2(n3858), 
        .ZN(n19167) );
  MOAI22 U28073 ( .A1(n27586), .A2(n3857), .B1(ram[14927]), .B2(n3858), 
        .ZN(n19168) );
  MOAI22 U28074 ( .A1(n29231), .A2(n3859), .B1(ram[14928]), .B2(n3860), 
        .ZN(n19169) );
  MOAI22 U28075 ( .A1(n28996), .A2(n3859), .B1(ram[14929]), .B2(n3860), 
        .ZN(n19170) );
  MOAI22 U28076 ( .A1(n28761), .A2(n3859), .B1(ram[14930]), .B2(n3860), 
        .ZN(n19171) );
  MOAI22 U28077 ( .A1(n28526), .A2(n3859), .B1(ram[14931]), .B2(n3860), 
        .ZN(n19172) );
  MOAI22 U28078 ( .A1(n28291), .A2(n3859), .B1(ram[14932]), .B2(n3860), 
        .ZN(n19173) );
  MOAI22 U28079 ( .A1(n28056), .A2(n3859), .B1(ram[14933]), .B2(n3860), 
        .ZN(n19174) );
  MOAI22 U28080 ( .A1(n27821), .A2(n3859), .B1(ram[14934]), .B2(n3860), 
        .ZN(n19175) );
  MOAI22 U28081 ( .A1(n27586), .A2(n3859), .B1(ram[14935]), .B2(n3860), 
        .ZN(n19176) );
  MOAI22 U28082 ( .A1(n29231), .A2(n3861), .B1(ram[14936]), .B2(n3862), 
        .ZN(n19177) );
  MOAI22 U28083 ( .A1(n28996), .A2(n3861), .B1(ram[14937]), .B2(n3862), 
        .ZN(n19178) );
  MOAI22 U28084 ( .A1(n28761), .A2(n3861), .B1(ram[14938]), .B2(n3862), 
        .ZN(n19179) );
  MOAI22 U28085 ( .A1(n28526), .A2(n3861), .B1(ram[14939]), .B2(n3862), 
        .ZN(n19180) );
  MOAI22 U28086 ( .A1(n28291), .A2(n3861), .B1(ram[14940]), .B2(n3862), 
        .ZN(n19181) );
  MOAI22 U28087 ( .A1(n28056), .A2(n3861), .B1(ram[14941]), .B2(n3862), 
        .ZN(n19182) );
  MOAI22 U28088 ( .A1(n27821), .A2(n3861), .B1(ram[14942]), .B2(n3862), 
        .ZN(n19183) );
  MOAI22 U28089 ( .A1(n27586), .A2(n3861), .B1(ram[14943]), .B2(n3862), 
        .ZN(n19184) );
  MOAI22 U28090 ( .A1(n29231), .A2(n3863), .B1(ram[14944]), .B2(n3864), 
        .ZN(n19185) );
  MOAI22 U28091 ( .A1(n28996), .A2(n3863), .B1(ram[14945]), .B2(n3864), 
        .ZN(n19186) );
  MOAI22 U28092 ( .A1(n28761), .A2(n3863), .B1(ram[14946]), .B2(n3864), 
        .ZN(n19187) );
  MOAI22 U28093 ( .A1(n28526), .A2(n3863), .B1(ram[14947]), .B2(n3864), 
        .ZN(n19188) );
  MOAI22 U28094 ( .A1(n28291), .A2(n3863), .B1(ram[14948]), .B2(n3864), 
        .ZN(n19189) );
  MOAI22 U28095 ( .A1(n28056), .A2(n3863), .B1(ram[14949]), .B2(n3864), 
        .ZN(n19190) );
  MOAI22 U28096 ( .A1(n27821), .A2(n3863), .B1(ram[14950]), .B2(n3864), 
        .ZN(n19191) );
  MOAI22 U28097 ( .A1(n27586), .A2(n3863), .B1(ram[14951]), .B2(n3864), 
        .ZN(n19192) );
  MOAI22 U28098 ( .A1(n29231), .A2(n3865), .B1(ram[14952]), .B2(n3866), 
        .ZN(n19193) );
  MOAI22 U28099 ( .A1(n28996), .A2(n3865), .B1(ram[14953]), .B2(n3866), 
        .ZN(n19194) );
  MOAI22 U28100 ( .A1(n28761), .A2(n3865), .B1(ram[14954]), .B2(n3866), 
        .ZN(n19195) );
  MOAI22 U28101 ( .A1(n28526), .A2(n3865), .B1(ram[14955]), .B2(n3866), 
        .ZN(n19196) );
  MOAI22 U28102 ( .A1(n28291), .A2(n3865), .B1(ram[14956]), .B2(n3866), 
        .ZN(n19197) );
  MOAI22 U28103 ( .A1(n28056), .A2(n3865), .B1(ram[14957]), .B2(n3866), 
        .ZN(n19198) );
  MOAI22 U28104 ( .A1(n27821), .A2(n3865), .B1(ram[14958]), .B2(n3866), 
        .ZN(n19199) );
  MOAI22 U28105 ( .A1(n27586), .A2(n3865), .B1(ram[14959]), .B2(n3866), 
        .ZN(n19200) );
  MOAI22 U28106 ( .A1(n29231), .A2(n3867), .B1(ram[14960]), .B2(n3868), 
        .ZN(n19201) );
  MOAI22 U28107 ( .A1(n28996), .A2(n3867), .B1(ram[14961]), .B2(n3868), 
        .ZN(n19202) );
  MOAI22 U28108 ( .A1(n28761), .A2(n3867), .B1(ram[14962]), .B2(n3868), 
        .ZN(n19203) );
  MOAI22 U28109 ( .A1(n28526), .A2(n3867), .B1(ram[14963]), .B2(n3868), 
        .ZN(n19204) );
  MOAI22 U28110 ( .A1(n28291), .A2(n3867), .B1(ram[14964]), .B2(n3868), 
        .ZN(n19205) );
  MOAI22 U28111 ( .A1(n28056), .A2(n3867), .B1(ram[14965]), .B2(n3868), 
        .ZN(n19206) );
  MOAI22 U28112 ( .A1(n27821), .A2(n3867), .B1(ram[14966]), .B2(n3868), 
        .ZN(n19207) );
  MOAI22 U28113 ( .A1(n27586), .A2(n3867), .B1(ram[14967]), .B2(n3868), 
        .ZN(n19208) );
  MOAI22 U28114 ( .A1(n29231), .A2(n3869), .B1(ram[14968]), .B2(n3870), 
        .ZN(n19209) );
  MOAI22 U28115 ( .A1(n28996), .A2(n3869), .B1(ram[14969]), .B2(n3870), 
        .ZN(n19210) );
  MOAI22 U28116 ( .A1(n28761), .A2(n3869), .B1(ram[14970]), .B2(n3870), 
        .ZN(n19211) );
  MOAI22 U28117 ( .A1(n28526), .A2(n3869), .B1(ram[14971]), .B2(n3870), 
        .ZN(n19212) );
  MOAI22 U28118 ( .A1(n28291), .A2(n3869), .B1(ram[14972]), .B2(n3870), 
        .ZN(n19213) );
  MOAI22 U28119 ( .A1(n28056), .A2(n3869), .B1(ram[14973]), .B2(n3870), 
        .ZN(n19214) );
  MOAI22 U28120 ( .A1(n27821), .A2(n3869), .B1(ram[14974]), .B2(n3870), 
        .ZN(n19215) );
  MOAI22 U28121 ( .A1(n27586), .A2(n3869), .B1(ram[14975]), .B2(n3870), 
        .ZN(n19216) );
  MOAI22 U28122 ( .A1(n29232), .A2(n3871), .B1(ram[14976]), .B2(n3872), 
        .ZN(n19217) );
  MOAI22 U28123 ( .A1(n28997), .A2(n3871), .B1(ram[14977]), .B2(n3872), 
        .ZN(n19218) );
  MOAI22 U28124 ( .A1(n28762), .A2(n3871), .B1(ram[14978]), .B2(n3872), 
        .ZN(n19219) );
  MOAI22 U28125 ( .A1(n28527), .A2(n3871), .B1(ram[14979]), .B2(n3872), 
        .ZN(n19220) );
  MOAI22 U28126 ( .A1(n28292), .A2(n3871), .B1(ram[14980]), .B2(n3872), 
        .ZN(n19221) );
  MOAI22 U28127 ( .A1(n28057), .A2(n3871), .B1(ram[14981]), .B2(n3872), 
        .ZN(n19222) );
  MOAI22 U28128 ( .A1(n27822), .A2(n3871), .B1(ram[14982]), .B2(n3872), 
        .ZN(n19223) );
  MOAI22 U28129 ( .A1(n27587), .A2(n3871), .B1(ram[14983]), .B2(n3872), 
        .ZN(n19224) );
  MOAI22 U28130 ( .A1(n29232), .A2(n3873), .B1(ram[14984]), .B2(n3874), 
        .ZN(n19225) );
  MOAI22 U28131 ( .A1(n28997), .A2(n3873), .B1(ram[14985]), .B2(n3874), 
        .ZN(n19226) );
  MOAI22 U28132 ( .A1(n28762), .A2(n3873), .B1(ram[14986]), .B2(n3874), 
        .ZN(n19227) );
  MOAI22 U28133 ( .A1(n28527), .A2(n3873), .B1(ram[14987]), .B2(n3874), 
        .ZN(n19228) );
  MOAI22 U28134 ( .A1(n28292), .A2(n3873), .B1(ram[14988]), .B2(n3874), 
        .ZN(n19229) );
  MOAI22 U28135 ( .A1(n28057), .A2(n3873), .B1(ram[14989]), .B2(n3874), 
        .ZN(n19230) );
  MOAI22 U28136 ( .A1(n27822), .A2(n3873), .B1(ram[14990]), .B2(n3874), 
        .ZN(n19231) );
  MOAI22 U28137 ( .A1(n27587), .A2(n3873), .B1(ram[14991]), .B2(n3874), 
        .ZN(n19232) );
  MOAI22 U28138 ( .A1(n29232), .A2(n3875), .B1(ram[14992]), .B2(n3876), 
        .ZN(n19233) );
  MOAI22 U28139 ( .A1(n28997), .A2(n3875), .B1(ram[14993]), .B2(n3876), 
        .ZN(n19234) );
  MOAI22 U28140 ( .A1(n28762), .A2(n3875), .B1(ram[14994]), .B2(n3876), 
        .ZN(n19235) );
  MOAI22 U28141 ( .A1(n28527), .A2(n3875), .B1(ram[14995]), .B2(n3876), 
        .ZN(n19236) );
  MOAI22 U28142 ( .A1(n28292), .A2(n3875), .B1(ram[14996]), .B2(n3876), 
        .ZN(n19237) );
  MOAI22 U28143 ( .A1(n28057), .A2(n3875), .B1(ram[14997]), .B2(n3876), 
        .ZN(n19238) );
  MOAI22 U28144 ( .A1(n27822), .A2(n3875), .B1(ram[14998]), .B2(n3876), 
        .ZN(n19239) );
  MOAI22 U28145 ( .A1(n27587), .A2(n3875), .B1(ram[14999]), .B2(n3876), 
        .ZN(n19240) );
  MOAI22 U28146 ( .A1(n29232), .A2(n3877), .B1(ram[15000]), .B2(n3878), 
        .ZN(n19241) );
  MOAI22 U28147 ( .A1(n28997), .A2(n3877), .B1(ram[15001]), .B2(n3878), 
        .ZN(n19242) );
  MOAI22 U28148 ( .A1(n28762), .A2(n3877), .B1(ram[15002]), .B2(n3878), 
        .ZN(n19243) );
  MOAI22 U28149 ( .A1(n28527), .A2(n3877), .B1(ram[15003]), .B2(n3878), 
        .ZN(n19244) );
  MOAI22 U28150 ( .A1(n28292), .A2(n3877), .B1(ram[15004]), .B2(n3878), 
        .ZN(n19245) );
  MOAI22 U28151 ( .A1(n28057), .A2(n3877), .B1(ram[15005]), .B2(n3878), 
        .ZN(n19246) );
  MOAI22 U28152 ( .A1(n27822), .A2(n3877), .B1(ram[15006]), .B2(n3878), 
        .ZN(n19247) );
  MOAI22 U28153 ( .A1(n27587), .A2(n3877), .B1(ram[15007]), .B2(n3878), 
        .ZN(n19248) );
  MOAI22 U28154 ( .A1(n29232), .A2(n3879), .B1(ram[15008]), .B2(n3880), 
        .ZN(n19249) );
  MOAI22 U28155 ( .A1(n28997), .A2(n3879), .B1(ram[15009]), .B2(n3880), 
        .ZN(n19250) );
  MOAI22 U28156 ( .A1(n28762), .A2(n3879), .B1(ram[15010]), .B2(n3880), 
        .ZN(n19251) );
  MOAI22 U28157 ( .A1(n28527), .A2(n3879), .B1(ram[15011]), .B2(n3880), 
        .ZN(n19252) );
  MOAI22 U28158 ( .A1(n28292), .A2(n3879), .B1(ram[15012]), .B2(n3880), 
        .ZN(n19253) );
  MOAI22 U28159 ( .A1(n28057), .A2(n3879), .B1(ram[15013]), .B2(n3880), 
        .ZN(n19254) );
  MOAI22 U28160 ( .A1(n27822), .A2(n3879), .B1(ram[15014]), .B2(n3880), 
        .ZN(n19255) );
  MOAI22 U28161 ( .A1(n27587), .A2(n3879), .B1(ram[15015]), .B2(n3880), 
        .ZN(n19256) );
  MOAI22 U28162 ( .A1(n29232), .A2(n3881), .B1(ram[15016]), .B2(n3882), 
        .ZN(n19257) );
  MOAI22 U28163 ( .A1(n28997), .A2(n3881), .B1(ram[15017]), .B2(n3882), 
        .ZN(n19258) );
  MOAI22 U28164 ( .A1(n28762), .A2(n3881), .B1(ram[15018]), .B2(n3882), 
        .ZN(n19259) );
  MOAI22 U28165 ( .A1(n28527), .A2(n3881), .B1(ram[15019]), .B2(n3882), 
        .ZN(n19260) );
  MOAI22 U28166 ( .A1(n28292), .A2(n3881), .B1(ram[15020]), .B2(n3882), 
        .ZN(n19261) );
  MOAI22 U28167 ( .A1(n28057), .A2(n3881), .B1(ram[15021]), .B2(n3882), 
        .ZN(n19262) );
  MOAI22 U28168 ( .A1(n27822), .A2(n3881), .B1(ram[15022]), .B2(n3882), 
        .ZN(n19263) );
  MOAI22 U28169 ( .A1(n27587), .A2(n3881), .B1(ram[15023]), .B2(n3882), 
        .ZN(n19264) );
  MOAI22 U28170 ( .A1(n29232), .A2(n3883), .B1(ram[15024]), .B2(n3884), 
        .ZN(n19265) );
  MOAI22 U28171 ( .A1(n28997), .A2(n3883), .B1(ram[15025]), .B2(n3884), 
        .ZN(n19266) );
  MOAI22 U28172 ( .A1(n28762), .A2(n3883), .B1(ram[15026]), .B2(n3884), 
        .ZN(n19267) );
  MOAI22 U28173 ( .A1(n28527), .A2(n3883), .B1(ram[15027]), .B2(n3884), 
        .ZN(n19268) );
  MOAI22 U28174 ( .A1(n28292), .A2(n3883), .B1(ram[15028]), .B2(n3884), 
        .ZN(n19269) );
  MOAI22 U28175 ( .A1(n28057), .A2(n3883), .B1(ram[15029]), .B2(n3884), 
        .ZN(n19270) );
  MOAI22 U28176 ( .A1(n27822), .A2(n3883), .B1(ram[15030]), .B2(n3884), 
        .ZN(n19271) );
  MOAI22 U28177 ( .A1(n27587), .A2(n3883), .B1(ram[15031]), .B2(n3884), 
        .ZN(n19272) );
  MOAI22 U28178 ( .A1(n29232), .A2(n3885), .B1(ram[15032]), .B2(n3886), 
        .ZN(n19273) );
  MOAI22 U28179 ( .A1(n28997), .A2(n3885), .B1(ram[15033]), .B2(n3886), 
        .ZN(n19274) );
  MOAI22 U28180 ( .A1(n28762), .A2(n3885), .B1(ram[15034]), .B2(n3886), 
        .ZN(n19275) );
  MOAI22 U28181 ( .A1(n28527), .A2(n3885), .B1(ram[15035]), .B2(n3886), 
        .ZN(n19276) );
  MOAI22 U28182 ( .A1(n28292), .A2(n3885), .B1(ram[15036]), .B2(n3886), 
        .ZN(n19277) );
  MOAI22 U28183 ( .A1(n28057), .A2(n3885), .B1(ram[15037]), .B2(n3886), 
        .ZN(n19278) );
  MOAI22 U28184 ( .A1(n27822), .A2(n3885), .B1(ram[15038]), .B2(n3886), 
        .ZN(n19279) );
  MOAI22 U28185 ( .A1(n27587), .A2(n3885), .B1(ram[15039]), .B2(n3886), 
        .ZN(n19280) );
  MOAI22 U28186 ( .A1(n29232), .A2(n3887), .B1(ram[15040]), .B2(n3888), 
        .ZN(n19281) );
  MOAI22 U28187 ( .A1(n28997), .A2(n3887), .B1(ram[15041]), .B2(n3888), 
        .ZN(n19282) );
  MOAI22 U28188 ( .A1(n28762), .A2(n3887), .B1(ram[15042]), .B2(n3888), 
        .ZN(n19283) );
  MOAI22 U28189 ( .A1(n28527), .A2(n3887), .B1(ram[15043]), .B2(n3888), 
        .ZN(n19284) );
  MOAI22 U28190 ( .A1(n28292), .A2(n3887), .B1(ram[15044]), .B2(n3888), 
        .ZN(n19285) );
  MOAI22 U28191 ( .A1(n28057), .A2(n3887), .B1(ram[15045]), .B2(n3888), 
        .ZN(n19286) );
  MOAI22 U28192 ( .A1(n27822), .A2(n3887), .B1(ram[15046]), .B2(n3888), 
        .ZN(n19287) );
  MOAI22 U28193 ( .A1(n27587), .A2(n3887), .B1(ram[15047]), .B2(n3888), 
        .ZN(n19288) );
  MOAI22 U28194 ( .A1(n29232), .A2(n3889), .B1(ram[15048]), .B2(n3890), 
        .ZN(n19289) );
  MOAI22 U28195 ( .A1(n28997), .A2(n3889), .B1(ram[15049]), .B2(n3890), 
        .ZN(n19290) );
  MOAI22 U28196 ( .A1(n28762), .A2(n3889), .B1(ram[15050]), .B2(n3890), 
        .ZN(n19291) );
  MOAI22 U28197 ( .A1(n28527), .A2(n3889), .B1(ram[15051]), .B2(n3890), 
        .ZN(n19292) );
  MOAI22 U28198 ( .A1(n28292), .A2(n3889), .B1(ram[15052]), .B2(n3890), 
        .ZN(n19293) );
  MOAI22 U28199 ( .A1(n28057), .A2(n3889), .B1(ram[15053]), .B2(n3890), 
        .ZN(n19294) );
  MOAI22 U28200 ( .A1(n27822), .A2(n3889), .B1(ram[15054]), .B2(n3890), 
        .ZN(n19295) );
  MOAI22 U28201 ( .A1(n27587), .A2(n3889), .B1(ram[15055]), .B2(n3890), 
        .ZN(n19296) );
  MOAI22 U28202 ( .A1(n29232), .A2(n3891), .B1(ram[15056]), .B2(n3892), 
        .ZN(n19297) );
  MOAI22 U28203 ( .A1(n28997), .A2(n3891), .B1(ram[15057]), .B2(n3892), 
        .ZN(n19298) );
  MOAI22 U28204 ( .A1(n28762), .A2(n3891), .B1(ram[15058]), .B2(n3892), 
        .ZN(n19299) );
  MOAI22 U28205 ( .A1(n28527), .A2(n3891), .B1(ram[15059]), .B2(n3892), 
        .ZN(n19300) );
  MOAI22 U28206 ( .A1(n28292), .A2(n3891), .B1(ram[15060]), .B2(n3892), 
        .ZN(n19301) );
  MOAI22 U28207 ( .A1(n28057), .A2(n3891), .B1(ram[15061]), .B2(n3892), 
        .ZN(n19302) );
  MOAI22 U28208 ( .A1(n27822), .A2(n3891), .B1(ram[15062]), .B2(n3892), 
        .ZN(n19303) );
  MOAI22 U28209 ( .A1(n27587), .A2(n3891), .B1(ram[15063]), .B2(n3892), 
        .ZN(n19304) );
  MOAI22 U28210 ( .A1(n29232), .A2(n3893), .B1(ram[15064]), .B2(n3894), 
        .ZN(n19305) );
  MOAI22 U28211 ( .A1(n28997), .A2(n3893), .B1(ram[15065]), .B2(n3894), 
        .ZN(n19306) );
  MOAI22 U28212 ( .A1(n28762), .A2(n3893), .B1(ram[15066]), .B2(n3894), 
        .ZN(n19307) );
  MOAI22 U28213 ( .A1(n28527), .A2(n3893), .B1(ram[15067]), .B2(n3894), 
        .ZN(n19308) );
  MOAI22 U28214 ( .A1(n28292), .A2(n3893), .B1(ram[15068]), .B2(n3894), 
        .ZN(n19309) );
  MOAI22 U28215 ( .A1(n28057), .A2(n3893), .B1(ram[15069]), .B2(n3894), 
        .ZN(n19310) );
  MOAI22 U28216 ( .A1(n27822), .A2(n3893), .B1(ram[15070]), .B2(n3894), 
        .ZN(n19311) );
  MOAI22 U28217 ( .A1(n27587), .A2(n3893), .B1(ram[15071]), .B2(n3894), 
        .ZN(n19312) );
  MOAI22 U28218 ( .A1(n29232), .A2(n3895), .B1(ram[15072]), .B2(n3896), 
        .ZN(n19313) );
  MOAI22 U28219 ( .A1(n28997), .A2(n3895), .B1(ram[15073]), .B2(n3896), 
        .ZN(n19314) );
  MOAI22 U28220 ( .A1(n28762), .A2(n3895), .B1(ram[15074]), .B2(n3896), 
        .ZN(n19315) );
  MOAI22 U28221 ( .A1(n28527), .A2(n3895), .B1(ram[15075]), .B2(n3896), 
        .ZN(n19316) );
  MOAI22 U28222 ( .A1(n28292), .A2(n3895), .B1(ram[15076]), .B2(n3896), 
        .ZN(n19317) );
  MOAI22 U28223 ( .A1(n28057), .A2(n3895), .B1(ram[15077]), .B2(n3896), 
        .ZN(n19318) );
  MOAI22 U28224 ( .A1(n27822), .A2(n3895), .B1(ram[15078]), .B2(n3896), 
        .ZN(n19319) );
  MOAI22 U28225 ( .A1(n27587), .A2(n3895), .B1(ram[15079]), .B2(n3896), 
        .ZN(n19320) );
  MOAI22 U28226 ( .A1(n29233), .A2(n3897), .B1(ram[15080]), .B2(n3898), 
        .ZN(n19321) );
  MOAI22 U28227 ( .A1(n28998), .A2(n3897), .B1(ram[15081]), .B2(n3898), 
        .ZN(n19322) );
  MOAI22 U28228 ( .A1(n28763), .A2(n3897), .B1(ram[15082]), .B2(n3898), 
        .ZN(n19323) );
  MOAI22 U28229 ( .A1(n28528), .A2(n3897), .B1(ram[15083]), .B2(n3898), 
        .ZN(n19324) );
  MOAI22 U28230 ( .A1(n28293), .A2(n3897), .B1(ram[15084]), .B2(n3898), 
        .ZN(n19325) );
  MOAI22 U28231 ( .A1(n28058), .A2(n3897), .B1(ram[15085]), .B2(n3898), 
        .ZN(n19326) );
  MOAI22 U28232 ( .A1(n27823), .A2(n3897), .B1(ram[15086]), .B2(n3898), 
        .ZN(n19327) );
  MOAI22 U28233 ( .A1(n27588), .A2(n3897), .B1(ram[15087]), .B2(n3898), 
        .ZN(n19328) );
  MOAI22 U28234 ( .A1(n29233), .A2(n3899), .B1(ram[15088]), .B2(n3900), 
        .ZN(n19329) );
  MOAI22 U28235 ( .A1(n28998), .A2(n3899), .B1(ram[15089]), .B2(n3900), 
        .ZN(n19330) );
  MOAI22 U28236 ( .A1(n28763), .A2(n3899), .B1(ram[15090]), .B2(n3900), 
        .ZN(n19331) );
  MOAI22 U28237 ( .A1(n28528), .A2(n3899), .B1(ram[15091]), .B2(n3900), 
        .ZN(n19332) );
  MOAI22 U28238 ( .A1(n28293), .A2(n3899), .B1(ram[15092]), .B2(n3900), 
        .ZN(n19333) );
  MOAI22 U28239 ( .A1(n28058), .A2(n3899), .B1(ram[15093]), .B2(n3900), 
        .ZN(n19334) );
  MOAI22 U28240 ( .A1(n27823), .A2(n3899), .B1(ram[15094]), .B2(n3900), 
        .ZN(n19335) );
  MOAI22 U28241 ( .A1(n27588), .A2(n3899), .B1(ram[15095]), .B2(n3900), 
        .ZN(n19336) );
  MOAI22 U28242 ( .A1(n29233), .A2(n3901), .B1(ram[15096]), .B2(n3902), 
        .ZN(n19337) );
  MOAI22 U28243 ( .A1(n28998), .A2(n3901), .B1(ram[15097]), .B2(n3902), 
        .ZN(n19338) );
  MOAI22 U28244 ( .A1(n28763), .A2(n3901), .B1(ram[15098]), .B2(n3902), 
        .ZN(n19339) );
  MOAI22 U28245 ( .A1(n28528), .A2(n3901), .B1(ram[15099]), .B2(n3902), 
        .ZN(n19340) );
  MOAI22 U28246 ( .A1(n28293), .A2(n3901), .B1(ram[15100]), .B2(n3902), 
        .ZN(n19341) );
  MOAI22 U28247 ( .A1(n28058), .A2(n3901), .B1(ram[15101]), .B2(n3902), 
        .ZN(n19342) );
  MOAI22 U28248 ( .A1(n27823), .A2(n3901), .B1(ram[15102]), .B2(n3902), 
        .ZN(n19343) );
  MOAI22 U28249 ( .A1(n27588), .A2(n3901), .B1(ram[15103]), .B2(n3902), 
        .ZN(n19344) );
  MOAI22 U28250 ( .A1(n29233), .A2(n3903), .B1(ram[15104]), .B2(n3904), 
        .ZN(n19345) );
  MOAI22 U28251 ( .A1(n28998), .A2(n3903), .B1(ram[15105]), .B2(n3904), 
        .ZN(n19346) );
  MOAI22 U28252 ( .A1(n28763), .A2(n3903), .B1(ram[15106]), .B2(n3904), 
        .ZN(n19347) );
  MOAI22 U28253 ( .A1(n28528), .A2(n3903), .B1(ram[15107]), .B2(n3904), 
        .ZN(n19348) );
  MOAI22 U28254 ( .A1(n28293), .A2(n3903), .B1(ram[15108]), .B2(n3904), 
        .ZN(n19349) );
  MOAI22 U28255 ( .A1(n28058), .A2(n3903), .B1(ram[15109]), .B2(n3904), 
        .ZN(n19350) );
  MOAI22 U28256 ( .A1(n27823), .A2(n3903), .B1(ram[15110]), .B2(n3904), 
        .ZN(n19351) );
  MOAI22 U28257 ( .A1(n27588), .A2(n3903), .B1(ram[15111]), .B2(n3904), 
        .ZN(n19352) );
  MOAI22 U28258 ( .A1(n29233), .A2(n3905), .B1(ram[15112]), .B2(n3906), 
        .ZN(n19353) );
  MOAI22 U28259 ( .A1(n28998), .A2(n3905), .B1(ram[15113]), .B2(n3906), 
        .ZN(n19354) );
  MOAI22 U28260 ( .A1(n28763), .A2(n3905), .B1(ram[15114]), .B2(n3906), 
        .ZN(n19355) );
  MOAI22 U28261 ( .A1(n28528), .A2(n3905), .B1(ram[15115]), .B2(n3906), 
        .ZN(n19356) );
  MOAI22 U28262 ( .A1(n28293), .A2(n3905), .B1(ram[15116]), .B2(n3906), 
        .ZN(n19357) );
  MOAI22 U28263 ( .A1(n28058), .A2(n3905), .B1(ram[15117]), .B2(n3906), 
        .ZN(n19358) );
  MOAI22 U28264 ( .A1(n27823), .A2(n3905), .B1(ram[15118]), .B2(n3906), 
        .ZN(n19359) );
  MOAI22 U28265 ( .A1(n27588), .A2(n3905), .B1(ram[15119]), .B2(n3906), 
        .ZN(n19360) );
  MOAI22 U28266 ( .A1(n29233), .A2(n3907), .B1(ram[15120]), .B2(n3908), 
        .ZN(n19361) );
  MOAI22 U28267 ( .A1(n28998), .A2(n3907), .B1(ram[15121]), .B2(n3908), 
        .ZN(n19362) );
  MOAI22 U28268 ( .A1(n28763), .A2(n3907), .B1(ram[15122]), .B2(n3908), 
        .ZN(n19363) );
  MOAI22 U28269 ( .A1(n28528), .A2(n3907), .B1(ram[15123]), .B2(n3908), 
        .ZN(n19364) );
  MOAI22 U28270 ( .A1(n28293), .A2(n3907), .B1(ram[15124]), .B2(n3908), 
        .ZN(n19365) );
  MOAI22 U28271 ( .A1(n28058), .A2(n3907), .B1(ram[15125]), .B2(n3908), 
        .ZN(n19366) );
  MOAI22 U28272 ( .A1(n27823), .A2(n3907), .B1(ram[15126]), .B2(n3908), 
        .ZN(n19367) );
  MOAI22 U28273 ( .A1(n27588), .A2(n3907), .B1(ram[15127]), .B2(n3908), 
        .ZN(n19368) );
  MOAI22 U28274 ( .A1(n29233), .A2(n3909), .B1(ram[15128]), .B2(n3910), 
        .ZN(n19369) );
  MOAI22 U28275 ( .A1(n28998), .A2(n3909), .B1(ram[15129]), .B2(n3910), 
        .ZN(n19370) );
  MOAI22 U28276 ( .A1(n28763), .A2(n3909), .B1(ram[15130]), .B2(n3910), 
        .ZN(n19371) );
  MOAI22 U28277 ( .A1(n28528), .A2(n3909), .B1(ram[15131]), .B2(n3910), 
        .ZN(n19372) );
  MOAI22 U28278 ( .A1(n28293), .A2(n3909), .B1(ram[15132]), .B2(n3910), 
        .ZN(n19373) );
  MOAI22 U28279 ( .A1(n28058), .A2(n3909), .B1(ram[15133]), .B2(n3910), 
        .ZN(n19374) );
  MOAI22 U28280 ( .A1(n27823), .A2(n3909), .B1(ram[15134]), .B2(n3910), 
        .ZN(n19375) );
  MOAI22 U28281 ( .A1(n27588), .A2(n3909), .B1(ram[15135]), .B2(n3910), 
        .ZN(n19376) );
  MOAI22 U28282 ( .A1(n29233), .A2(n3911), .B1(ram[15136]), .B2(n3912), 
        .ZN(n19377) );
  MOAI22 U28283 ( .A1(n28998), .A2(n3911), .B1(ram[15137]), .B2(n3912), 
        .ZN(n19378) );
  MOAI22 U28284 ( .A1(n28763), .A2(n3911), .B1(ram[15138]), .B2(n3912), 
        .ZN(n19379) );
  MOAI22 U28285 ( .A1(n28528), .A2(n3911), .B1(ram[15139]), .B2(n3912), 
        .ZN(n19380) );
  MOAI22 U28286 ( .A1(n28293), .A2(n3911), .B1(ram[15140]), .B2(n3912), 
        .ZN(n19381) );
  MOAI22 U28287 ( .A1(n28058), .A2(n3911), .B1(ram[15141]), .B2(n3912), 
        .ZN(n19382) );
  MOAI22 U28288 ( .A1(n27823), .A2(n3911), .B1(ram[15142]), .B2(n3912), 
        .ZN(n19383) );
  MOAI22 U28289 ( .A1(n27588), .A2(n3911), .B1(ram[15143]), .B2(n3912), 
        .ZN(n19384) );
  MOAI22 U28290 ( .A1(n29233), .A2(n3913), .B1(ram[15144]), .B2(n3914), 
        .ZN(n19385) );
  MOAI22 U28291 ( .A1(n28998), .A2(n3913), .B1(ram[15145]), .B2(n3914), 
        .ZN(n19386) );
  MOAI22 U28292 ( .A1(n28763), .A2(n3913), .B1(ram[15146]), .B2(n3914), 
        .ZN(n19387) );
  MOAI22 U28293 ( .A1(n28528), .A2(n3913), .B1(ram[15147]), .B2(n3914), 
        .ZN(n19388) );
  MOAI22 U28294 ( .A1(n28293), .A2(n3913), .B1(ram[15148]), .B2(n3914), 
        .ZN(n19389) );
  MOAI22 U28295 ( .A1(n28058), .A2(n3913), .B1(ram[15149]), .B2(n3914), 
        .ZN(n19390) );
  MOAI22 U28296 ( .A1(n27823), .A2(n3913), .B1(ram[15150]), .B2(n3914), 
        .ZN(n19391) );
  MOAI22 U28297 ( .A1(n27588), .A2(n3913), .B1(ram[15151]), .B2(n3914), 
        .ZN(n19392) );
  MOAI22 U28298 ( .A1(n29233), .A2(n3915), .B1(ram[15152]), .B2(n3916), 
        .ZN(n19393) );
  MOAI22 U28299 ( .A1(n28998), .A2(n3915), .B1(ram[15153]), .B2(n3916), 
        .ZN(n19394) );
  MOAI22 U28300 ( .A1(n28763), .A2(n3915), .B1(ram[15154]), .B2(n3916), 
        .ZN(n19395) );
  MOAI22 U28301 ( .A1(n28528), .A2(n3915), .B1(ram[15155]), .B2(n3916), 
        .ZN(n19396) );
  MOAI22 U28302 ( .A1(n28293), .A2(n3915), .B1(ram[15156]), .B2(n3916), 
        .ZN(n19397) );
  MOAI22 U28303 ( .A1(n28058), .A2(n3915), .B1(ram[15157]), .B2(n3916), 
        .ZN(n19398) );
  MOAI22 U28304 ( .A1(n27823), .A2(n3915), .B1(ram[15158]), .B2(n3916), 
        .ZN(n19399) );
  MOAI22 U28305 ( .A1(n27588), .A2(n3915), .B1(ram[15159]), .B2(n3916), 
        .ZN(n19400) );
  MOAI22 U28306 ( .A1(n29233), .A2(n3917), .B1(ram[15160]), .B2(n3918), 
        .ZN(n19401) );
  MOAI22 U28307 ( .A1(n28998), .A2(n3917), .B1(ram[15161]), .B2(n3918), 
        .ZN(n19402) );
  MOAI22 U28308 ( .A1(n28763), .A2(n3917), .B1(ram[15162]), .B2(n3918), 
        .ZN(n19403) );
  MOAI22 U28309 ( .A1(n28528), .A2(n3917), .B1(ram[15163]), .B2(n3918), 
        .ZN(n19404) );
  MOAI22 U28310 ( .A1(n28293), .A2(n3917), .B1(ram[15164]), .B2(n3918), 
        .ZN(n19405) );
  MOAI22 U28311 ( .A1(n28058), .A2(n3917), .B1(ram[15165]), .B2(n3918), 
        .ZN(n19406) );
  MOAI22 U28312 ( .A1(n27823), .A2(n3917), .B1(ram[15166]), .B2(n3918), 
        .ZN(n19407) );
  MOAI22 U28313 ( .A1(n27588), .A2(n3917), .B1(ram[15167]), .B2(n3918), 
        .ZN(n19408) );
  MOAI22 U28314 ( .A1(n29233), .A2(n3919), .B1(ram[15168]), .B2(n3920), 
        .ZN(n19409) );
  MOAI22 U28315 ( .A1(n28998), .A2(n3919), .B1(ram[15169]), .B2(n3920), 
        .ZN(n19410) );
  MOAI22 U28316 ( .A1(n28763), .A2(n3919), .B1(ram[15170]), .B2(n3920), 
        .ZN(n19411) );
  MOAI22 U28317 ( .A1(n28528), .A2(n3919), .B1(ram[15171]), .B2(n3920), 
        .ZN(n19412) );
  MOAI22 U28318 ( .A1(n28293), .A2(n3919), .B1(ram[15172]), .B2(n3920), 
        .ZN(n19413) );
  MOAI22 U28319 ( .A1(n28058), .A2(n3919), .B1(ram[15173]), .B2(n3920), 
        .ZN(n19414) );
  MOAI22 U28320 ( .A1(n27823), .A2(n3919), .B1(ram[15174]), .B2(n3920), 
        .ZN(n19415) );
  MOAI22 U28321 ( .A1(n27588), .A2(n3919), .B1(ram[15175]), .B2(n3920), 
        .ZN(n19416) );
  MOAI22 U28322 ( .A1(n29233), .A2(n3921), .B1(ram[15176]), .B2(n3922), 
        .ZN(n19417) );
  MOAI22 U28323 ( .A1(n28998), .A2(n3921), .B1(ram[15177]), .B2(n3922), 
        .ZN(n19418) );
  MOAI22 U28324 ( .A1(n28763), .A2(n3921), .B1(ram[15178]), .B2(n3922), 
        .ZN(n19419) );
  MOAI22 U28325 ( .A1(n28528), .A2(n3921), .B1(ram[15179]), .B2(n3922), 
        .ZN(n19420) );
  MOAI22 U28326 ( .A1(n28293), .A2(n3921), .B1(ram[15180]), .B2(n3922), 
        .ZN(n19421) );
  MOAI22 U28327 ( .A1(n28058), .A2(n3921), .B1(ram[15181]), .B2(n3922), 
        .ZN(n19422) );
  MOAI22 U28328 ( .A1(n27823), .A2(n3921), .B1(ram[15182]), .B2(n3922), 
        .ZN(n19423) );
  MOAI22 U28329 ( .A1(n27588), .A2(n3921), .B1(ram[15183]), .B2(n3922), 
        .ZN(n19424) );
  MOAI22 U28330 ( .A1(n29234), .A2(n3923), .B1(ram[15184]), .B2(n3924), 
        .ZN(n19425) );
  MOAI22 U28331 ( .A1(n28999), .A2(n3923), .B1(ram[15185]), .B2(n3924), 
        .ZN(n19426) );
  MOAI22 U28332 ( .A1(n28764), .A2(n3923), .B1(ram[15186]), .B2(n3924), 
        .ZN(n19427) );
  MOAI22 U28333 ( .A1(n28529), .A2(n3923), .B1(ram[15187]), .B2(n3924), 
        .ZN(n19428) );
  MOAI22 U28334 ( .A1(n28294), .A2(n3923), .B1(ram[15188]), .B2(n3924), 
        .ZN(n19429) );
  MOAI22 U28335 ( .A1(n28059), .A2(n3923), .B1(ram[15189]), .B2(n3924), 
        .ZN(n19430) );
  MOAI22 U28336 ( .A1(n27824), .A2(n3923), .B1(ram[15190]), .B2(n3924), 
        .ZN(n19431) );
  MOAI22 U28337 ( .A1(n27589), .A2(n3923), .B1(ram[15191]), .B2(n3924), 
        .ZN(n19432) );
  MOAI22 U28338 ( .A1(n29234), .A2(n3925), .B1(ram[15192]), .B2(n3926), 
        .ZN(n19433) );
  MOAI22 U28339 ( .A1(n28999), .A2(n3925), .B1(ram[15193]), .B2(n3926), 
        .ZN(n19434) );
  MOAI22 U28340 ( .A1(n28764), .A2(n3925), .B1(ram[15194]), .B2(n3926), 
        .ZN(n19435) );
  MOAI22 U28341 ( .A1(n28529), .A2(n3925), .B1(ram[15195]), .B2(n3926), 
        .ZN(n19436) );
  MOAI22 U28342 ( .A1(n28294), .A2(n3925), .B1(ram[15196]), .B2(n3926), 
        .ZN(n19437) );
  MOAI22 U28343 ( .A1(n28059), .A2(n3925), .B1(ram[15197]), .B2(n3926), 
        .ZN(n19438) );
  MOAI22 U28344 ( .A1(n27824), .A2(n3925), .B1(ram[15198]), .B2(n3926), 
        .ZN(n19439) );
  MOAI22 U28345 ( .A1(n27589), .A2(n3925), .B1(ram[15199]), .B2(n3926), 
        .ZN(n19440) );
  MOAI22 U28346 ( .A1(n29234), .A2(n3927), .B1(ram[15200]), .B2(n3928), 
        .ZN(n19441) );
  MOAI22 U28347 ( .A1(n28999), .A2(n3927), .B1(ram[15201]), .B2(n3928), 
        .ZN(n19442) );
  MOAI22 U28348 ( .A1(n28764), .A2(n3927), .B1(ram[15202]), .B2(n3928), 
        .ZN(n19443) );
  MOAI22 U28349 ( .A1(n28529), .A2(n3927), .B1(ram[15203]), .B2(n3928), 
        .ZN(n19444) );
  MOAI22 U28350 ( .A1(n28294), .A2(n3927), .B1(ram[15204]), .B2(n3928), 
        .ZN(n19445) );
  MOAI22 U28351 ( .A1(n28059), .A2(n3927), .B1(ram[15205]), .B2(n3928), 
        .ZN(n19446) );
  MOAI22 U28352 ( .A1(n27824), .A2(n3927), .B1(ram[15206]), .B2(n3928), 
        .ZN(n19447) );
  MOAI22 U28353 ( .A1(n27589), .A2(n3927), .B1(ram[15207]), .B2(n3928), 
        .ZN(n19448) );
  MOAI22 U28354 ( .A1(n29234), .A2(n3929), .B1(ram[15208]), .B2(n3930), 
        .ZN(n19449) );
  MOAI22 U28355 ( .A1(n28999), .A2(n3929), .B1(ram[15209]), .B2(n3930), 
        .ZN(n19450) );
  MOAI22 U28356 ( .A1(n28764), .A2(n3929), .B1(ram[15210]), .B2(n3930), 
        .ZN(n19451) );
  MOAI22 U28357 ( .A1(n28529), .A2(n3929), .B1(ram[15211]), .B2(n3930), 
        .ZN(n19452) );
  MOAI22 U28358 ( .A1(n28294), .A2(n3929), .B1(ram[15212]), .B2(n3930), 
        .ZN(n19453) );
  MOAI22 U28359 ( .A1(n28059), .A2(n3929), .B1(ram[15213]), .B2(n3930), 
        .ZN(n19454) );
  MOAI22 U28360 ( .A1(n27824), .A2(n3929), .B1(ram[15214]), .B2(n3930), 
        .ZN(n19455) );
  MOAI22 U28361 ( .A1(n27589), .A2(n3929), .B1(ram[15215]), .B2(n3930), 
        .ZN(n19456) );
  MOAI22 U28362 ( .A1(n29234), .A2(n3931), .B1(ram[15216]), .B2(n3932), 
        .ZN(n19457) );
  MOAI22 U28363 ( .A1(n28999), .A2(n3931), .B1(ram[15217]), .B2(n3932), 
        .ZN(n19458) );
  MOAI22 U28364 ( .A1(n28764), .A2(n3931), .B1(ram[15218]), .B2(n3932), 
        .ZN(n19459) );
  MOAI22 U28365 ( .A1(n28529), .A2(n3931), .B1(ram[15219]), .B2(n3932), 
        .ZN(n19460) );
  MOAI22 U28366 ( .A1(n28294), .A2(n3931), .B1(ram[15220]), .B2(n3932), 
        .ZN(n19461) );
  MOAI22 U28367 ( .A1(n28059), .A2(n3931), .B1(ram[15221]), .B2(n3932), 
        .ZN(n19462) );
  MOAI22 U28368 ( .A1(n27824), .A2(n3931), .B1(ram[15222]), .B2(n3932), 
        .ZN(n19463) );
  MOAI22 U28369 ( .A1(n27589), .A2(n3931), .B1(ram[15223]), .B2(n3932), 
        .ZN(n19464) );
  MOAI22 U28370 ( .A1(n29234), .A2(n3933), .B1(ram[15224]), .B2(n3934), 
        .ZN(n19465) );
  MOAI22 U28371 ( .A1(n28999), .A2(n3933), .B1(ram[15225]), .B2(n3934), 
        .ZN(n19466) );
  MOAI22 U28372 ( .A1(n28764), .A2(n3933), .B1(ram[15226]), .B2(n3934), 
        .ZN(n19467) );
  MOAI22 U28373 ( .A1(n28529), .A2(n3933), .B1(ram[15227]), .B2(n3934), 
        .ZN(n19468) );
  MOAI22 U28374 ( .A1(n28294), .A2(n3933), .B1(ram[15228]), .B2(n3934), 
        .ZN(n19469) );
  MOAI22 U28375 ( .A1(n28059), .A2(n3933), .B1(ram[15229]), .B2(n3934), 
        .ZN(n19470) );
  MOAI22 U28376 ( .A1(n27824), .A2(n3933), .B1(ram[15230]), .B2(n3934), 
        .ZN(n19471) );
  MOAI22 U28377 ( .A1(n27589), .A2(n3933), .B1(ram[15231]), .B2(n3934), 
        .ZN(n19472) );
  MOAI22 U28378 ( .A1(n29234), .A2(n3935), .B1(ram[15232]), .B2(n3936), 
        .ZN(n19473) );
  MOAI22 U28379 ( .A1(n28999), .A2(n3935), .B1(ram[15233]), .B2(n3936), 
        .ZN(n19474) );
  MOAI22 U28380 ( .A1(n28764), .A2(n3935), .B1(ram[15234]), .B2(n3936), 
        .ZN(n19475) );
  MOAI22 U28381 ( .A1(n28529), .A2(n3935), .B1(ram[15235]), .B2(n3936), 
        .ZN(n19476) );
  MOAI22 U28382 ( .A1(n28294), .A2(n3935), .B1(ram[15236]), .B2(n3936), 
        .ZN(n19477) );
  MOAI22 U28383 ( .A1(n28059), .A2(n3935), .B1(ram[15237]), .B2(n3936), 
        .ZN(n19478) );
  MOAI22 U28384 ( .A1(n27824), .A2(n3935), .B1(ram[15238]), .B2(n3936), 
        .ZN(n19479) );
  MOAI22 U28385 ( .A1(n27589), .A2(n3935), .B1(ram[15239]), .B2(n3936), 
        .ZN(n19480) );
  MOAI22 U28386 ( .A1(n29234), .A2(n3937), .B1(ram[15240]), .B2(n3938), 
        .ZN(n19481) );
  MOAI22 U28387 ( .A1(n28999), .A2(n3937), .B1(ram[15241]), .B2(n3938), 
        .ZN(n19482) );
  MOAI22 U28388 ( .A1(n28764), .A2(n3937), .B1(ram[15242]), .B2(n3938), 
        .ZN(n19483) );
  MOAI22 U28389 ( .A1(n28529), .A2(n3937), .B1(ram[15243]), .B2(n3938), 
        .ZN(n19484) );
  MOAI22 U28390 ( .A1(n28294), .A2(n3937), .B1(ram[15244]), .B2(n3938), 
        .ZN(n19485) );
  MOAI22 U28391 ( .A1(n28059), .A2(n3937), .B1(ram[15245]), .B2(n3938), 
        .ZN(n19486) );
  MOAI22 U28392 ( .A1(n27824), .A2(n3937), .B1(ram[15246]), .B2(n3938), 
        .ZN(n19487) );
  MOAI22 U28393 ( .A1(n27589), .A2(n3937), .B1(ram[15247]), .B2(n3938), 
        .ZN(n19488) );
  MOAI22 U28394 ( .A1(n29234), .A2(n3939), .B1(ram[15248]), .B2(n3940), 
        .ZN(n19489) );
  MOAI22 U28395 ( .A1(n28999), .A2(n3939), .B1(ram[15249]), .B2(n3940), 
        .ZN(n19490) );
  MOAI22 U28396 ( .A1(n28764), .A2(n3939), .B1(ram[15250]), .B2(n3940), 
        .ZN(n19491) );
  MOAI22 U28397 ( .A1(n28529), .A2(n3939), .B1(ram[15251]), .B2(n3940), 
        .ZN(n19492) );
  MOAI22 U28398 ( .A1(n28294), .A2(n3939), .B1(ram[15252]), .B2(n3940), 
        .ZN(n19493) );
  MOAI22 U28399 ( .A1(n28059), .A2(n3939), .B1(ram[15253]), .B2(n3940), 
        .ZN(n19494) );
  MOAI22 U28400 ( .A1(n27824), .A2(n3939), .B1(ram[15254]), .B2(n3940), 
        .ZN(n19495) );
  MOAI22 U28401 ( .A1(n27589), .A2(n3939), .B1(ram[15255]), .B2(n3940), 
        .ZN(n19496) );
  MOAI22 U28402 ( .A1(n29234), .A2(n3941), .B1(ram[15256]), .B2(n3942), 
        .ZN(n19497) );
  MOAI22 U28403 ( .A1(n28999), .A2(n3941), .B1(ram[15257]), .B2(n3942), 
        .ZN(n19498) );
  MOAI22 U28404 ( .A1(n28764), .A2(n3941), .B1(ram[15258]), .B2(n3942), 
        .ZN(n19499) );
  MOAI22 U28405 ( .A1(n28529), .A2(n3941), .B1(ram[15259]), .B2(n3942), 
        .ZN(n19500) );
  MOAI22 U28406 ( .A1(n28294), .A2(n3941), .B1(ram[15260]), .B2(n3942), 
        .ZN(n19501) );
  MOAI22 U28407 ( .A1(n28059), .A2(n3941), .B1(ram[15261]), .B2(n3942), 
        .ZN(n19502) );
  MOAI22 U28408 ( .A1(n27824), .A2(n3941), .B1(ram[15262]), .B2(n3942), 
        .ZN(n19503) );
  MOAI22 U28409 ( .A1(n27589), .A2(n3941), .B1(ram[15263]), .B2(n3942), 
        .ZN(n19504) );
  MOAI22 U28410 ( .A1(n29234), .A2(n3943), .B1(ram[15264]), .B2(n3944), 
        .ZN(n19505) );
  MOAI22 U28411 ( .A1(n28999), .A2(n3943), .B1(ram[15265]), .B2(n3944), 
        .ZN(n19506) );
  MOAI22 U28412 ( .A1(n28764), .A2(n3943), .B1(ram[15266]), .B2(n3944), 
        .ZN(n19507) );
  MOAI22 U28413 ( .A1(n28529), .A2(n3943), .B1(ram[15267]), .B2(n3944), 
        .ZN(n19508) );
  MOAI22 U28414 ( .A1(n28294), .A2(n3943), .B1(ram[15268]), .B2(n3944), 
        .ZN(n19509) );
  MOAI22 U28415 ( .A1(n28059), .A2(n3943), .B1(ram[15269]), .B2(n3944), 
        .ZN(n19510) );
  MOAI22 U28416 ( .A1(n27824), .A2(n3943), .B1(ram[15270]), .B2(n3944), 
        .ZN(n19511) );
  MOAI22 U28417 ( .A1(n27589), .A2(n3943), .B1(ram[15271]), .B2(n3944), 
        .ZN(n19512) );
  MOAI22 U28418 ( .A1(n29234), .A2(n3945), .B1(ram[15272]), .B2(n3946), 
        .ZN(n19513) );
  MOAI22 U28419 ( .A1(n28999), .A2(n3945), .B1(ram[15273]), .B2(n3946), 
        .ZN(n19514) );
  MOAI22 U28420 ( .A1(n28764), .A2(n3945), .B1(ram[15274]), .B2(n3946), 
        .ZN(n19515) );
  MOAI22 U28421 ( .A1(n28529), .A2(n3945), .B1(ram[15275]), .B2(n3946), 
        .ZN(n19516) );
  MOAI22 U28422 ( .A1(n28294), .A2(n3945), .B1(ram[15276]), .B2(n3946), 
        .ZN(n19517) );
  MOAI22 U28423 ( .A1(n28059), .A2(n3945), .B1(ram[15277]), .B2(n3946), 
        .ZN(n19518) );
  MOAI22 U28424 ( .A1(n27824), .A2(n3945), .B1(ram[15278]), .B2(n3946), 
        .ZN(n19519) );
  MOAI22 U28425 ( .A1(n27589), .A2(n3945), .B1(ram[15279]), .B2(n3946), 
        .ZN(n19520) );
  MOAI22 U28426 ( .A1(n29234), .A2(n3947), .B1(ram[15280]), .B2(n3948), 
        .ZN(n19521) );
  MOAI22 U28427 ( .A1(n28999), .A2(n3947), .B1(ram[15281]), .B2(n3948), 
        .ZN(n19522) );
  MOAI22 U28428 ( .A1(n28764), .A2(n3947), .B1(ram[15282]), .B2(n3948), 
        .ZN(n19523) );
  MOAI22 U28429 ( .A1(n28529), .A2(n3947), .B1(ram[15283]), .B2(n3948), 
        .ZN(n19524) );
  MOAI22 U28430 ( .A1(n28294), .A2(n3947), .B1(ram[15284]), .B2(n3948), 
        .ZN(n19525) );
  MOAI22 U28431 ( .A1(n28059), .A2(n3947), .B1(ram[15285]), .B2(n3948), 
        .ZN(n19526) );
  MOAI22 U28432 ( .A1(n27824), .A2(n3947), .B1(ram[15286]), .B2(n3948), 
        .ZN(n19527) );
  MOAI22 U28433 ( .A1(n27589), .A2(n3947), .B1(ram[15287]), .B2(n3948), 
        .ZN(n19528) );
  MOAI22 U28434 ( .A1(n29235), .A2(n3949), .B1(ram[15288]), .B2(n3950), 
        .ZN(n19529) );
  MOAI22 U28435 ( .A1(n29000), .A2(n3949), .B1(ram[15289]), .B2(n3950), 
        .ZN(n19530) );
  MOAI22 U28436 ( .A1(n28765), .A2(n3949), .B1(ram[15290]), .B2(n3950), 
        .ZN(n19531) );
  MOAI22 U28437 ( .A1(n28530), .A2(n3949), .B1(ram[15291]), .B2(n3950), 
        .ZN(n19532) );
  MOAI22 U28438 ( .A1(n28295), .A2(n3949), .B1(ram[15292]), .B2(n3950), 
        .ZN(n19533) );
  MOAI22 U28439 ( .A1(n28060), .A2(n3949), .B1(ram[15293]), .B2(n3950), 
        .ZN(n19534) );
  MOAI22 U28440 ( .A1(n27825), .A2(n3949), .B1(ram[15294]), .B2(n3950), 
        .ZN(n19535) );
  MOAI22 U28441 ( .A1(n27590), .A2(n3949), .B1(ram[15295]), .B2(n3950), 
        .ZN(n19536) );
  MOAI22 U28442 ( .A1(n29235), .A2(n3951), .B1(ram[15296]), .B2(n3952), 
        .ZN(n19537) );
  MOAI22 U28443 ( .A1(n29000), .A2(n3951), .B1(ram[15297]), .B2(n3952), 
        .ZN(n19538) );
  MOAI22 U28444 ( .A1(n28765), .A2(n3951), .B1(ram[15298]), .B2(n3952), 
        .ZN(n19539) );
  MOAI22 U28445 ( .A1(n28530), .A2(n3951), .B1(ram[15299]), .B2(n3952), 
        .ZN(n19540) );
  MOAI22 U28446 ( .A1(n28295), .A2(n3951), .B1(ram[15300]), .B2(n3952), 
        .ZN(n19541) );
  MOAI22 U28447 ( .A1(n28060), .A2(n3951), .B1(ram[15301]), .B2(n3952), 
        .ZN(n19542) );
  MOAI22 U28448 ( .A1(n27825), .A2(n3951), .B1(ram[15302]), .B2(n3952), 
        .ZN(n19543) );
  MOAI22 U28449 ( .A1(n27590), .A2(n3951), .B1(ram[15303]), .B2(n3952), 
        .ZN(n19544) );
  MOAI22 U28450 ( .A1(n29235), .A2(n3953), .B1(ram[15304]), .B2(n3954), 
        .ZN(n19545) );
  MOAI22 U28451 ( .A1(n29000), .A2(n3953), .B1(ram[15305]), .B2(n3954), 
        .ZN(n19546) );
  MOAI22 U28452 ( .A1(n28765), .A2(n3953), .B1(ram[15306]), .B2(n3954), 
        .ZN(n19547) );
  MOAI22 U28453 ( .A1(n28530), .A2(n3953), .B1(ram[15307]), .B2(n3954), 
        .ZN(n19548) );
  MOAI22 U28454 ( .A1(n28295), .A2(n3953), .B1(ram[15308]), .B2(n3954), 
        .ZN(n19549) );
  MOAI22 U28455 ( .A1(n28060), .A2(n3953), .B1(ram[15309]), .B2(n3954), 
        .ZN(n19550) );
  MOAI22 U28456 ( .A1(n27825), .A2(n3953), .B1(ram[15310]), .B2(n3954), 
        .ZN(n19551) );
  MOAI22 U28457 ( .A1(n27590), .A2(n3953), .B1(ram[15311]), .B2(n3954), 
        .ZN(n19552) );
  MOAI22 U28458 ( .A1(n29235), .A2(n3955), .B1(ram[15312]), .B2(n3956), 
        .ZN(n19553) );
  MOAI22 U28459 ( .A1(n29000), .A2(n3955), .B1(ram[15313]), .B2(n3956), 
        .ZN(n19554) );
  MOAI22 U28460 ( .A1(n28765), .A2(n3955), .B1(ram[15314]), .B2(n3956), 
        .ZN(n19555) );
  MOAI22 U28461 ( .A1(n28530), .A2(n3955), .B1(ram[15315]), .B2(n3956), 
        .ZN(n19556) );
  MOAI22 U28462 ( .A1(n28295), .A2(n3955), .B1(ram[15316]), .B2(n3956), 
        .ZN(n19557) );
  MOAI22 U28463 ( .A1(n28060), .A2(n3955), .B1(ram[15317]), .B2(n3956), 
        .ZN(n19558) );
  MOAI22 U28464 ( .A1(n27825), .A2(n3955), .B1(ram[15318]), .B2(n3956), 
        .ZN(n19559) );
  MOAI22 U28465 ( .A1(n27590), .A2(n3955), .B1(ram[15319]), .B2(n3956), 
        .ZN(n19560) );
  MOAI22 U28466 ( .A1(n29235), .A2(n3957), .B1(ram[15320]), .B2(n3958), 
        .ZN(n19561) );
  MOAI22 U28467 ( .A1(n29000), .A2(n3957), .B1(ram[15321]), .B2(n3958), 
        .ZN(n19562) );
  MOAI22 U28468 ( .A1(n28765), .A2(n3957), .B1(ram[15322]), .B2(n3958), 
        .ZN(n19563) );
  MOAI22 U28469 ( .A1(n28530), .A2(n3957), .B1(ram[15323]), .B2(n3958), 
        .ZN(n19564) );
  MOAI22 U28470 ( .A1(n28295), .A2(n3957), .B1(ram[15324]), .B2(n3958), 
        .ZN(n19565) );
  MOAI22 U28471 ( .A1(n28060), .A2(n3957), .B1(ram[15325]), .B2(n3958), 
        .ZN(n19566) );
  MOAI22 U28472 ( .A1(n27825), .A2(n3957), .B1(ram[15326]), .B2(n3958), 
        .ZN(n19567) );
  MOAI22 U28473 ( .A1(n27590), .A2(n3957), .B1(ram[15327]), .B2(n3958), 
        .ZN(n19568) );
  MOAI22 U28474 ( .A1(n29235), .A2(n3959), .B1(ram[15328]), .B2(n3960), 
        .ZN(n19569) );
  MOAI22 U28475 ( .A1(n29000), .A2(n3959), .B1(ram[15329]), .B2(n3960), 
        .ZN(n19570) );
  MOAI22 U28476 ( .A1(n28765), .A2(n3959), .B1(ram[15330]), .B2(n3960), 
        .ZN(n19571) );
  MOAI22 U28477 ( .A1(n28530), .A2(n3959), .B1(ram[15331]), .B2(n3960), 
        .ZN(n19572) );
  MOAI22 U28478 ( .A1(n28295), .A2(n3959), .B1(ram[15332]), .B2(n3960), 
        .ZN(n19573) );
  MOAI22 U28479 ( .A1(n28060), .A2(n3959), .B1(ram[15333]), .B2(n3960), 
        .ZN(n19574) );
  MOAI22 U28480 ( .A1(n27825), .A2(n3959), .B1(ram[15334]), .B2(n3960), 
        .ZN(n19575) );
  MOAI22 U28481 ( .A1(n27590), .A2(n3959), .B1(ram[15335]), .B2(n3960), 
        .ZN(n19576) );
  MOAI22 U28482 ( .A1(n29235), .A2(n3961), .B1(ram[15336]), .B2(n3962), 
        .ZN(n19577) );
  MOAI22 U28483 ( .A1(n29000), .A2(n3961), .B1(ram[15337]), .B2(n3962), 
        .ZN(n19578) );
  MOAI22 U28484 ( .A1(n28765), .A2(n3961), .B1(ram[15338]), .B2(n3962), 
        .ZN(n19579) );
  MOAI22 U28485 ( .A1(n28530), .A2(n3961), .B1(ram[15339]), .B2(n3962), 
        .ZN(n19580) );
  MOAI22 U28486 ( .A1(n28295), .A2(n3961), .B1(ram[15340]), .B2(n3962), 
        .ZN(n19581) );
  MOAI22 U28487 ( .A1(n28060), .A2(n3961), .B1(ram[15341]), .B2(n3962), 
        .ZN(n19582) );
  MOAI22 U28488 ( .A1(n27825), .A2(n3961), .B1(ram[15342]), .B2(n3962), 
        .ZN(n19583) );
  MOAI22 U28489 ( .A1(n27590), .A2(n3961), .B1(ram[15343]), .B2(n3962), 
        .ZN(n19584) );
  MOAI22 U28490 ( .A1(n29235), .A2(n3963), .B1(ram[15344]), .B2(n3964), 
        .ZN(n19585) );
  MOAI22 U28491 ( .A1(n29000), .A2(n3963), .B1(ram[15345]), .B2(n3964), 
        .ZN(n19586) );
  MOAI22 U28492 ( .A1(n28765), .A2(n3963), .B1(ram[15346]), .B2(n3964), 
        .ZN(n19587) );
  MOAI22 U28493 ( .A1(n28530), .A2(n3963), .B1(ram[15347]), .B2(n3964), 
        .ZN(n19588) );
  MOAI22 U28494 ( .A1(n28295), .A2(n3963), .B1(ram[15348]), .B2(n3964), 
        .ZN(n19589) );
  MOAI22 U28495 ( .A1(n28060), .A2(n3963), .B1(ram[15349]), .B2(n3964), 
        .ZN(n19590) );
  MOAI22 U28496 ( .A1(n27825), .A2(n3963), .B1(ram[15350]), .B2(n3964), 
        .ZN(n19591) );
  MOAI22 U28497 ( .A1(n27590), .A2(n3963), .B1(ram[15351]), .B2(n3964), 
        .ZN(n19592) );
  MOAI22 U28498 ( .A1(n29235), .A2(n3965), .B1(ram[15352]), .B2(n3966), 
        .ZN(n19593) );
  MOAI22 U28499 ( .A1(n29000), .A2(n3965), .B1(ram[15353]), .B2(n3966), 
        .ZN(n19594) );
  MOAI22 U28500 ( .A1(n28765), .A2(n3965), .B1(ram[15354]), .B2(n3966), 
        .ZN(n19595) );
  MOAI22 U28501 ( .A1(n28530), .A2(n3965), .B1(ram[15355]), .B2(n3966), 
        .ZN(n19596) );
  MOAI22 U28502 ( .A1(n28295), .A2(n3965), .B1(ram[15356]), .B2(n3966), 
        .ZN(n19597) );
  MOAI22 U28503 ( .A1(n28060), .A2(n3965), .B1(ram[15357]), .B2(n3966), 
        .ZN(n19598) );
  MOAI22 U28504 ( .A1(n27825), .A2(n3965), .B1(ram[15358]), .B2(n3966), 
        .ZN(n19599) );
  MOAI22 U28505 ( .A1(n27590), .A2(n3965), .B1(ram[15359]), .B2(n3966), 
        .ZN(n19600) );
  MOAI22 U28506 ( .A1(n29235), .A2(n3967), .B1(ram[15360]), .B2(n3968), 
        .ZN(n19601) );
  MOAI22 U28507 ( .A1(n29000), .A2(n3967), .B1(ram[15361]), .B2(n3968), 
        .ZN(n19602) );
  MOAI22 U28508 ( .A1(n28765), .A2(n3967), .B1(ram[15362]), .B2(n3968), 
        .ZN(n19603) );
  MOAI22 U28509 ( .A1(n28530), .A2(n3967), .B1(ram[15363]), .B2(n3968), 
        .ZN(n19604) );
  MOAI22 U28510 ( .A1(n28295), .A2(n3967), .B1(ram[15364]), .B2(n3968), 
        .ZN(n19605) );
  MOAI22 U28511 ( .A1(n28060), .A2(n3967), .B1(ram[15365]), .B2(n3968), 
        .ZN(n19606) );
  MOAI22 U28512 ( .A1(n27825), .A2(n3967), .B1(ram[15366]), .B2(n3968), 
        .ZN(n19607) );
  MOAI22 U28513 ( .A1(n27590), .A2(n3967), .B1(ram[15367]), .B2(n3968), 
        .ZN(n19608) );
  MOAI22 U28514 ( .A1(n29235), .A2(n3970), .B1(ram[15368]), .B2(n3971), 
        .ZN(n19609) );
  MOAI22 U28515 ( .A1(n29000), .A2(n3970), .B1(ram[15369]), .B2(n3971), 
        .ZN(n19610) );
  MOAI22 U28516 ( .A1(n28765), .A2(n3970), .B1(ram[15370]), .B2(n3971), 
        .ZN(n19611) );
  MOAI22 U28517 ( .A1(n28530), .A2(n3970), .B1(ram[15371]), .B2(n3971), 
        .ZN(n19612) );
  MOAI22 U28518 ( .A1(n28295), .A2(n3970), .B1(ram[15372]), .B2(n3971), 
        .ZN(n19613) );
  MOAI22 U28519 ( .A1(n28060), .A2(n3970), .B1(ram[15373]), .B2(n3971), 
        .ZN(n19614) );
  MOAI22 U28520 ( .A1(n27825), .A2(n3970), .B1(ram[15374]), .B2(n3971), 
        .ZN(n19615) );
  MOAI22 U28521 ( .A1(n27590), .A2(n3970), .B1(ram[15375]), .B2(n3971), 
        .ZN(n19616) );
  MOAI22 U28522 ( .A1(n29235), .A2(n3972), .B1(ram[15376]), .B2(n3973), 
        .ZN(n19617) );
  MOAI22 U28523 ( .A1(n29000), .A2(n3972), .B1(ram[15377]), .B2(n3973), 
        .ZN(n19618) );
  MOAI22 U28524 ( .A1(n28765), .A2(n3972), .B1(ram[15378]), .B2(n3973), 
        .ZN(n19619) );
  MOAI22 U28525 ( .A1(n28530), .A2(n3972), .B1(ram[15379]), .B2(n3973), 
        .ZN(n19620) );
  MOAI22 U28526 ( .A1(n28295), .A2(n3972), .B1(ram[15380]), .B2(n3973), 
        .ZN(n19621) );
  MOAI22 U28527 ( .A1(n28060), .A2(n3972), .B1(ram[15381]), .B2(n3973), 
        .ZN(n19622) );
  MOAI22 U28528 ( .A1(n27825), .A2(n3972), .B1(ram[15382]), .B2(n3973), 
        .ZN(n19623) );
  MOAI22 U28529 ( .A1(n27590), .A2(n3972), .B1(ram[15383]), .B2(n3973), 
        .ZN(n19624) );
  MOAI22 U28530 ( .A1(n29235), .A2(n3974), .B1(ram[15384]), .B2(n3975), 
        .ZN(n19625) );
  MOAI22 U28531 ( .A1(n29000), .A2(n3974), .B1(ram[15385]), .B2(n3975), 
        .ZN(n19626) );
  MOAI22 U28532 ( .A1(n28765), .A2(n3974), .B1(ram[15386]), .B2(n3975), 
        .ZN(n19627) );
  MOAI22 U28533 ( .A1(n28530), .A2(n3974), .B1(ram[15387]), .B2(n3975), 
        .ZN(n19628) );
  MOAI22 U28534 ( .A1(n28295), .A2(n3974), .B1(ram[15388]), .B2(n3975), 
        .ZN(n19629) );
  MOAI22 U28535 ( .A1(n28060), .A2(n3974), .B1(ram[15389]), .B2(n3975), 
        .ZN(n19630) );
  MOAI22 U28536 ( .A1(n27825), .A2(n3974), .B1(ram[15390]), .B2(n3975), 
        .ZN(n19631) );
  MOAI22 U28537 ( .A1(n27590), .A2(n3974), .B1(ram[15391]), .B2(n3975), 
        .ZN(n19632) );
  MOAI22 U28538 ( .A1(n29236), .A2(n3976), .B1(ram[15392]), .B2(n3977), 
        .ZN(n19633) );
  MOAI22 U28539 ( .A1(n29001), .A2(n3976), .B1(ram[15393]), .B2(n3977), 
        .ZN(n19634) );
  MOAI22 U28540 ( .A1(n28766), .A2(n3976), .B1(ram[15394]), .B2(n3977), 
        .ZN(n19635) );
  MOAI22 U28541 ( .A1(n28531), .A2(n3976), .B1(ram[15395]), .B2(n3977), 
        .ZN(n19636) );
  MOAI22 U28542 ( .A1(n28296), .A2(n3976), .B1(ram[15396]), .B2(n3977), 
        .ZN(n19637) );
  MOAI22 U28543 ( .A1(n28061), .A2(n3976), .B1(ram[15397]), .B2(n3977), 
        .ZN(n19638) );
  MOAI22 U28544 ( .A1(n27826), .A2(n3976), .B1(ram[15398]), .B2(n3977), 
        .ZN(n19639) );
  MOAI22 U28545 ( .A1(n27591), .A2(n3976), .B1(ram[15399]), .B2(n3977), 
        .ZN(n19640) );
  MOAI22 U28546 ( .A1(n29236), .A2(n3978), .B1(ram[15400]), .B2(n3979), 
        .ZN(n19641) );
  MOAI22 U28547 ( .A1(n29001), .A2(n3978), .B1(ram[15401]), .B2(n3979), 
        .ZN(n19642) );
  MOAI22 U28548 ( .A1(n28766), .A2(n3978), .B1(ram[15402]), .B2(n3979), 
        .ZN(n19643) );
  MOAI22 U28549 ( .A1(n28531), .A2(n3978), .B1(ram[15403]), .B2(n3979), 
        .ZN(n19644) );
  MOAI22 U28550 ( .A1(n28296), .A2(n3978), .B1(ram[15404]), .B2(n3979), 
        .ZN(n19645) );
  MOAI22 U28551 ( .A1(n28061), .A2(n3978), .B1(ram[15405]), .B2(n3979), 
        .ZN(n19646) );
  MOAI22 U28552 ( .A1(n27826), .A2(n3978), .B1(ram[15406]), .B2(n3979), 
        .ZN(n19647) );
  MOAI22 U28553 ( .A1(n27591), .A2(n3978), .B1(ram[15407]), .B2(n3979), 
        .ZN(n19648) );
  MOAI22 U28554 ( .A1(n29236), .A2(n3980), .B1(ram[15408]), .B2(n3981), 
        .ZN(n19649) );
  MOAI22 U28555 ( .A1(n29001), .A2(n3980), .B1(ram[15409]), .B2(n3981), 
        .ZN(n19650) );
  MOAI22 U28556 ( .A1(n28766), .A2(n3980), .B1(ram[15410]), .B2(n3981), 
        .ZN(n19651) );
  MOAI22 U28557 ( .A1(n28531), .A2(n3980), .B1(ram[15411]), .B2(n3981), 
        .ZN(n19652) );
  MOAI22 U28558 ( .A1(n28296), .A2(n3980), .B1(ram[15412]), .B2(n3981), 
        .ZN(n19653) );
  MOAI22 U28559 ( .A1(n28061), .A2(n3980), .B1(ram[15413]), .B2(n3981), 
        .ZN(n19654) );
  MOAI22 U28560 ( .A1(n27826), .A2(n3980), .B1(ram[15414]), .B2(n3981), 
        .ZN(n19655) );
  MOAI22 U28561 ( .A1(n27591), .A2(n3980), .B1(ram[15415]), .B2(n3981), 
        .ZN(n19656) );
  MOAI22 U28562 ( .A1(n29236), .A2(n3982), .B1(ram[15416]), .B2(n3983), 
        .ZN(n19657) );
  MOAI22 U28563 ( .A1(n29001), .A2(n3982), .B1(ram[15417]), .B2(n3983), 
        .ZN(n19658) );
  MOAI22 U28564 ( .A1(n28766), .A2(n3982), .B1(ram[15418]), .B2(n3983), 
        .ZN(n19659) );
  MOAI22 U28565 ( .A1(n28531), .A2(n3982), .B1(ram[15419]), .B2(n3983), 
        .ZN(n19660) );
  MOAI22 U28566 ( .A1(n28296), .A2(n3982), .B1(ram[15420]), .B2(n3983), 
        .ZN(n19661) );
  MOAI22 U28567 ( .A1(n28061), .A2(n3982), .B1(ram[15421]), .B2(n3983), 
        .ZN(n19662) );
  MOAI22 U28568 ( .A1(n27826), .A2(n3982), .B1(ram[15422]), .B2(n3983), 
        .ZN(n19663) );
  MOAI22 U28569 ( .A1(n27591), .A2(n3982), .B1(ram[15423]), .B2(n3983), 
        .ZN(n19664) );
  MOAI22 U28570 ( .A1(n29236), .A2(n3984), .B1(ram[15424]), .B2(n3985), 
        .ZN(n19665) );
  MOAI22 U28571 ( .A1(n29001), .A2(n3984), .B1(ram[15425]), .B2(n3985), 
        .ZN(n19666) );
  MOAI22 U28572 ( .A1(n28766), .A2(n3984), .B1(ram[15426]), .B2(n3985), 
        .ZN(n19667) );
  MOAI22 U28573 ( .A1(n28531), .A2(n3984), .B1(ram[15427]), .B2(n3985), 
        .ZN(n19668) );
  MOAI22 U28574 ( .A1(n28296), .A2(n3984), .B1(ram[15428]), .B2(n3985), 
        .ZN(n19669) );
  MOAI22 U28575 ( .A1(n28061), .A2(n3984), .B1(ram[15429]), .B2(n3985), 
        .ZN(n19670) );
  MOAI22 U28576 ( .A1(n27826), .A2(n3984), .B1(ram[15430]), .B2(n3985), 
        .ZN(n19671) );
  MOAI22 U28577 ( .A1(n27591), .A2(n3984), .B1(ram[15431]), .B2(n3985), 
        .ZN(n19672) );
  MOAI22 U28578 ( .A1(n29236), .A2(n3986), .B1(ram[15432]), .B2(n3987), 
        .ZN(n19673) );
  MOAI22 U28579 ( .A1(n29001), .A2(n3986), .B1(ram[15433]), .B2(n3987), 
        .ZN(n19674) );
  MOAI22 U28580 ( .A1(n28766), .A2(n3986), .B1(ram[15434]), .B2(n3987), 
        .ZN(n19675) );
  MOAI22 U28581 ( .A1(n28531), .A2(n3986), .B1(ram[15435]), .B2(n3987), 
        .ZN(n19676) );
  MOAI22 U28582 ( .A1(n28296), .A2(n3986), .B1(ram[15436]), .B2(n3987), 
        .ZN(n19677) );
  MOAI22 U28583 ( .A1(n28061), .A2(n3986), .B1(ram[15437]), .B2(n3987), 
        .ZN(n19678) );
  MOAI22 U28584 ( .A1(n27826), .A2(n3986), .B1(ram[15438]), .B2(n3987), 
        .ZN(n19679) );
  MOAI22 U28585 ( .A1(n27591), .A2(n3986), .B1(ram[15439]), .B2(n3987), 
        .ZN(n19680) );
  MOAI22 U28586 ( .A1(n29236), .A2(n3988), .B1(ram[15440]), .B2(n3989), 
        .ZN(n19681) );
  MOAI22 U28587 ( .A1(n29001), .A2(n3988), .B1(ram[15441]), .B2(n3989), 
        .ZN(n19682) );
  MOAI22 U28588 ( .A1(n28766), .A2(n3988), .B1(ram[15442]), .B2(n3989), 
        .ZN(n19683) );
  MOAI22 U28589 ( .A1(n28531), .A2(n3988), .B1(ram[15443]), .B2(n3989), 
        .ZN(n19684) );
  MOAI22 U28590 ( .A1(n28296), .A2(n3988), .B1(ram[15444]), .B2(n3989), 
        .ZN(n19685) );
  MOAI22 U28591 ( .A1(n28061), .A2(n3988), .B1(ram[15445]), .B2(n3989), 
        .ZN(n19686) );
  MOAI22 U28592 ( .A1(n27826), .A2(n3988), .B1(ram[15446]), .B2(n3989), 
        .ZN(n19687) );
  MOAI22 U28593 ( .A1(n27591), .A2(n3988), .B1(ram[15447]), .B2(n3989), 
        .ZN(n19688) );
  MOAI22 U28594 ( .A1(n29236), .A2(n3990), .B1(ram[15448]), .B2(n3991), 
        .ZN(n19689) );
  MOAI22 U28595 ( .A1(n29001), .A2(n3990), .B1(ram[15449]), .B2(n3991), 
        .ZN(n19690) );
  MOAI22 U28596 ( .A1(n28766), .A2(n3990), .B1(ram[15450]), .B2(n3991), 
        .ZN(n19691) );
  MOAI22 U28597 ( .A1(n28531), .A2(n3990), .B1(ram[15451]), .B2(n3991), 
        .ZN(n19692) );
  MOAI22 U28598 ( .A1(n28296), .A2(n3990), .B1(ram[15452]), .B2(n3991), 
        .ZN(n19693) );
  MOAI22 U28599 ( .A1(n28061), .A2(n3990), .B1(ram[15453]), .B2(n3991), 
        .ZN(n19694) );
  MOAI22 U28600 ( .A1(n27826), .A2(n3990), .B1(ram[15454]), .B2(n3991), 
        .ZN(n19695) );
  MOAI22 U28601 ( .A1(n27591), .A2(n3990), .B1(ram[15455]), .B2(n3991), 
        .ZN(n19696) );
  MOAI22 U28602 ( .A1(n29236), .A2(n3992), .B1(ram[15456]), .B2(n3993), 
        .ZN(n19697) );
  MOAI22 U28603 ( .A1(n29001), .A2(n3992), .B1(ram[15457]), .B2(n3993), 
        .ZN(n19698) );
  MOAI22 U28604 ( .A1(n28766), .A2(n3992), .B1(ram[15458]), .B2(n3993), 
        .ZN(n19699) );
  MOAI22 U28605 ( .A1(n28531), .A2(n3992), .B1(ram[15459]), .B2(n3993), 
        .ZN(n19700) );
  MOAI22 U28606 ( .A1(n28296), .A2(n3992), .B1(ram[15460]), .B2(n3993), 
        .ZN(n19701) );
  MOAI22 U28607 ( .A1(n28061), .A2(n3992), .B1(ram[15461]), .B2(n3993), 
        .ZN(n19702) );
  MOAI22 U28608 ( .A1(n27826), .A2(n3992), .B1(ram[15462]), .B2(n3993), 
        .ZN(n19703) );
  MOAI22 U28609 ( .A1(n27591), .A2(n3992), .B1(ram[15463]), .B2(n3993), 
        .ZN(n19704) );
  MOAI22 U28610 ( .A1(n29236), .A2(n3994), .B1(ram[15464]), .B2(n3995), 
        .ZN(n19705) );
  MOAI22 U28611 ( .A1(n29001), .A2(n3994), .B1(ram[15465]), .B2(n3995), 
        .ZN(n19706) );
  MOAI22 U28612 ( .A1(n28766), .A2(n3994), .B1(ram[15466]), .B2(n3995), 
        .ZN(n19707) );
  MOAI22 U28613 ( .A1(n28531), .A2(n3994), .B1(ram[15467]), .B2(n3995), 
        .ZN(n19708) );
  MOAI22 U28614 ( .A1(n28296), .A2(n3994), .B1(ram[15468]), .B2(n3995), 
        .ZN(n19709) );
  MOAI22 U28615 ( .A1(n28061), .A2(n3994), .B1(ram[15469]), .B2(n3995), 
        .ZN(n19710) );
  MOAI22 U28616 ( .A1(n27826), .A2(n3994), .B1(ram[15470]), .B2(n3995), 
        .ZN(n19711) );
  MOAI22 U28617 ( .A1(n27591), .A2(n3994), .B1(ram[15471]), .B2(n3995), 
        .ZN(n19712) );
  MOAI22 U28618 ( .A1(n29236), .A2(n3996), .B1(ram[15472]), .B2(n3997), 
        .ZN(n19713) );
  MOAI22 U28619 ( .A1(n29001), .A2(n3996), .B1(ram[15473]), .B2(n3997), 
        .ZN(n19714) );
  MOAI22 U28620 ( .A1(n28766), .A2(n3996), .B1(ram[15474]), .B2(n3997), 
        .ZN(n19715) );
  MOAI22 U28621 ( .A1(n28531), .A2(n3996), .B1(ram[15475]), .B2(n3997), 
        .ZN(n19716) );
  MOAI22 U28622 ( .A1(n28296), .A2(n3996), .B1(ram[15476]), .B2(n3997), 
        .ZN(n19717) );
  MOAI22 U28623 ( .A1(n28061), .A2(n3996), .B1(ram[15477]), .B2(n3997), 
        .ZN(n19718) );
  MOAI22 U28624 ( .A1(n27826), .A2(n3996), .B1(ram[15478]), .B2(n3997), 
        .ZN(n19719) );
  MOAI22 U28625 ( .A1(n27591), .A2(n3996), .B1(ram[15479]), .B2(n3997), 
        .ZN(n19720) );
  MOAI22 U28626 ( .A1(n29236), .A2(n3998), .B1(ram[15480]), .B2(n3999), 
        .ZN(n19721) );
  MOAI22 U28627 ( .A1(n29001), .A2(n3998), .B1(ram[15481]), .B2(n3999), 
        .ZN(n19722) );
  MOAI22 U28628 ( .A1(n28766), .A2(n3998), .B1(ram[15482]), .B2(n3999), 
        .ZN(n19723) );
  MOAI22 U28629 ( .A1(n28531), .A2(n3998), .B1(ram[15483]), .B2(n3999), 
        .ZN(n19724) );
  MOAI22 U28630 ( .A1(n28296), .A2(n3998), .B1(ram[15484]), .B2(n3999), 
        .ZN(n19725) );
  MOAI22 U28631 ( .A1(n28061), .A2(n3998), .B1(ram[15485]), .B2(n3999), 
        .ZN(n19726) );
  MOAI22 U28632 ( .A1(n27826), .A2(n3998), .B1(ram[15486]), .B2(n3999), 
        .ZN(n19727) );
  MOAI22 U28633 ( .A1(n27591), .A2(n3998), .B1(ram[15487]), .B2(n3999), 
        .ZN(n19728) );
  MOAI22 U28634 ( .A1(n29236), .A2(n4000), .B1(ram[15488]), .B2(n4001), 
        .ZN(n19729) );
  MOAI22 U28635 ( .A1(n29001), .A2(n4000), .B1(ram[15489]), .B2(n4001), 
        .ZN(n19730) );
  MOAI22 U28636 ( .A1(n28766), .A2(n4000), .B1(ram[15490]), .B2(n4001), 
        .ZN(n19731) );
  MOAI22 U28637 ( .A1(n28531), .A2(n4000), .B1(ram[15491]), .B2(n4001), 
        .ZN(n19732) );
  MOAI22 U28638 ( .A1(n28296), .A2(n4000), .B1(ram[15492]), .B2(n4001), 
        .ZN(n19733) );
  MOAI22 U28639 ( .A1(n28061), .A2(n4000), .B1(ram[15493]), .B2(n4001), 
        .ZN(n19734) );
  MOAI22 U28640 ( .A1(n27826), .A2(n4000), .B1(ram[15494]), .B2(n4001), 
        .ZN(n19735) );
  MOAI22 U28641 ( .A1(n27591), .A2(n4000), .B1(ram[15495]), .B2(n4001), 
        .ZN(n19736) );
  MOAI22 U28642 ( .A1(n29237), .A2(n4002), .B1(ram[15496]), .B2(n4003), 
        .ZN(n19737) );
  MOAI22 U28643 ( .A1(n29002), .A2(n4002), .B1(ram[15497]), .B2(n4003), 
        .ZN(n19738) );
  MOAI22 U28644 ( .A1(n28767), .A2(n4002), .B1(ram[15498]), .B2(n4003), 
        .ZN(n19739) );
  MOAI22 U28645 ( .A1(n28532), .A2(n4002), .B1(ram[15499]), .B2(n4003), 
        .ZN(n19740) );
  MOAI22 U28646 ( .A1(n28297), .A2(n4002), .B1(ram[15500]), .B2(n4003), 
        .ZN(n19741) );
  MOAI22 U28647 ( .A1(n28062), .A2(n4002), .B1(ram[15501]), .B2(n4003), 
        .ZN(n19742) );
  MOAI22 U28648 ( .A1(n27827), .A2(n4002), .B1(ram[15502]), .B2(n4003), 
        .ZN(n19743) );
  MOAI22 U28649 ( .A1(n27592), .A2(n4002), .B1(ram[15503]), .B2(n4003), 
        .ZN(n19744) );
  MOAI22 U28650 ( .A1(n29237), .A2(n4004), .B1(ram[15504]), .B2(n4005), 
        .ZN(n19745) );
  MOAI22 U28651 ( .A1(n29002), .A2(n4004), .B1(ram[15505]), .B2(n4005), 
        .ZN(n19746) );
  MOAI22 U28652 ( .A1(n28767), .A2(n4004), .B1(ram[15506]), .B2(n4005), 
        .ZN(n19747) );
  MOAI22 U28653 ( .A1(n28532), .A2(n4004), .B1(ram[15507]), .B2(n4005), 
        .ZN(n19748) );
  MOAI22 U28654 ( .A1(n28297), .A2(n4004), .B1(ram[15508]), .B2(n4005), 
        .ZN(n19749) );
  MOAI22 U28655 ( .A1(n28062), .A2(n4004), .B1(ram[15509]), .B2(n4005), 
        .ZN(n19750) );
  MOAI22 U28656 ( .A1(n27827), .A2(n4004), .B1(ram[15510]), .B2(n4005), 
        .ZN(n19751) );
  MOAI22 U28657 ( .A1(n27592), .A2(n4004), .B1(ram[15511]), .B2(n4005), 
        .ZN(n19752) );
  MOAI22 U28658 ( .A1(n29237), .A2(n4006), .B1(ram[15512]), .B2(n4007), 
        .ZN(n19753) );
  MOAI22 U28659 ( .A1(n29002), .A2(n4006), .B1(ram[15513]), .B2(n4007), 
        .ZN(n19754) );
  MOAI22 U28660 ( .A1(n28767), .A2(n4006), .B1(ram[15514]), .B2(n4007), 
        .ZN(n19755) );
  MOAI22 U28661 ( .A1(n28532), .A2(n4006), .B1(ram[15515]), .B2(n4007), 
        .ZN(n19756) );
  MOAI22 U28662 ( .A1(n28297), .A2(n4006), .B1(ram[15516]), .B2(n4007), 
        .ZN(n19757) );
  MOAI22 U28663 ( .A1(n28062), .A2(n4006), .B1(ram[15517]), .B2(n4007), 
        .ZN(n19758) );
  MOAI22 U28664 ( .A1(n27827), .A2(n4006), .B1(ram[15518]), .B2(n4007), 
        .ZN(n19759) );
  MOAI22 U28665 ( .A1(n27592), .A2(n4006), .B1(ram[15519]), .B2(n4007), 
        .ZN(n19760) );
  MOAI22 U28666 ( .A1(n29237), .A2(n4008), .B1(ram[15520]), .B2(n4009), 
        .ZN(n19761) );
  MOAI22 U28667 ( .A1(n29002), .A2(n4008), .B1(ram[15521]), .B2(n4009), 
        .ZN(n19762) );
  MOAI22 U28668 ( .A1(n28767), .A2(n4008), .B1(ram[15522]), .B2(n4009), 
        .ZN(n19763) );
  MOAI22 U28669 ( .A1(n28532), .A2(n4008), .B1(ram[15523]), .B2(n4009), 
        .ZN(n19764) );
  MOAI22 U28670 ( .A1(n28297), .A2(n4008), .B1(ram[15524]), .B2(n4009), 
        .ZN(n19765) );
  MOAI22 U28671 ( .A1(n28062), .A2(n4008), .B1(ram[15525]), .B2(n4009), 
        .ZN(n19766) );
  MOAI22 U28672 ( .A1(n27827), .A2(n4008), .B1(ram[15526]), .B2(n4009), 
        .ZN(n19767) );
  MOAI22 U28673 ( .A1(n27592), .A2(n4008), .B1(ram[15527]), .B2(n4009), 
        .ZN(n19768) );
  MOAI22 U28674 ( .A1(n29237), .A2(n4010), .B1(ram[15528]), .B2(n4011), 
        .ZN(n19769) );
  MOAI22 U28675 ( .A1(n29002), .A2(n4010), .B1(ram[15529]), .B2(n4011), 
        .ZN(n19770) );
  MOAI22 U28676 ( .A1(n28767), .A2(n4010), .B1(ram[15530]), .B2(n4011), 
        .ZN(n19771) );
  MOAI22 U28677 ( .A1(n28532), .A2(n4010), .B1(ram[15531]), .B2(n4011), 
        .ZN(n19772) );
  MOAI22 U28678 ( .A1(n28297), .A2(n4010), .B1(ram[15532]), .B2(n4011), 
        .ZN(n19773) );
  MOAI22 U28679 ( .A1(n28062), .A2(n4010), .B1(ram[15533]), .B2(n4011), 
        .ZN(n19774) );
  MOAI22 U28680 ( .A1(n27827), .A2(n4010), .B1(ram[15534]), .B2(n4011), 
        .ZN(n19775) );
  MOAI22 U28681 ( .A1(n27592), .A2(n4010), .B1(ram[15535]), .B2(n4011), 
        .ZN(n19776) );
  MOAI22 U28682 ( .A1(n29237), .A2(n4012), .B1(ram[15536]), .B2(n4013), 
        .ZN(n19777) );
  MOAI22 U28683 ( .A1(n29002), .A2(n4012), .B1(ram[15537]), .B2(n4013), 
        .ZN(n19778) );
  MOAI22 U28684 ( .A1(n28767), .A2(n4012), .B1(ram[15538]), .B2(n4013), 
        .ZN(n19779) );
  MOAI22 U28685 ( .A1(n28532), .A2(n4012), .B1(ram[15539]), .B2(n4013), 
        .ZN(n19780) );
  MOAI22 U28686 ( .A1(n28297), .A2(n4012), .B1(ram[15540]), .B2(n4013), 
        .ZN(n19781) );
  MOAI22 U28687 ( .A1(n28062), .A2(n4012), .B1(ram[15541]), .B2(n4013), 
        .ZN(n19782) );
  MOAI22 U28688 ( .A1(n27827), .A2(n4012), .B1(ram[15542]), .B2(n4013), 
        .ZN(n19783) );
  MOAI22 U28689 ( .A1(n27592), .A2(n4012), .B1(ram[15543]), .B2(n4013), 
        .ZN(n19784) );
  MOAI22 U28690 ( .A1(n29237), .A2(n4014), .B1(ram[15544]), .B2(n4015), 
        .ZN(n19785) );
  MOAI22 U28691 ( .A1(n29002), .A2(n4014), .B1(ram[15545]), .B2(n4015), 
        .ZN(n19786) );
  MOAI22 U28692 ( .A1(n28767), .A2(n4014), .B1(ram[15546]), .B2(n4015), 
        .ZN(n19787) );
  MOAI22 U28693 ( .A1(n28532), .A2(n4014), .B1(ram[15547]), .B2(n4015), 
        .ZN(n19788) );
  MOAI22 U28694 ( .A1(n28297), .A2(n4014), .B1(ram[15548]), .B2(n4015), 
        .ZN(n19789) );
  MOAI22 U28695 ( .A1(n28062), .A2(n4014), .B1(ram[15549]), .B2(n4015), 
        .ZN(n19790) );
  MOAI22 U28696 ( .A1(n27827), .A2(n4014), .B1(ram[15550]), .B2(n4015), 
        .ZN(n19791) );
  MOAI22 U28697 ( .A1(n27592), .A2(n4014), .B1(ram[15551]), .B2(n4015), 
        .ZN(n19792) );
  MOAI22 U28698 ( .A1(n29237), .A2(n4016), .B1(ram[15552]), .B2(n4017), 
        .ZN(n19793) );
  MOAI22 U28699 ( .A1(n29002), .A2(n4016), .B1(ram[15553]), .B2(n4017), 
        .ZN(n19794) );
  MOAI22 U28700 ( .A1(n28767), .A2(n4016), .B1(ram[15554]), .B2(n4017), 
        .ZN(n19795) );
  MOAI22 U28701 ( .A1(n28532), .A2(n4016), .B1(ram[15555]), .B2(n4017), 
        .ZN(n19796) );
  MOAI22 U28702 ( .A1(n28297), .A2(n4016), .B1(ram[15556]), .B2(n4017), 
        .ZN(n19797) );
  MOAI22 U28703 ( .A1(n28062), .A2(n4016), .B1(ram[15557]), .B2(n4017), 
        .ZN(n19798) );
  MOAI22 U28704 ( .A1(n27827), .A2(n4016), .B1(ram[15558]), .B2(n4017), 
        .ZN(n19799) );
  MOAI22 U28705 ( .A1(n27592), .A2(n4016), .B1(ram[15559]), .B2(n4017), 
        .ZN(n19800) );
  MOAI22 U28706 ( .A1(n29237), .A2(n4018), .B1(ram[15560]), .B2(n4019), 
        .ZN(n19801) );
  MOAI22 U28707 ( .A1(n29002), .A2(n4018), .B1(ram[15561]), .B2(n4019), 
        .ZN(n19802) );
  MOAI22 U28708 ( .A1(n28767), .A2(n4018), .B1(ram[15562]), .B2(n4019), 
        .ZN(n19803) );
  MOAI22 U28709 ( .A1(n28532), .A2(n4018), .B1(ram[15563]), .B2(n4019), 
        .ZN(n19804) );
  MOAI22 U28710 ( .A1(n28297), .A2(n4018), .B1(ram[15564]), .B2(n4019), 
        .ZN(n19805) );
  MOAI22 U28711 ( .A1(n28062), .A2(n4018), .B1(ram[15565]), .B2(n4019), 
        .ZN(n19806) );
  MOAI22 U28712 ( .A1(n27827), .A2(n4018), .B1(ram[15566]), .B2(n4019), 
        .ZN(n19807) );
  MOAI22 U28713 ( .A1(n27592), .A2(n4018), .B1(ram[15567]), .B2(n4019), 
        .ZN(n19808) );
  MOAI22 U28714 ( .A1(n29237), .A2(n4020), .B1(ram[15568]), .B2(n4021), 
        .ZN(n19809) );
  MOAI22 U28715 ( .A1(n29002), .A2(n4020), .B1(ram[15569]), .B2(n4021), 
        .ZN(n19810) );
  MOAI22 U28716 ( .A1(n28767), .A2(n4020), .B1(ram[15570]), .B2(n4021), 
        .ZN(n19811) );
  MOAI22 U28717 ( .A1(n28532), .A2(n4020), .B1(ram[15571]), .B2(n4021), 
        .ZN(n19812) );
  MOAI22 U28718 ( .A1(n28297), .A2(n4020), .B1(ram[15572]), .B2(n4021), 
        .ZN(n19813) );
  MOAI22 U28719 ( .A1(n28062), .A2(n4020), .B1(ram[15573]), .B2(n4021), 
        .ZN(n19814) );
  MOAI22 U28720 ( .A1(n27827), .A2(n4020), .B1(ram[15574]), .B2(n4021), 
        .ZN(n19815) );
  MOAI22 U28721 ( .A1(n27592), .A2(n4020), .B1(ram[15575]), .B2(n4021), 
        .ZN(n19816) );
  MOAI22 U28722 ( .A1(n29237), .A2(n4022), .B1(ram[15576]), .B2(n4023), 
        .ZN(n19817) );
  MOAI22 U28723 ( .A1(n29002), .A2(n4022), .B1(ram[15577]), .B2(n4023), 
        .ZN(n19818) );
  MOAI22 U28724 ( .A1(n28767), .A2(n4022), .B1(ram[15578]), .B2(n4023), 
        .ZN(n19819) );
  MOAI22 U28725 ( .A1(n28532), .A2(n4022), .B1(ram[15579]), .B2(n4023), 
        .ZN(n19820) );
  MOAI22 U28726 ( .A1(n28297), .A2(n4022), .B1(ram[15580]), .B2(n4023), 
        .ZN(n19821) );
  MOAI22 U28727 ( .A1(n28062), .A2(n4022), .B1(ram[15581]), .B2(n4023), 
        .ZN(n19822) );
  MOAI22 U28728 ( .A1(n27827), .A2(n4022), .B1(ram[15582]), .B2(n4023), 
        .ZN(n19823) );
  MOAI22 U28729 ( .A1(n27592), .A2(n4022), .B1(ram[15583]), .B2(n4023), 
        .ZN(n19824) );
  MOAI22 U28730 ( .A1(n29237), .A2(n4024), .B1(ram[15584]), .B2(n4025), 
        .ZN(n19825) );
  MOAI22 U28731 ( .A1(n29002), .A2(n4024), .B1(ram[15585]), .B2(n4025), 
        .ZN(n19826) );
  MOAI22 U28732 ( .A1(n28767), .A2(n4024), .B1(ram[15586]), .B2(n4025), 
        .ZN(n19827) );
  MOAI22 U28733 ( .A1(n28532), .A2(n4024), .B1(ram[15587]), .B2(n4025), 
        .ZN(n19828) );
  MOAI22 U28734 ( .A1(n28297), .A2(n4024), .B1(ram[15588]), .B2(n4025), 
        .ZN(n19829) );
  MOAI22 U28735 ( .A1(n28062), .A2(n4024), .B1(ram[15589]), .B2(n4025), 
        .ZN(n19830) );
  MOAI22 U28736 ( .A1(n27827), .A2(n4024), .B1(ram[15590]), .B2(n4025), 
        .ZN(n19831) );
  MOAI22 U28737 ( .A1(n27592), .A2(n4024), .B1(ram[15591]), .B2(n4025), 
        .ZN(n19832) );
  MOAI22 U28738 ( .A1(n29237), .A2(n4026), .B1(ram[15592]), .B2(n4027), 
        .ZN(n19833) );
  MOAI22 U28739 ( .A1(n29002), .A2(n4026), .B1(ram[15593]), .B2(n4027), 
        .ZN(n19834) );
  MOAI22 U28740 ( .A1(n28767), .A2(n4026), .B1(ram[15594]), .B2(n4027), 
        .ZN(n19835) );
  MOAI22 U28741 ( .A1(n28532), .A2(n4026), .B1(ram[15595]), .B2(n4027), 
        .ZN(n19836) );
  MOAI22 U28742 ( .A1(n28297), .A2(n4026), .B1(ram[15596]), .B2(n4027), 
        .ZN(n19837) );
  MOAI22 U28743 ( .A1(n28062), .A2(n4026), .B1(ram[15597]), .B2(n4027), 
        .ZN(n19838) );
  MOAI22 U28744 ( .A1(n27827), .A2(n4026), .B1(ram[15598]), .B2(n4027), 
        .ZN(n19839) );
  MOAI22 U28745 ( .A1(n27592), .A2(n4026), .B1(ram[15599]), .B2(n4027), 
        .ZN(n19840) );
  MOAI22 U28746 ( .A1(n29238), .A2(n4028), .B1(ram[15600]), .B2(n4029), 
        .ZN(n19841) );
  MOAI22 U28747 ( .A1(n29003), .A2(n4028), .B1(ram[15601]), .B2(n4029), 
        .ZN(n19842) );
  MOAI22 U28748 ( .A1(n28768), .A2(n4028), .B1(ram[15602]), .B2(n4029), 
        .ZN(n19843) );
  MOAI22 U28749 ( .A1(n28533), .A2(n4028), .B1(ram[15603]), .B2(n4029), 
        .ZN(n19844) );
  MOAI22 U28750 ( .A1(n28298), .A2(n4028), .B1(ram[15604]), .B2(n4029), 
        .ZN(n19845) );
  MOAI22 U28751 ( .A1(n28063), .A2(n4028), .B1(ram[15605]), .B2(n4029), 
        .ZN(n19846) );
  MOAI22 U28752 ( .A1(n27828), .A2(n4028), .B1(ram[15606]), .B2(n4029), 
        .ZN(n19847) );
  MOAI22 U28753 ( .A1(n27593), .A2(n4028), .B1(ram[15607]), .B2(n4029), 
        .ZN(n19848) );
  MOAI22 U28754 ( .A1(n29238), .A2(n4030), .B1(ram[15608]), .B2(n4031), 
        .ZN(n19849) );
  MOAI22 U28755 ( .A1(n29003), .A2(n4030), .B1(ram[15609]), .B2(n4031), 
        .ZN(n19850) );
  MOAI22 U28756 ( .A1(n28768), .A2(n4030), .B1(ram[15610]), .B2(n4031), 
        .ZN(n19851) );
  MOAI22 U28757 ( .A1(n28533), .A2(n4030), .B1(ram[15611]), .B2(n4031), 
        .ZN(n19852) );
  MOAI22 U28758 ( .A1(n28298), .A2(n4030), .B1(ram[15612]), .B2(n4031), 
        .ZN(n19853) );
  MOAI22 U28759 ( .A1(n28063), .A2(n4030), .B1(ram[15613]), .B2(n4031), 
        .ZN(n19854) );
  MOAI22 U28760 ( .A1(n27828), .A2(n4030), .B1(ram[15614]), .B2(n4031), 
        .ZN(n19855) );
  MOAI22 U28761 ( .A1(n27593), .A2(n4030), .B1(ram[15615]), .B2(n4031), 
        .ZN(n19856) );
  MOAI22 U28762 ( .A1(n29238), .A2(n4032), .B1(ram[15616]), .B2(n4033), 
        .ZN(n19857) );
  MOAI22 U28763 ( .A1(n29003), .A2(n4032), .B1(ram[15617]), .B2(n4033), 
        .ZN(n19858) );
  MOAI22 U28764 ( .A1(n28768), .A2(n4032), .B1(ram[15618]), .B2(n4033), 
        .ZN(n19859) );
  MOAI22 U28765 ( .A1(n28533), .A2(n4032), .B1(ram[15619]), .B2(n4033), 
        .ZN(n19860) );
  MOAI22 U28766 ( .A1(n28298), .A2(n4032), .B1(ram[15620]), .B2(n4033), 
        .ZN(n19861) );
  MOAI22 U28767 ( .A1(n28063), .A2(n4032), .B1(ram[15621]), .B2(n4033), 
        .ZN(n19862) );
  MOAI22 U28768 ( .A1(n27828), .A2(n4032), .B1(ram[15622]), .B2(n4033), 
        .ZN(n19863) );
  MOAI22 U28769 ( .A1(n27593), .A2(n4032), .B1(ram[15623]), .B2(n4033), 
        .ZN(n19864) );
  MOAI22 U28770 ( .A1(n29238), .A2(n4034), .B1(ram[15624]), .B2(n4035), 
        .ZN(n19865) );
  MOAI22 U28771 ( .A1(n29003), .A2(n4034), .B1(ram[15625]), .B2(n4035), 
        .ZN(n19866) );
  MOAI22 U28772 ( .A1(n28768), .A2(n4034), .B1(ram[15626]), .B2(n4035), 
        .ZN(n19867) );
  MOAI22 U28773 ( .A1(n28533), .A2(n4034), .B1(ram[15627]), .B2(n4035), 
        .ZN(n19868) );
  MOAI22 U28774 ( .A1(n28298), .A2(n4034), .B1(ram[15628]), .B2(n4035), 
        .ZN(n19869) );
  MOAI22 U28775 ( .A1(n28063), .A2(n4034), .B1(ram[15629]), .B2(n4035), 
        .ZN(n19870) );
  MOAI22 U28776 ( .A1(n27828), .A2(n4034), .B1(ram[15630]), .B2(n4035), 
        .ZN(n19871) );
  MOAI22 U28777 ( .A1(n27593), .A2(n4034), .B1(ram[15631]), .B2(n4035), 
        .ZN(n19872) );
  MOAI22 U28778 ( .A1(n29238), .A2(n4036), .B1(ram[15632]), .B2(n4037), 
        .ZN(n19873) );
  MOAI22 U28779 ( .A1(n29003), .A2(n4036), .B1(ram[15633]), .B2(n4037), 
        .ZN(n19874) );
  MOAI22 U28780 ( .A1(n28768), .A2(n4036), .B1(ram[15634]), .B2(n4037), 
        .ZN(n19875) );
  MOAI22 U28781 ( .A1(n28533), .A2(n4036), .B1(ram[15635]), .B2(n4037), 
        .ZN(n19876) );
  MOAI22 U28782 ( .A1(n28298), .A2(n4036), .B1(ram[15636]), .B2(n4037), 
        .ZN(n19877) );
  MOAI22 U28783 ( .A1(n28063), .A2(n4036), .B1(ram[15637]), .B2(n4037), 
        .ZN(n19878) );
  MOAI22 U28784 ( .A1(n27828), .A2(n4036), .B1(ram[15638]), .B2(n4037), 
        .ZN(n19879) );
  MOAI22 U28785 ( .A1(n27593), .A2(n4036), .B1(ram[15639]), .B2(n4037), 
        .ZN(n19880) );
  MOAI22 U28786 ( .A1(n29238), .A2(n4038), .B1(ram[15640]), .B2(n4039), 
        .ZN(n19881) );
  MOAI22 U28787 ( .A1(n29003), .A2(n4038), .B1(ram[15641]), .B2(n4039), 
        .ZN(n19882) );
  MOAI22 U28788 ( .A1(n28768), .A2(n4038), .B1(ram[15642]), .B2(n4039), 
        .ZN(n19883) );
  MOAI22 U28789 ( .A1(n28533), .A2(n4038), .B1(ram[15643]), .B2(n4039), 
        .ZN(n19884) );
  MOAI22 U28790 ( .A1(n28298), .A2(n4038), .B1(ram[15644]), .B2(n4039), 
        .ZN(n19885) );
  MOAI22 U28791 ( .A1(n28063), .A2(n4038), .B1(ram[15645]), .B2(n4039), 
        .ZN(n19886) );
  MOAI22 U28792 ( .A1(n27828), .A2(n4038), .B1(ram[15646]), .B2(n4039), 
        .ZN(n19887) );
  MOAI22 U28793 ( .A1(n27593), .A2(n4038), .B1(ram[15647]), .B2(n4039), 
        .ZN(n19888) );
  MOAI22 U28794 ( .A1(n29238), .A2(n4040), .B1(ram[15648]), .B2(n4041), 
        .ZN(n19889) );
  MOAI22 U28795 ( .A1(n29003), .A2(n4040), .B1(ram[15649]), .B2(n4041), 
        .ZN(n19890) );
  MOAI22 U28796 ( .A1(n28768), .A2(n4040), .B1(ram[15650]), .B2(n4041), 
        .ZN(n19891) );
  MOAI22 U28797 ( .A1(n28533), .A2(n4040), .B1(ram[15651]), .B2(n4041), 
        .ZN(n19892) );
  MOAI22 U28798 ( .A1(n28298), .A2(n4040), .B1(ram[15652]), .B2(n4041), 
        .ZN(n19893) );
  MOAI22 U28799 ( .A1(n28063), .A2(n4040), .B1(ram[15653]), .B2(n4041), 
        .ZN(n19894) );
  MOAI22 U28800 ( .A1(n27828), .A2(n4040), .B1(ram[15654]), .B2(n4041), 
        .ZN(n19895) );
  MOAI22 U28801 ( .A1(n27593), .A2(n4040), .B1(ram[15655]), .B2(n4041), 
        .ZN(n19896) );
  MOAI22 U28802 ( .A1(n29238), .A2(n4042), .B1(ram[15656]), .B2(n4043), 
        .ZN(n19897) );
  MOAI22 U28803 ( .A1(n29003), .A2(n4042), .B1(ram[15657]), .B2(n4043), 
        .ZN(n19898) );
  MOAI22 U28804 ( .A1(n28768), .A2(n4042), .B1(ram[15658]), .B2(n4043), 
        .ZN(n19899) );
  MOAI22 U28805 ( .A1(n28533), .A2(n4042), .B1(ram[15659]), .B2(n4043), 
        .ZN(n19900) );
  MOAI22 U28806 ( .A1(n28298), .A2(n4042), .B1(ram[15660]), .B2(n4043), 
        .ZN(n19901) );
  MOAI22 U28807 ( .A1(n28063), .A2(n4042), .B1(ram[15661]), .B2(n4043), 
        .ZN(n19902) );
  MOAI22 U28808 ( .A1(n27828), .A2(n4042), .B1(ram[15662]), .B2(n4043), 
        .ZN(n19903) );
  MOAI22 U28809 ( .A1(n27593), .A2(n4042), .B1(ram[15663]), .B2(n4043), 
        .ZN(n19904) );
  MOAI22 U28810 ( .A1(n29238), .A2(n4044), .B1(ram[15664]), .B2(n4045), 
        .ZN(n19905) );
  MOAI22 U28811 ( .A1(n29003), .A2(n4044), .B1(ram[15665]), .B2(n4045), 
        .ZN(n19906) );
  MOAI22 U28812 ( .A1(n28768), .A2(n4044), .B1(ram[15666]), .B2(n4045), 
        .ZN(n19907) );
  MOAI22 U28813 ( .A1(n28533), .A2(n4044), .B1(ram[15667]), .B2(n4045), 
        .ZN(n19908) );
  MOAI22 U28814 ( .A1(n28298), .A2(n4044), .B1(ram[15668]), .B2(n4045), 
        .ZN(n19909) );
  MOAI22 U28815 ( .A1(n28063), .A2(n4044), .B1(ram[15669]), .B2(n4045), 
        .ZN(n19910) );
  MOAI22 U28816 ( .A1(n27828), .A2(n4044), .B1(ram[15670]), .B2(n4045), 
        .ZN(n19911) );
  MOAI22 U28817 ( .A1(n27593), .A2(n4044), .B1(ram[15671]), .B2(n4045), 
        .ZN(n19912) );
  MOAI22 U28818 ( .A1(n29238), .A2(n4046), .B1(ram[15672]), .B2(n4047), 
        .ZN(n19913) );
  MOAI22 U28819 ( .A1(n29003), .A2(n4046), .B1(ram[15673]), .B2(n4047), 
        .ZN(n19914) );
  MOAI22 U28820 ( .A1(n28768), .A2(n4046), .B1(ram[15674]), .B2(n4047), 
        .ZN(n19915) );
  MOAI22 U28821 ( .A1(n28533), .A2(n4046), .B1(ram[15675]), .B2(n4047), 
        .ZN(n19916) );
  MOAI22 U28822 ( .A1(n28298), .A2(n4046), .B1(ram[15676]), .B2(n4047), 
        .ZN(n19917) );
  MOAI22 U28823 ( .A1(n28063), .A2(n4046), .B1(ram[15677]), .B2(n4047), 
        .ZN(n19918) );
  MOAI22 U28824 ( .A1(n27828), .A2(n4046), .B1(ram[15678]), .B2(n4047), 
        .ZN(n19919) );
  MOAI22 U28825 ( .A1(n27593), .A2(n4046), .B1(ram[15679]), .B2(n4047), 
        .ZN(n19920) );
  MOAI22 U28826 ( .A1(n29238), .A2(n4048), .B1(ram[15680]), .B2(n4049), 
        .ZN(n19921) );
  MOAI22 U28827 ( .A1(n29003), .A2(n4048), .B1(ram[15681]), .B2(n4049), 
        .ZN(n19922) );
  MOAI22 U28828 ( .A1(n28768), .A2(n4048), .B1(ram[15682]), .B2(n4049), 
        .ZN(n19923) );
  MOAI22 U28829 ( .A1(n28533), .A2(n4048), .B1(ram[15683]), .B2(n4049), 
        .ZN(n19924) );
  MOAI22 U28830 ( .A1(n28298), .A2(n4048), .B1(ram[15684]), .B2(n4049), 
        .ZN(n19925) );
  MOAI22 U28831 ( .A1(n28063), .A2(n4048), .B1(ram[15685]), .B2(n4049), 
        .ZN(n19926) );
  MOAI22 U28832 ( .A1(n27828), .A2(n4048), .B1(ram[15686]), .B2(n4049), 
        .ZN(n19927) );
  MOAI22 U28833 ( .A1(n27593), .A2(n4048), .B1(ram[15687]), .B2(n4049), 
        .ZN(n19928) );
  MOAI22 U28834 ( .A1(n29238), .A2(n4050), .B1(ram[15688]), .B2(n4051), 
        .ZN(n19929) );
  MOAI22 U28835 ( .A1(n29003), .A2(n4050), .B1(ram[15689]), .B2(n4051), 
        .ZN(n19930) );
  MOAI22 U28836 ( .A1(n28768), .A2(n4050), .B1(ram[15690]), .B2(n4051), 
        .ZN(n19931) );
  MOAI22 U28837 ( .A1(n28533), .A2(n4050), .B1(ram[15691]), .B2(n4051), 
        .ZN(n19932) );
  MOAI22 U28838 ( .A1(n28298), .A2(n4050), .B1(ram[15692]), .B2(n4051), 
        .ZN(n19933) );
  MOAI22 U28839 ( .A1(n28063), .A2(n4050), .B1(ram[15693]), .B2(n4051), 
        .ZN(n19934) );
  MOAI22 U28840 ( .A1(n27828), .A2(n4050), .B1(ram[15694]), .B2(n4051), 
        .ZN(n19935) );
  MOAI22 U28841 ( .A1(n27593), .A2(n4050), .B1(ram[15695]), .B2(n4051), 
        .ZN(n19936) );
  MOAI22 U28842 ( .A1(n29238), .A2(n4052), .B1(ram[15696]), .B2(n4053), 
        .ZN(n19937) );
  MOAI22 U28843 ( .A1(n29003), .A2(n4052), .B1(ram[15697]), .B2(n4053), 
        .ZN(n19938) );
  MOAI22 U28844 ( .A1(n28768), .A2(n4052), .B1(ram[15698]), .B2(n4053), 
        .ZN(n19939) );
  MOAI22 U28845 ( .A1(n28533), .A2(n4052), .B1(ram[15699]), .B2(n4053), 
        .ZN(n19940) );
  MOAI22 U28846 ( .A1(n28298), .A2(n4052), .B1(ram[15700]), .B2(n4053), 
        .ZN(n19941) );
  MOAI22 U28847 ( .A1(n28063), .A2(n4052), .B1(ram[15701]), .B2(n4053), 
        .ZN(n19942) );
  MOAI22 U28848 ( .A1(n27828), .A2(n4052), .B1(ram[15702]), .B2(n4053), 
        .ZN(n19943) );
  MOAI22 U28849 ( .A1(n27593), .A2(n4052), .B1(ram[15703]), .B2(n4053), 
        .ZN(n19944) );
  MOAI22 U28850 ( .A1(n29239), .A2(n4054), .B1(ram[15704]), .B2(n4055), 
        .ZN(n19945) );
  MOAI22 U28851 ( .A1(n29004), .A2(n4054), .B1(ram[15705]), .B2(n4055), 
        .ZN(n19946) );
  MOAI22 U28852 ( .A1(n28769), .A2(n4054), .B1(ram[15706]), .B2(n4055), 
        .ZN(n19947) );
  MOAI22 U28853 ( .A1(n28534), .A2(n4054), .B1(ram[15707]), .B2(n4055), 
        .ZN(n19948) );
  MOAI22 U28854 ( .A1(n28299), .A2(n4054), .B1(ram[15708]), .B2(n4055), 
        .ZN(n19949) );
  MOAI22 U28855 ( .A1(n28064), .A2(n4054), .B1(ram[15709]), .B2(n4055), 
        .ZN(n19950) );
  MOAI22 U28856 ( .A1(n27829), .A2(n4054), .B1(ram[15710]), .B2(n4055), 
        .ZN(n19951) );
  MOAI22 U28857 ( .A1(n27594), .A2(n4054), .B1(ram[15711]), .B2(n4055), 
        .ZN(n19952) );
  MOAI22 U28858 ( .A1(n29239), .A2(n4056), .B1(ram[15712]), .B2(n4057), 
        .ZN(n19953) );
  MOAI22 U28859 ( .A1(n29004), .A2(n4056), .B1(ram[15713]), .B2(n4057), 
        .ZN(n19954) );
  MOAI22 U28860 ( .A1(n28769), .A2(n4056), .B1(ram[15714]), .B2(n4057), 
        .ZN(n19955) );
  MOAI22 U28861 ( .A1(n28534), .A2(n4056), .B1(ram[15715]), .B2(n4057), 
        .ZN(n19956) );
  MOAI22 U28862 ( .A1(n28299), .A2(n4056), .B1(ram[15716]), .B2(n4057), 
        .ZN(n19957) );
  MOAI22 U28863 ( .A1(n28064), .A2(n4056), .B1(ram[15717]), .B2(n4057), 
        .ZN(n19958) );
  MOAI22 U28864 ( .A1(n27829), .A2(n4056), .B1(ram[15718]), .B2(n4057), 
        .ZN(n19959) );
  MOAI22 U28865 ( .A1(n27594), .A2(n4056), .B1(ram[15719]), .B2(n4057), 
        .ZN(n19960) );
  MOAI22 U28866 ( .A1(n29239), .A2(n4058), .B1(ram[15720]), .B2(n4059), 
        .ZN(n19961) );
  MOAI22 U28867 ( .A1(n29004), .A2(n4058), .B1(ram[15721]), .B2(n4059), 
        .ZN(n19962) );
  MOAI22 U28868 ( .A1(n28769), .A2(n4058), .B1(ram[15722]), .B2(n4059), 
        .ZN(n19963) );
  MOAI22 U28869 ( .A1(n28534), .A2(n4058), .B1(ram[15723]), .B2(n4059), 
        .ZN(n19964) );
  MOAI22 U28870 ( .A1(n28299), .A2(n4058), .B1(ram[15724]), .B2(n4059), 
        .ZN(n19965) );
  MOAI22 U28871 ( .A1(n28064), .A2(n4058), .B1(ram[15725]), .B2(n4059), 
        .ZN(n19966) );
  MOAI22 U28872 ( .A1(n27829), .A2(n4058), .B1(ram[15726]), .B2(n4059), 
        .ZN(n19967) );
  MOAI22 U28873 ( .A1(n27594), .A2(n4058), .B1(ram[15727]), .B2(n4059), 
        .ZN(n19968) );
  MOAI22 U28874 ( .A1(n29239), .A2(n4060), .B1(ram[15728]), .B2(n4061), 
        .ZN(n19969) );
  MOAI22 U28875 ( .A1(n29004), .A2(n4060), .B1(ram[15729]), .B2(n4061), 
        .ZN(n19970) );
  MOAI22 U28876 ( .A1(n28769), .A2(n4060), .B1(ram[15730]), .B2(n4061), 
        .ZN(n19971) );
  MOAI22 U28877 ( .A1(n28534), .A2(n4060), .B1(ram[15731]), .B2(n4061), 
        .ZN(n19972) );
  MOAI22 U28878 ( .A1(n28299), .A2(n4060), .B1(ram[15732]), .B2(n4061), 
        .ZN(n19973) );
  MOAI22 U28879 ( .A1(n28064), .A2(n4060), .B1(ram[15733]), .B2(n4061), 
        .ZN(n19974) );
  MOAI22 U28880 ( .A1(n27829), .A2(n4060), .B1(ram[15734]), .B2(n4061), 
        .ZN(n19975) );
  MOAI22 U28881 ( .A1(n27594), .A2(n4060), .B1(ram[15735]), .B2(n4061), 
        .ZN(n19976) );
  MOAI22 U28882 ( .A1(n29239), .A2(n4062), .B1(ram[15736]), .B2(n4063), 
        .ZN(n19977) );
  MOAI22 U28883 ( .A1(n29004), .A2(n4062), .B1(ram[15737]), .B2(n4063), 
        .ZN(n19978) );
  MOAI22 U28884 ( .A1(n28769), .A2(n4062), .B1(ram[15738]), .B2(n4063), 
        .ZN(n19979) );
  MOAI22 U28885 ( .A1(n28534), .A2(n4062), .B1(ram[15739]), .B2(n4063), 
        .ZN(n19980) );
  MOAI22 U28886 ( .A1(n28299), .A2(n4062), .B1(ram[15740]), .B2(n4063), 
        .ZN(n19981) );
  MOAI22 U28887 ( .A1(n28064), .A2(n4062), .B1(ram[15741]), .B2(n4063), 
        .ZN(n19982) );
  MOAI22 U28888 ( .A1(n27829), .A2(n4062), .B1(ram[15742]), .B2(n4063), 
        .ZN(n19983) );
  MOAI22 U28889 ( .A1(n27594), .A2(n4062), .B1(ram[15743]), .B2(n4063), 
        .ZN(n19984) );
  MOAI22 U28890 ( .A1(n29239), .A2(n4064), .B1(ram[15744]), .B2(n4065), 
        .ZN(n19985) );
  MOAI22 U28891 ( .A1(n29004), .A2(n4064), .B1(ram[15745]), .B2(n4065), 
        .ZN(n19986) );
  MOAI22 U28892 ( .A1(n28769), .A2(n4064), .B1(ram[15746]), .B2(n4065), 
        .ZN(n19987) );
  MOAI22 U28893 ( .A1(n28534), .A2(n4064), .B1(ram[15747]), .B2(n4065), 
        .ZN(n19988) );
  MOAI22 U28894 ( .A1(n28299), .A2(n4064), .B1(ram[15748]), .B2(n4065), 
        .ZN(n19989) );
  MOAI22 U28895 ( .A1(n28064), .A2(n4064), .B1(ram[15749]), .B2(n4065), 
        .ZN(n19990) );
  MOAI22 U28896 ( .A1(n27829), .A2(n4064), .B1(ram[15750]), .B2(n4065), 
        .ZN(n19991) );
  MOAI22 U28897 ( .A1(n27594), .A2(n4064), .B1(ram[15751]), .B2(n4065), 
        .ZN(n19992) );
  MOAI22 U28898 ( .A1(n29239), .A2(n4066), .B1(ram[15752]), .B2(n4067), 
        .ZN(n19993) );
  MOAI22 U28899 ( .A1(n29004), .A2(n4066), .B1(ram[15753]), .B2(n4067), 
        .ZN(n19994) );
  MOAI22 U28900 ( .A1(n28769), .A2(n4066), .B1(ram[15754]), .B2(n4067), 
        .ZN(n19995) );
  MOAI22 U28901 ( .A1(n28534), .A2(n4066), .B1(ram[15755]), .B2(n4067), 
        .ZN(n19996) );
  MOAI22 U28902 ( .A1(n28299), .A2(n4066), .B1(ram[15756]), .B2(n4067), 
        .ZN(n19997) );
  MOAI22 U28903 ( .A1(n28064), .A2(n4066), .B1(ram[15757]), .B2(n4067), 
        .ZN(n19998) );
  MOAI22 U28904 ( .A1(n27829), .A2(n4066), .B1(ram[15758]), .B2(n4067), 
        .ZN(n19999) );
  MOAI22 U28905 ( .A1(n27594), .A2(n4066), .B1(ram[15759]), .B2(n4067), 
        .ZN(n20000) );
  MOAI22 U28906 ( .A1(n29239), .A2(n4068), .B1(ram[15760]), .B2(n4069), 
        .ZN(n20001) );
  MOAI22 U28907 ( .A1(n29004), .A2(n4068), .B1(ram[15761]), .B2(n4069), 
        .ZN(n20002) );
  MOAI22 U28908 ( .A1(n28769), .A2(n4068), .B1(ram[15762]), .B2(n4069), 
        .ZN(n20003) );
  MOAI22 U28909 ( .A1(n28534), .A2(n4068), .B1(ram[15763]), .B2(n4069), 
        .ZN(n20004) );
  MOAI22 U28910 ( .A1(n28299), .A2(n4068), .B1(ram[15764]), .B2(n4069), 
        .ZN(n20005) );
  MOAI22 U28911 ( .A1(n28064), .A2(n4068), .B1(ram[15765]), .B2(n4069), 
        .ZN(n20006) );
  MOAI22 U28912 ( .A1(n27829), .A2(n4068), .B1(ram[15766]), .B2(n4069), 
        .ZN(n20007) );
  MOAI22 U28913 ( .A1(n27594), .A2(n4068), .B1(ram[15767]), .B2(n4069), 
        .ZN(n20008) );
  MOAI22 U28914 ( .A1(n29239), .A2(n4070), .B1(ram[15768]), .B2(n4071), 
        .ZN(n20009) );
  MOAI22 U28915 ( .A1(n29004), .A2(n4070), .B1(ram[15769]), .B2(n4071), 
        .ZN(n20010) );
  MOAI22 U28916 ( .A1(n28769), .A2(n4070), .B1(ram[15770]), .B2(n4071), 
        .ZN(n20011) );
  MOAI22 U28917 ( .A1(n28534), .A2(n4070), .B1(ram[15771]), .B2(n4071), 
        .ZN(n20012) );
  MOAI22 U28918 ( .A1(n28299), .A2(n4070), .B1(ram[15772]), .B2(n4071), 
        .ZN(n20013) );
  MOAI22 U28919 ( .A1(n28064), .A2(n4070), .B1(ram[15773]), .B2(n4071), 
        .ZN(n20014) );
  MOAI22 U28920 ( .A1(n27829), .A2(n4070), .B1(ram[15774]), .B2(n4071), 
        .ZN(n20015) );
  MOAI22 U28921 ( .A1(n27594), .A2(n4070), .B1(ram[15775]), .B2(n4071), 
        .ZN(n20016) );
  MOAI22 U28922 ( .A1(n29239), .A2(n4072), .B1(ram[15776]), .B2(n4073), 
        .ZN(n20017) );
  MOAI22 U28923 ( .A1(n29004), .A2(n4072), .B1(ram[15777]), .B2(n4073), 
        .ZN(n20018) );
  MOAI22 U28924 ( .A1(n28769), .A2(n4072), .B1(ram[15778]), .B2(n4073), 
        .ZN(n20019) );
  MOAI22 U28925 ( .A1(n28534), .A2(n4072), .B1(ram[15779]), .B2(n4073), 
        .ZN(n20020) );
  MOAI22 U28926 ( .A1(n28299), .A2(n4072), .B1(ram[15780]), .B2(n4073), 
        .ZN(n20021) );
  MOAI22 U28927 ( .A1(n28064), .A2(n4072), .B1(ram[15781]), .B2(n4073), 
        .ZN(n20022) );
  MOAI22 U28928 ( .A1(n27829), .A2(n4072), .B1(ram[15782]), .B2(n4073), 
        .ZN(n20023) );
  MOAI22 U28929 ( .A1(n27594), .A2(n4072), .B1(ram[15783]), .B2(n4073), 
        .ZN(n20024) );
  MOAI22 U28930 ( .A1(n29239), .A2(n4074), .B1(ram[15784]), .B2(n4075), 
        .ZN(n20025) );
  MOAI22 U28931 ( .A1(n29004), .A2(n4074), .B1(ram[15785]), .B2(n4075), 
        .ZN(n20026) );
  MOAI22 U28932 ( .A1(n28769), .A2(n4074), .B1(ram[15786]), .B2(n4075), 
        .ZN(n20027) );
  MOAI22 U28933 ( .A1(n28534), .A2(n4074), .B1(ram[15787]), .B2(n4075), 
        .ZN(n20028) );
  MOAI22 U28934 ( .A1(n28299), .A2(n4074), .B1(ram[15788]), .B2(n4075), 
        .ZN(n20029) );
  MOAI22 U28935 ( .A1(n28064), .A2(n4074), .B1(ram[15789]), .B2(n4075), 
        .ZN(n20030) );
  MOAI22 U28936 ( .A1(n27829), .A2(n4074), .B1(ram[15790]), .B2(n4075), 
        .ZN(n20031) );
  MOAI22 U28937 ( .A1(n27594), .A2(n4074), .B1(ram[15791]), .B2(n4075), 
        .ZN(n20032) );
  MOAI22 U28938 ( .A1(n29239), .A2(n4076), .B1(ram[15792]), .B2(n4077), 
        .ZN(n20033) );
  MOAI22 U28939 ( .A1(n29004), .A2(n4076), .B1(ram[15793]), .B2(n4077), 
        .ZN(n20034) );
  MOAI22 U28940 ( .A1(n28769), .A2(n4076), .B1(ram[15794]), .B2(n4077), 
        .ZN(n20035) );
  MOAI22 U28941 ( .A1(n28534), .A2(n4076), .B1(ram[15795]), .B2(n4077), 
        .ZN(n20036) );
  MOAI22 U28942 ( .A1(n28299), .A2(n4076), .B1(ram[15796]), .B2(n4077), 
        .ZN(n20037) );
  MOAI22 U28943 ( .A1(n28064), .A2(n4076), .B1(ram[15797]), .B2(n4077), 
        .ZN(n20038) );
  MOAI22 U28944 ( .A1(n27829), .A2(n4076), .B1(ram[15798]), .B2(n4077), 
        .ZN(n20039) );
  MOAI22 U28945 ( .A1(n27594), .A2(n4076), .B1(ram[15799]), .B2(n4077), 
        .ZN(n20040) );
  MOAI22 U28946 ( .A1(n29239), .A2(n4078), .B1(ram[15800]), .B2(n4079), 
        .ZN(n20041) );
  MOAI22 U28947 ( .A1(n29004), .A2(n4078), .B1(ram[15801]), .B2(n4079), 
        .ZN(n20042) );
  MOAI22 U28948 ( .A1(n28769), .A2(n4078), .B1(ram[15802]), .B2(n4079), 
        .ZN(n20043) );
  MOAI22 U28949 ( .A1(n28534), .A2(n4078), .B1(ram[15803]), .B2(n4079), 
        .ZN(n20044) );
  MOAI22 U28950 ( .A1(n28299), .A2(n4078), .B1(ram[15804]), .B2(n4079), 
        .ZN(n20045) );
  MOAI22 U28951 ( .A1(n28064), .A2(n4078), .B1(ram[15805]), .B2(n4079), 
        .ZN(n20046) );
  MOAI22 U28952 ( .A1(n27829), .A2(n4078), .B1(ram[15806]), .B2(n4079), 
        .ZN(n20047) );
  MOAI22 U28953 ( .A1(n27594), .A2(n4078), .B1(ram[15807]), .B2(n4079), 
        .ZN(n20048) );
  MOAI22 U28954 ( .A1(n29240), .A2(n4080), .B1(ram[15808]), .B2(n4081), 
        .ZN(n20049) );
  MOAI22 U28955 ( .A1(n29005), .A2(n4080), .B1(ram[15809]), .B2(n4081), 
        .ZN(n20050) );
  MOAI22 U28956 ( .A1(n28770), .A2(n4080), .B1(ram[15810]), .B2(n4081), 
        .ZN(n20051) );
  MOAI22 U28957 ( .A1(n28535), .A2(n4080), .B1(ram[15811]), .B2(n4081), 
        .ZN(n20052) );
  MOAI22 U28958 ( .A1(n28300), .A2(n4080), .B1(ram[15812]), .B2(n4081), 
        .ZN(n20053) );
  MOAI22 U28959 ( .A1(n28065), .A2(n4080), .B1(ram[15813]), .B2(n4081), 
        .ZN(n20054) );
  MOAI22 U28960 ( .A1(n27830), .A2(n4080), .B1(ram[15814]), .B2(n4081), 
        .ZN(n20055) );
  MOAI22 U28961 ( .A1(n27595), .A2(n4080), .B1(ram[15815]), .B2(n4081), 
        .ZN(n20056) );
  MOAI22 U28962 ( .A1(n29240), .A2(n4082), .B1(ram[15816]), .B2(n4083), 
        .ZN(n20057) );
  MOAI22 U28963 ( .A1(n29005), .A2(n4082), .B1(ram[15817]), .B2(n4083), 
        .ZN(n20058) );
  MOAI22 U28964 ( .A1(n28770), .A2(n4082), .B1(ram[15818]), .B2(n4083), 
        .ZN(n20059) );
  MOAI22 U28965 ( .A1(n28535), .A2(n4082), .B1(ram[15819]), .B2(n4083), 
        .ZN(n20060) );
  MOAI22 U28966 ( .A1(n28300), .A2(n4082), .B1(ram[15820]), .B2(n4083), 
        .ZN(n20061) );
  MOAI22 U28967 ( .A1(n28065), .A2(n4082), .B1(ram[15821]), .B2(n4083), 
        .ZN(n20062) );
  MOAI22 U28968 ( .A1(n27830), .A2(n4082), .B1(ram[15822]), .B2(n4083), 
        .ZN(n20063) );
  MOAI22 U28969 ( .A1(n27595), .A2(n4082), .B1(ram[15823]), .B2(n4083), 
        .ZN(n20064) );
  MOAI22 U28970 ( .A1(n29240), .A2(n4084), .B1(ram[15824]), .B2(n4085), 
        .ZN(n20065) );
  MOAI22 U28971 ( .A1(n29005), .A2(n4084), .B1(ram[15825]), .B2(n4085), 
        .ZN(n20066) );
  MOAI22 U28972 ( .A1(n28770), .A2(n4084), .B1(ram[15826]), .B2(n4085), 
        .ZN(n20067) );
  MOAI22 U28973 ( .A1(n28535), .A2(n4084), .B1(ram[15827]), .B2(n4085), 
        .ZN(n20068) );
  MOAI22 U28974 ( .A1(n28300), .A2(n4084), .B1(ram[15828]), .B2(n4085), 
        .ZN(n20069) );
  MOAI22 U28975 ( .A1(n28065), .A2(n4084), .B1(ram[15829]), .B2(n4085), 
        .ZN(n20070) );
  MOAI22 U28976 ( .A1(n27830), .A2(n4084), .B1(ram[15830]), .B2(n4085), 
        .ZN(n20071) );
  MOAI22 U28977 ( .A1(n27595), .A2(n4084), .B1(ram[15831]), .B2(n4085), 
        .ZN(n20072) );
  MOAI22 U28978 ( .A1(n29240), .A2(n4086), .B1(ram[15832]), .B2(n4087), 
        .ZN(n20073) );
  MOAI22 U28979 ( .A1(n29005), .A2(n4086), .B1(ram[15833]), .B2(n4087), 
        .ZN(n20074) );
  MOAI22 U28980 ( .A1(n28770), .A2(n4086), .B1(ram[15834]), .B2(n4087), 
        .ZN(n20075) );
  MOAI22 U28981 ( .A1(n28535), .A2(n4086), .B1(ram[15835]), .B2(n4087), 
        .ZN(n20076) );
  MOAI22 U28982 ( .A1(n28300), .A2(n4086), .B1(ram[15836]), .B2(n4087), 
        .ZN(n20077) );
  MOAI22 U28983 ( .A1(n28065), .A2(n4086), .B1(ram[15837]), .B2(n4087), 
        .ZN(n20078) );
  MOAI22 U28984 ( .A1(n27830), .A2(n4086), .B1(ram[15838]), .B2(n4087), 
        .ZN(n20079) );
  MOAI22 U28985 ( .A1(n27595), .A2(n4086), .B1(ram[15839]), .B2(n4087), 
        .ZN(n20080) );
  MOAI22 U28986 ( .A1(n29240), .A2(n4088), .B1(ram[15840]), .B2(n4089), 
        .ZN(n20081) );
  MOAI22 U28987 ( .A1(n29005), .A2(n4088), .B1(ram[15841]), .B2(n4089), 
        .ZN(n20082) );
  MOAI22 U28988 ( .A1(n28770), .A2(n4088), .B1(ram[15842]), .B2(n4089), 
        .ZN(n20083) );
  MOAI22 U28989 ( .A1(n28535), .A2(n4088), .B1(ram[15843]), .B2(n4089), 
        .ZN(n20084) );
  MOAI22 U28990 ( .A1(n28300), .A2(n4088), .B1(ram[15844]), .B2(n4089), 
        .ZN(n20085) );
  MOAI22 U28991 ( .A1(n28065), .A2(n4088), .B1(ram[15845]), .B2(n4089), 
        .ZN(n20086) );
  MOAI22 U28992 ( .A1(n27830), .A2(n4088), .B1(ram[15846]), .B2(n4089), 
        .ZN(n20087) );
  MOAI22 U28993 ( .A1(n27595), .A2(n4088), .B1(ram[15847]), .B2(n4089), 
        .ZN(n20088) );
  MOAI22 U28994 ( .A1(n29240), .A2(n4090), .B1(ram[15848]), .B2(n4091), 
        .ZN(n20089) );
  MOAI22 U28995 ( .A1(n29005), .A2(n4090), .B1(ram[15849]), .B2(n4091), 
        .ZN(n20090) );
  MOAI22 U28996 ( .A1(n28770), .A2(n4090), .B1(ram[15850]), .B2(n4091), 
        .ZN(n20091) );
  MOAI22 U28997 ( .A1(n28535), .A2(n4090), .B1(ram[15851]), .B2(n4091), 
        .ZN(n20092) );
  MOAI22 U28998 ( .A1(n28300), .A2(n4090), .B1(ram[15852]), .B2(n4091), 
        .ZN(n20093) );
  MOAI22 U28999 ( .A1(n28065), .A2(n4090), .B1(ram[15853]), .B2(n4091), 
        .ZN(n20094) );
  MOAI22 U29000 ( .A1(n27830), .A2(n4090), .B1(ram[15854]), .B2(n4091), 
        .ZN(n20095) );
  MOAI22 U29001 ( .A1(n27595), .A2(n4090), .B1(ram[15855]), .B2(n4091), 
        .ZN(n20096) );
  MOAI22 U29002 ( .A1(n29240), .A2(n4092), .B1(ram[15856]), .B2(n4093), 
        .ZN(n20097) );
  MOAI22 U29003 ( .A1(n29005), .A2(n4092), .B1(ram[15857]), .B2(n4093), 
        .ZN(n20098) );
  MOAI22 U29004 ( .A1(n28770), .A2(n4092), .B1(ram[15858]), .B2(n4093), 
        .ZN(n20099) );
  MOAI22 U29005 ( .A1(n28535), .A2(n4092), .B1(ram[15859]), .B2(n4093), 
        .ZN(n20100) );
  MOAI22 U29006 ( .A1(n28300), .A2(n4092), .B1(ram[15860]), .B2(n4093), 
        .ZN(n20101) );
  MOAI22 U29007 ( .A1(n28065), .A2(n4092), .B1(ram[15861]), .B2(n4093), 
        .ZN(n20102) );
  MOAI22 U29008 ( .A1(n27830), .A2(n4092), .B1(ram[15862]), .B2(n4093), 
        .ZN(n20103) );
  MOAI22 U29009 ( .A1(n27595), .A2(n4092), .B1(ram[15863]), .B2(n4093), 
        .ZN(n20104) );
  MOAI22 U29010 ( .A1(n29240), .A2(n4094), .B1(ram[15864]), .B2(n4095), 
        .ZN(n20105) );
  MOAI22 U29011 ( .A1(n29005), .A2(n4094), .B1(ram[15865]), .B2(n4095), 
        .ZN(n20106) );
  MOAI22 U29012 ( .A1(n28770), .A2(n4094), .B1(ram[15866]), .B2(n4095), 
        .ZN(n20107) );
  MOAI22 U29013 ( .A1(n28535), .A2(n4094), .B1(ram[15867]), .B2(n4095), 
        .ZN(n20108) );
  MOAI22 U29014 ( .A1(n28300), .A2(n4094), .B1(ram[15868]), .B2(n4095), 
        .ZN(n20109) );
  MOAI22 U29015 ( .A1(n28065), .A2(n4094), .B1(ram[15869]), .B2(n4095), 
        .ZN(n20110) );
  MOAI22 U29016 ( .A1(n27830), .A2(n4094), .B1(ram[15870]), .B2(n4095), 
        .ZN(n20111) );
  MOAI22 U29017 ( .A1(n27595), .A2(n4094), .B1(ram[15871]), .B2(n4095), 
        .ZN(n20112) );
  MOAI22 U29018 ( .A1(n29240), .A2(n4096), .B1(ram[15872]), .B2(n4097), 
        .ZN(n20113) );
  MOAI22 U29019 ( .A1(n29005), .A2(n4096), .B1(ram[15873]), .B2(n4097), 
        .ZN(n20114) );
  MOAI22 U29020 ( .A1(n28770), .A2(n4096), .B1(ram[15874]), .B2(n4097), 
        .ZN(n20115) );
  MOAI22 U29021 ( .A1(n28535), .A2(n4096), .B1(ram[15875]), .B2(n4097), 
        .ZN(n20116) );
  MOAI22 U29022 ( .A1(n28300), .A2(n4096), .B1(ram[15876]), .B2(n4097), 
        .ZN(n20117) );
  MOAI22 U29023 ( .A1(n28065), .A2(n4096), .B1(ram[15877]), .B2(n4097), 
        .ZN(n20118) );
  MOAI22 U29024 ( .A1(n27830), .A2(n4096), .B1(ram[15878]), .B2(n4097), 
        .ZN(n20119) );
  MOAI22 U29025 ( .A1(n27595), .A2(n4096), .B1(ram[15879]), .B2(n4097), 
        .ZN(n20120) );
  MOAI22 U29026 ( .A1(n29240), .A2(n4101), .B1(ram[15880]), .B2(n4102), 
        .ZN(n20121) );
  MOAI22 U29027 ( .A1(n29005), .A2(n4101), .B1(ram[15881]), .B2(n4102), 
        .ZN(n20122) );
  MOAI22 U29028 ( .A1(n28770), .A2(n4101), .B1(ram[15882]), .B2(n4102), 
        .ZN(n20123) );
  MOAI22 U29029 ( .A1(n28535), .A2(n4101), .B1(ram[15883]), .B2(n4102), 
        .ZN(n20124) );
  MOAI22 U29030 ( .A1(n28300), .A2(n4101), .B1(ram[15884]), .B2(n4102), 
        .ZN(n20125) );
  MOAI22 U29031 ( .A1(n28065), .A2(n4101), .B1(ram[15885]), .B2(n4102), 
        .ZN(n20126) );
  MOAI22 U29032 ( .A1(n27830), .A2(n4101), .B1(ram[15886]), .B2(n4102), 
        .ZN(n20127) );
  MOAI22 U29033 ( .A1(n27595), .A2(n4101), .B1(ram[15887]), .B2(n4102), 
        .ZN(n20128) );
  MOAI22 U29034 ( .A1(n29240), .A2(n4104), .B1(ram[15888]), .B2(n4105), 
        .ZN(n20129) );
  MOAI22 U29035 ( .A1(n29005), .A2(n4104), .B1(ram[15889]), .B2(n4105), 
        .ZN(n20130) );
  MOAI22 U29036 ( .A1(n28770), .A2(n4104), .B1(ram[15890]), .B2(n4105), 
        .ZN(n20131) );
  MOAI22 U29037 ( .A1(n28535), .A2(n4104), .B1(ram[15891]), .B2(n4105), 
        .ZN(n20132) );
  MOAI22 U29038 ( .A1(n28300), .A2(n4104), .B1(ram[15892]), .B2(n4105), 
        .ZN(n20133) );
  MOAI22 U29039 ( .A1(n28065), .A2(n4104), .B1(ram[15893]), .B2(n4105), 
        .ZN(n20134) );
  MOAI22 U29040 ( .A1(n27830), .A2(n4104), .B1(ram[15894]), .B2(n4105), 
        .ZN(n20135) );
  MOAI22 U29041 ( .A1(n27595), .A2(n4104), .B1(ram[15895]), .B2(n4105), 
        .ZN(n20136) );
  MOAI22 U29042 ( .A1(n29240), .A2(n4107), .B1(ram[15896]), .B2(n4108), 
        .ZN(n20137) );
  MOAI22 U29043 ( .A1(n29005), .A2(n4107), .B1(ram[15897]), .B2(n4108), 
        .ZN(n20138) );
  MOAI22 U29044 ( .A1(n28770), .A2(n4107), .B1(ram[15898]), .B2(n4108), 
        .ZN(n20139) );
  MOAI22 U29045 ( .A1(n28535), .A2(n4107), .B1(ram[15899]), .B2(n4108), 
        .ZN(n20140) );
  MOAI22 U29046 ( .A1(n28300), .A2(n4107), .B1(ram[15900]), .B2(n4108), 
        .ZN(n20141) );
  MOAI22 U29047 ( .A1(n28065), .A2(n4107), .B1(ram[15901]), .B2(n4108), 
        .ZN(n20142) );
  MOAI22 U29048 ( .A1(n27830), .A2(n4107), .B1(ram[15902]), .B2(n4108), 
        .ZN(n20143) );
  MOAI22 U29049 ( .A1(n27595), .A2(n4107), .B1(ram[15903]), .B2(n4108), 
        .ZN(n20144) );
  MOAI22 U29050 ( .A1(n29240), .A2(n4110), .B1(ram[15904]), .B2(n4111), 
        .ZN(n20145) );
  MOAI22 U29051 ( .A1(n29005), .A2(n4110), .B1(ram[15905]), .B2(n4111), 
        .ZN(n20146) );
  MOAI22 U29052 ( .A1(n28770), .A2(n4110), .B1(ram[15906]), .B2(n4111), 
        .ZN(n20147) );
  MOAI22 U29053 ( .A1(n28535), .A2(n4110), .B1(ram[15907]), .B2(n4111), 
        .ZN(n20148) );
  MOAI22 U29054 ( .A1(n28300), .A2(n4110), .B1(ram[15908]), .B2(n4111), 
        .ZN(n20149) );
  MOAI22 U29055 ( .A1(n28065), .A2(n4110), .B1(ram[15909]), .B2(n4111), 
        .ZN(n20150) );
  MOAI22 U29056 ( .A1(n27830), .A2(n4110), .B1(ram[15910]), .B2(n4111), 
        .ZN(n20151) );
  MOAI22 U29057 ( .A1(n27595), .A2(n4110), .B1(ram[15911]), .B2(n4111), 
        .ZN(n20152) );
  MOAI22 U29058 ( .A1(n29241), .A2(n4113), .B1(ram[15912]), .B2(n4114), 
        .ZN(n20153) );
  MOAI22 U29059 ( .A1(n29006), .A2(n4113), .B1(ram[15913]), .B2(n4114), 
        .ZN(n20154) );
  MOAI22 U29060 ( .A1(n28771), .A2(n4113), .B1(ram[15914]), .B2(n4114), 
        .ZN(n20155) );
  MOAI22 U29061 ( .A1(n28536), .A2(n4113), .B1(ram[15915]), .B2(n4114), 
        .ZN(n20156) );
  MOAI22 U29062 ( .A1(n28301), .A2(n4113), .B1(ram[15916]), .B2(n4114), 
        .ZN(n20157) );
  MOAI22 U29063 ( .A1(n28066), .A2(n4113), .B1(ram[15917]), .B2(n4114), 
        .ZN(n20158) );
  MOAI22 U29064 ( .A1(n27831), .A2(n4113), .B1(ram[15918]), .B2(n4114), 
        .ZN(n20159) );
  MOAI22 U29065 ( .A1(n27596), .A2(n4113), .B1(ram[15919]), .B2(n4114), 
        .ZN(n20160) );
  MOAI22 U29066 ( .A1(n29241), .A2(n4116), .B1(ram[15920]), .B2(n4117), 
        .ZN(n20161) );
  MOAI22 U29067 ( .A1(n29006), .A2(n4116), .B1(ram[15921]), .B2(n4117), 
        .ZN(n20162) );
  MOAI22 U29068 ( .A1(n28771), .A2(n4116), .B1(ram[15922]), .B2(n4117), 
        .ZN(n20163) );
  MOAI22 U29069 ( .A1(n28536), .A2(n4116), .B1(ram[15923]), .B2(n4117), 
        .ZN(n20164) );
  MOAI22 U29070 ( .A1(n28301), .A2(n4116), .B1(ram[15924]), .B2(n4117), 
        .ZN(n20165) );
  MOAI22 U29071 ( .A1(n28066), .A2(n4116), .B1(ram[15925]), .B2(n4117), 
        .ZN(n20166) );
  MOAI22 U29072 ( .A1(n27831), .A2(n4116), .B1(ram[15926]), .B2(n4117), 
        .ZN(n20167) );
  MOAI22 U29073 ( .A1(n27596), .A2(n4116), .B1(ram[15927]), .B2(n4117), 
        .ZN(n20168) );
  MOAI22 U29074 ( .A1(n29241), .A2(n4119), .B1(ram[15928]), .B2(n4120), 
        .ZN(n20169) );
  MOAI22 U29075 ( .A1(n29006), .A2(n4119), .B1(ram[15929]), .B2(n4120), 
        .ZN(n20170) );
  MOAI22 U29076 ( .A1(n28771), .A2(n4119), .B1(ram[15930]), .B2(n4120), 
        .ZN(n20171) );
  MOAI22 U29077 ( .A1(n28536), .A2(n4119), .B1(ram[15931]), .B2(n4120), 
        .ZN(n20172) );
  MOAI22 U29078 ( .A1(n28301), .A2(n4119), .B1(ram[15932]), .B2(n4120), 
        .ZN(n20173) );
  MOAI22 U29079 ( .A1(n28066), .A2(n4119), .B1(ram[15933]), .B2(n4120), 
        .ZN(n20174) );
  MOAI22 U29080 ( .A1(n27831), .A2(n4119), .B1(ram[15934]), .B2(n4120), 
        .ZN(n20175) );
  MOAI22 U29081 ( .A1(n27596), .A2(n4119), .B1(ram[15935]), .B2(n4120), 
        .ZN(n20176) );
  MOAI22 U29082 ( .A1(n29241), .A2(n4122), .B1(ram[15936]), .B2(n4123), 
        .ZN(n20177) );
  MOAI22 U29083 ( .A1(n29006), .A2(n4122), .B1(ram[15937]), .B2(n4123), 
        .ZN(n20178) );
  MOAI22 U29084 ( .A1(n28771), .A2(n4122), .B1(ram[15938]), .B2(n4123), 
        .ZN(n20179) );
  MOAI22 U29085 ( .A1(n28536), .A2(n4122), .B1(ram[15939]), .B2(n4123), 
        .ZN(n20180) );
  MOAI22 U29086 ( .A1(n28301), .A2(n4122), .B1(ram[15940]), .B2(n4123), 
        .ZN(n20181) );
  MOAI22 U29087 ( .A1(n28066), .A2(n4122), .B1(ram[15941]), .B2(n4123), 
        .ZN(n20182) );
  MOAI22 U29088 ( .A1(n27831), .A2(n4122), .B1(ram[15942]), .B2(n4123), 
        .ZN(n20183) );
  MOAI22 U29089 ( .A1(n27596), .A2(n4122), .B1(ram[15943]), .B2(n4123), 
        .ZN(n20184) );
  MOAI22 U29090 ( .A1(n29241), .A2(n4125), .B1(ram[15944]), .B2(n4126), 
        .ZN(n20185) );
  MOAI22 U29091 ( .A1(n29006), .A2(n4125), .B1(ram[15945]), .B2(n4126), 
        .ZN(n20186) );
  MOAI22 U29092 ( .A1(n28771), .A2(n4125), .B1(ram[15946]), .B2(n4126), 
        .ZN(n20187) );
  MOAI22 U29093 ( .A1(n28536), .A2(n4125), .B1(ram[15947]), .B2(n4126), 
        .ZN(n20188) );
  MOAI22 U29094 ( .A1(n28301), .A2(n4125), .B1(ram[15948]), .B2(n4126), 
        .ZN(n20189) );
  MOAI22 U29095 ( .A1(n28066), .A2(n4125), .B1(ram[15949]), .B2(n4126), 
        .ZN(n20190) );
  MOAI22 U29096 ( .A1(n27831), .A2(n4125), .B1(ram[15950]), .B2(n4126), 
        .ZN(n20191) );
  MOAI22 U29097 ( .A1(n27596), .A2(n4125), .B1(ram[15951]), .B2(n4126), 
        .ZN(n20192) );
  MOAI22 U29098 ( .A1(n29241), .A2(n4127), .B1(ram[15952]), .B2(n4128), 
        .ZN(n20193) );
  MOAI22 U29099 ( .A1(n29006), .A2(n4127), .B1(ram[15953]), .B2(n4128), 
        .ZN(n20194) );
  MOAI22 U29100 ( .A1(n28771), .A2(n4127), .B1(ram[15954]), .B2(n4128), 
        .ZN(n20195) );
  MOAI22 U29101 ( .A1(n28536), .A2(n4127), .B1(ram[15955]), .B2(n4128), 
        .ZN(n20196) );
  MOAI22 U29102 ( .A1(n28301), .A2(n4127), .B1(ram[15956]), .B2(n4128), 
        .ZN(n20197) );
  MOAI22 U29103 ( .A1(n28066), .A2(n4127), .B1(ram[15957]), .B2(n4128), 
        .ZN(n20198) );
  MOAI22 U29104 ( .A1(n27831), .A2(n4127), .B1(ram[15958]), .B2(n4128), 
        .ZN(n20199) );
  MOAI22 U29105 ( .A1(n27596), .A2(n4127), .B1(ram[15959]), .B2(n4128), 
        .ZN(n20200) );
  MOAI22 U29106 ( .A1(n29241), .A2(n4129), .B1(ram[15960]), .B2(n4130), 
        .ZN(n20201) );
  MOAI22 U29107 ( .A1(n29006), .A2(n4129), .B1(ram[15961]), .B2(n4130), 
        .ZN(n20202) );
  MOAI22 U29108 ( .A1(n28771), .A2(n4129), .B1(ram[15962]), .B2(n4130), 
        .ZN(n20203) );
  MOAI22 U29109 ( .A1(n28536), .A2(n4129), .B1(ram[15963]), .B2(n4130), 
        .ZN(n20204) );
  MOAI22 U29110 ( .A1(n28301), .A2(n4129), .B1(ram[15964]), .B2(n4130), 
        .ZN(n20205) );
  MOAI22 U29111 ( .A1(n28066), .A2(n4129), .B1(ram[15965]), .B2(n4130), 
        .ZN(n20206) );
  MOAI22 U29112 ( .A1(n27831), .A2(n4129), .B1(ram[15966]), .B2(n4130), 
        .ZN(n20207) );
  MOAI22 U29113 ( .A1(n27596), .A2(n4129), .B1(ram[15967]), .B2(n4130), 
        .ZN(n20208) );
  MOAI22 U29114 ( .A1(n29241), .A2(n4131), .B1(ram[15968]), .B2(n4132), 
        .ZN(n20209) );
  MOAI22 U29115 ( .A1(n29006), .A2(n4131), .B1(ram[15969]), .B2(n4132), 
        .ZN(n20210) );
  MOAI22 U29116 ( .A1(n28771), .A2(n4131), .B1(ram[15970]), .B2(n4132), 
        .ZN(n20211) );
  MOAI22 U29117 ( .A1(n28536), .A2(n4131), .B1(ram[15971]), .B2(n4132), 
        .ZN(n20212) );
  MOAI22 U29118 ( .A1(n28301), .A2(n4131), .B1(ram[15972]), .B2(n4132), 
        .ZN(n20213) );
  MOAI22 U29119 ( .A1(n28066), .A2(n4131), .B1(ram[15973]), .B2(n4132), 
        .ZN(n20214) );
  MOAI22 U29120 ( .A1(n27831), .A2(n4131), .B1(ram[15974]), .B2(n4132), 
        .ZN(n20215) );
  MOAI22 U29121 ( .A1(n27596), .A2(n4131), .B1(ram[15975]), .B2(n4132), 
        .ZN(n20216) );
  MOAI22 U29122 ( .A1(n29241), .A2(n4133), .B1(ram[15976]), .B2(n4134), 
        .ZN(n20217) );
  MOAI22 U29123 ( .A1(n29006), .A2(n4133), .B1(ram[15977]), .B2(n4134), 
        .ZN(n20218) );
  MOAI22 U29124 ( .A1(n28771), .A2(n4133), .B1(ram[15978]), .B2(n4134), 
        .ZN(n20219) );
  MOAI22 U29125 ( .A1(n28536), .A2(n4133), .B1(ram[15979]), .B2(n4134), 
        .ZN(n20220) );
  MOAI22 U29126 ( .A1(n28301), .A2(n4133), .B1(ram[15980]), .B2(n4134), 
        .ZN(n20221) );
  MOAI22 U29127 ( .A1(n28066), .A2(n4133), .B1(ram[15981]), .B2(n4134), 
        .ZN(n20222) );
  MOAI22 U29128 ( .A1(n27831), .A2(n4133), .B1(ram[15982]), .B2(n4134), 
        .ZN(n20223) );
  MOAI22 U29129 ( .A1(n27596), .A2(n4133), .B1(ram[15983]), .B2(n4134), 
        .ZN(n20224) );
  MOAI22 U29130 ( .A1(n29241), .A2(n4135), .B1(ram[15984]), .B2(n4136), 
        .ZN(n20225) );
  MOAI22 U29131 ( .A1(n29006), .A2(n4135), .B1(ram[15985]), .B2(n4136), 
        .ZN(n20226) );
  MOAI22 U29132 ( .A1(n28771), .A2(n4135), .B1(ram[15986]), .B2(n4136), 
        .ZN(n20227) );
  MOAI22 U29133 ( .A1(n28536), .A2(n4135), .B1(ram[15987]), .B2(n4136), 
        .ZN(n20228) );
  MOAI22 U29134 ( .A1(n28301), .A2(n4135), .B1(ram[15988]), .B2(n4136), 
        .ZN(n20229) );
  MOAI22 U29135 ( .A1(n28066), .A2(n4135), .B1(ram[15989]), .B2(n4136), 
        .ZN(n20230) );
  MOAI22 U29136 ( .A1(n27831), .A2(n4135), .B1(ram[15990]), .B2(n4136), 
        .ZN(n20231) );
  MOAI22 U29137 ( .A1(n27596), .A2(n4135), .B1(ram[15991]), .B2(n4136), 
        .ZN(n20232) );
  MOAI22 U29138 ( .A1(n29241), .A2(n4137), .B1(ram[15992]), .B2(n4138), 
        .ZN(n20233) );
  MOAI22 U29139 ( .A1(n29006), .A2(n4137), .B1(ram[15993]), .B2(n4138), 
        .ZN(n20234) );
  MOAI22 U29140 ( .A1(n28771), .A2(n4137), .B1(ram[15994]), .B2(n4138), 
        .ZN(n20235) );
  MOAI22 U29141 ( .A1(n28536), .A2(n4137), .B1(ram[15995]), .B2(n4138), 
        .ZN(n20236) );
  MOAI22 U29142 ( .A1(n28301), .A2(n4137), .B1(ram[15996]), .B2(n4138), 
        .ZN(n20237) );
  MOAI22 U29143 ( .A1(n28066), .A2(n4137), .B1(ram[15997]), .B2(n4138), 
        .ZN(n20238) );
  MOAI22 U29144 ( .A1(n27831), .A2(n4137), .B1(ram[15998]), .B2(n4138), 
        .ZN(n20239) );
  MOAI22 U29145 ( .A1(n27596), .A2(n4137), .B1(ram[15999]), .B2(n4138), 
        .ZN(n20240) );
  MOAI22 U29146 ( .A1(n29241), .A2(n4139), .B1(ram[16000]), .B2(n4140), 
        .ZN(n20241) );
  MOAI22 U29147 ( .A1(n29006), .A2(n4139), .B1(ram[16001]), .B2(n4140), 
        .ZN(n20242) );
  MOAI22 U29148 ( .A1(n28771), .A2(n4139), .B1(ram[16002]), .B2(n4140), 
        .ZN(n20243) );
  MOAI22 U29149 ( .A1(n28536), .A2(n4139), .B1(ram[16003]), .B2(n4140), 
        .ZN(n20244) );
  MOAI22 U29150 ( .A1(n28301), .A2(n4139), .B1(ram[16004]), .B2(n4140), 
        .ZN(n20245) );
  MOAI22 U29151 ( .A1(n28066), .A2(n4139), .B1(ram[16005]), .B2(n4140), 
        .ZN(n20246) );
  MOAI22 U29152 ( .A1(n27831), .A2(n4139), .B1(ram[16006]), .B2(n4140), 
        .ZN(n20247) );
  MOAI22 U29153 ( .A1(n27596), .A2(n4139), .B1(ram[16007]), .B2(n4140), 
        .ZN(n20248) );
  MOAI22 U29154 ( .A1(n29241), .A2(n4142), .B1(ram[16008]), .B2(n4143), 
        .ZN(n20249) );
  MOAI22 U29155 ( .A1(n29006), .A2(n4142), .B1(ram[16009]), .B2(n4143), 
        .ZN(n20250) );
  MOAI22 U29156 ( .A1(n28771), .A2(n4142), .B1(ram[16010]), .B2(n4143), 
        .ZN(n20251) );
  MOAI22 U29157 ( .A1(n28536), .A2(n4142), .B1(ram[16011]), .B2(n4143), 
        .ZN(n20252) );
  MOAI22 U29158 ( .A1(n28301), .A2(n4142), .B1(ram[16012]), .B2(n4143), 
        .ZN(n20253) );
  MOAI22 U29159 ( .A1(n28066), .A2(n4142), .B1(ram[16013]), .B2(n4143), 
        .ZN(n20254) );
  MOAI22 U29160 ( .A1(n27831), .A2(n4142), .B1(ram[16014]), .B2(n4143), 
        .ZN(n20255) );
  MOAI22 U29161 ( .A1(n27596), .A2(n4142), .B1(ram[16015]), .B2(n4143), 
        .ZN(n20256) );
  MOAI22 U29162 ( .A1(n29242), .A2(n4144), .B1(ram[16016]), .B2(n4145), 
        .ZN(n20257) );
  MOAI22 U29163 ( .A1(n29007), .A2(n4144), .B1(ram[16017]), .B2(n4145), 
        .ZN(n20258) );
  MOAI22 U29164 ( .A1(n28772), .A2(n4144), .B1(ram[16018]), .B2(n4145), 
        .ZN(n20259) );
  MOAI22 U29165 ( .A1(n28537), .A2(n4144), .B1(ram[16019]), .B2(n4145), 
        .ZN(n20260) );
  MOAI22 U29166 ( .A1(n28302), .A2(n4144), .B1(ram[16020]), .B2(n4145), 
        .ZN(n20261) );
  MOAI22 U29167 ( .A1(n28067), .A2(n4144), .B1(ram[16021]), .B2(n4145), 
        .ZN(n20262) );
  MOAI22 U29168 ( .A1(n27832), .A2(n4144), .B1(ram[16022]), .B2(n4145), 
        .ZN(n20263) );
  MOAI22 U29169 ( .A1(n27597), .A2(n4144), .B1(ram[16023]), .B2(n4145), 
        .ZN(n20264) );
  MOAI22 U29170 ( .A1(n29242), .A2(n4146), .B1(ram[16024]), .B2(n4147), 
        .ZN(n20265) );
  MOAI22 U29171 ( .A1(n29007), .A2(n4146), .B1(ram[16025]), .B2(n4147), 
        .ZN(n20266) );
  MOAI22 U29172 ( .A1(n28772), .A2(n4146), .B1(ram[16026]), .B2(n4147), 
        .ZN(n20267) );
  MOAI22 U29173 ( .A1(n28537), .A2(n4146), .B1(ram[16027]), .B2(n4147), 
        .ZN(n20268) );
  MOAI22 U29174 ( .A1(n28302), .A2(n4146), .B1(ram[16028]), .B2(n4147), 
        .ZN(n20269) );
  MOAI22 U29175 ( .A1(n28067), .A2(n4146), .B1(ram[16029]), .B2(n4147), 
        .ZN(n20270) );
  MOAI22 U29176 ( .A1(n27832), .A2(n4146), .B1(ram[16030]), .B2(n4147), 
        .ZN(n20271) );
  MOAI22 U29177 ( .A1(n27597), .A2(n4146), .B1(ram[16031]), .B2(n4147), 
        .ZN(n20272) );
  MOAI22 U29178 ( .A1(n29242), .A2(n4148), .B1(ram[16032]), .B2(n4149), 
        .ZN(n20273) );
  MOAI22 U29179 ( .A1(n29007), .A2(n4148), .B1(ram[16033]), .B2(n4149), 
        .ZN(n20274) );
  MOAI22 U29180 ( .A1(n28772), .A2(n4148), .B1(ram[16034]), .B2(n4149), 
        .ZN(n20275) );
  MOAI22 U29181 ( .A1(n28537), .A2(n4148), .B1(ram[16035]), .B2(n4149), 
        .ZN(n20276) );
  MOAI22 U29182 ( .A1(n28302), .A2(n4148), .B1(ram[16036]), .B2(n4149), 
        .ZN(n20277) );
  MOAI22 U29183 ( .A1(n28067), .A2(n4148), .B1(ram[16037]), .B2(n4149), 
        .ZN(n20278) );
  MOAI22 U29184 ( .A1(n27832), .A2(n4148), .B1(ram[16038]), .B2(n4149), 
        .ZN(n20279) );
  MOAI22 U29185 ( .A1(n27597), .A2(n4148), .B1(ram[16039]), .B2(n4149), 
        .ZN(n20280) );
  MOAI22 U29186 ( .A1(n29242), .A2(n4150), .B1(ram[16040]), .B2(n4151), 
        .ZN(n20281) );
  MOAI22 U29187 ( .A1(n29007), .A2(n4150), .B1(ram[16041]), .B2(n4151), 
        .ZN(n20282) );
  MOAI22 U29188 ( .A1(n28772), .A2(n4150), .B1(ram[16042]), .B2(n4151), 
        .ZN(n20283) );
  MOAI22 U29189 ( .A1(n28537), .A2(n4150), .B1(ram[16043]), .B2(n4151), 
        .ZN(n20284) );
  MOAI22 U29190 ( .A1(n28302), .A2(n4150), .B1(ram[16044]), .B2(n4151), 
        .ZN(n20285) );
  MOAI22 U29191 ( .A1(n28067), .A2(n4150), .B1(ram[16045]), .B2(n4151), 
        .ZN(n20286) );
  MOAI22 U29192 ( .A1(n27832), .A2(n4150), .B1(ram[16046]), .B2(n4151), 
        .ZN(n20287) );
  MOAI22 U29193 ( .A1(n27597), .A2(n4150), .B1(ram[16047]), .B2(n4151), 
        .ZN(n20288) );
  MOAI22 U29194 ( .A1(n29242), .A2(n4152), .B1(ram[16048]), .B2(n4153), 
        .ZN(n20289) );
  MOAI22 U29195 ( .A1(n29007), .A2(n4152), .B1(ram[16049]), .B2(n4153), 
        .ZN(n20290) );
  MOAI22 U29196 ( .A1(n28772), .A2(n4152), .B1(ram[16050]), .B2(n4153), 
        .ZN(n20291) );
  MOAI22 U29197 ( .A1(n28537), .A2(n4152), .B1(ram[16051]), .B2(n4153), 
        .ZN(n20292) );
  MOAI22 U29198 ( .A1(n28302), .A2(n4152), .B1(ram[16052]), .B2(n4153), 
        .ZN(n20293) );
  MOAI22 U29199 ( .A1(n28067), .A2(n4152), .B1(ram[16053]), .B2(n4153), 
        .ZN(n20294) );
  MOAI22 U29200 ( .A1(n27832), .A2(n4152), .B1(ram[16054]), .B2(n4153), 
        .ZN(n20295) );
  MOAI22 U29201 ( .A1(n27597), .A2(n4152), .B1(ram[16055]), .B2(n4153), 
        .ZN(n20296) );
  MOAI22 U29202 ( .A1(n29242), .A2(n4154), .B1(ram[16056]), .B2(n4155), 
        .ZN(n20297) );
  MOAI22 U29203 ( .A1(n29007), .A2(n4154), .B1(ram[16057]), .B2(n4155), 
        .ZN(n20298) );
  MOAI22 U29204 ( .A1(n28772), .A2(n4154), .B1(ram[16058]), .B2(n4155), 
        .ZN(n20299) );
  MOAI22 U29205 ( .A1(n28537), .A2(n4154), .B1(ram[16059]), .B2(n4155), 
        .ZN(n20300) );
  MOAI22 U29206 ( .A1(n28302), .A2(n4154), .B1(ram[16060]), .B2(n4155), 
        .ZN(n20301) );
  MOAI22 U29207 ( .A1(n28067), .A2(n4154), .B1(ram[16061]), .B2(n4155), 
        .ZN(n20302) );
  MOAI22 U29208 ( .A1(n27832), .A2(n4154), .B1(ram[16062]), .B2(n4155), 
        .ZN(n20303) );
  MOAI22 U29209 ( .A1(n27597), .A2(n4154), .B1(ram[16063]), .B2(n4155), 
        .ZN(n20304) );
  MOAI22 U29210 ( .A1(n29242), .A2(n4156), .B1(ram[16064]), .B2(n4157), 
        .ZN(n20305) );
  MOAI22 U29211 ( .A1(n29007), .A2(n4156), .B1(ram[16065]), .B2(n4157), 
        .ZN(n20306) );
  MOAI22 U29212 ( .A1(n28772), .A2(n4156), .B1(ram[16066]), .B2(n4157), 
        .ZN(n20307) );
  MOAI22 U29213 ( .A1(n28537), .A2(n4156), .B1(ram[16067]), .B2(n4157), 
        .ZN(n20308) );
  MOAI22 U29214 ( .A1(n28302), .A2(n4156), .B1(ram[16068]), .B2(n4157), 
        .ZN(n20309) );
  MOAI22 U29215 ( .A1(n28067), .A2(n4156), .B1(ram[16069]), .B2(n4157), 
        .ZN(n20310) );
  MOAI22 U29216 ( .A1(n27832), .A2(n4156), .B1(ram[16070]), .B2(n4157), 
        .ZN(n20311) );
  MOAI22 U29217 ( .A1(n27597), .A2(n4156), .B1(ram[16071]), .B2(n4157), 
        .ZN(n20312) );
  MOAI22 U29218 ( .A1(n29242), .A2(n4159), .B1(ram[16072]), .B2(n4160), 
        .ZN(n20313) );
  MOAI22 U29219 ( .A1(n29007), .A2(n4159), .B1(ram[16073]), .B2(n4160), 
        .ZN(n20314) );
  MOAI22 U29220 ( .A1(n28772), .A2(n4159), .B1(ram[16074]), .B2(n4160), 
        .ZN(n20315) );
  MOAI22 U29221 ( .A1(n28537), .A2(n4159), .B1(ram[16075]), .B2(n4160), 
        .ZN(n20316) );
  MOAI22 U29222 ( .A1(n28302), .A2(n4159), .B1(ram[16076]), .B2(n4160), 
        .ZN(n20317) );
  MOAI22 U29223 ( .A1(n28067), .A2(n4159), .B1(ram[16077]), .B2(n4160), 
        .ZN(n20318) );
  MOAI22 U29224 ( .A1(n27832), .A2(n4159), .B1(ram[16078]), .B2(n4160), 
        .ZN(n20319) );
  MOAI22 U29225 ( .A1(n27597), .A2(n4159), .B1(ram[16079]), .B2(n4160), 
        .ZN(n20320) );
  MOAI22 U29226 ( .A1(n29242), .A2(n4161), .B1(ram[16080]), .B2(n4162), 
        .ZN(n20321) );
  MOAI22 U29227 ( .A1(n29007), .A2(n4161), .B1(ram[16081]), .B2(n4162), 
        .ZN(n20322) );
  MOAI22 U29228 ( .A1(n28772), .A2(n4161), .B1(ram[16082]), .B2(n4162), 
        .ZN(n20323) );
  MOAI22 U29229 ( .A1(n28537), .A2(n4161), .B1(ram[16083]), .B2(n4162), 
        .ZN(n20324) );
  MOAI22 U29230 ( .A1(n28302), .A2(n4161), .B1(ram[16084]), .B2(n4162), 
        .ZN(n20325) );
  MOAI22 U29231 ( .A1(n28067), .A2(n4161), .B1(ram[16085]), .B2(n4162), 
        .ZN(n20326) );
  MOAI22 U29232 ( .A1(n27832), .A2(n4161), .B1(ram[16086]), .B2(n4162), 
        .ZN(n20327) );
  MOAI22 U29233 ( .A1(n27597), .A2(n4161), .B1(ram[16087]), .B2(n4162), 
        .ZN(n20328) );
  MOAI22 U29234 ( .A1(n29242), .A2(n4163), .B1(ram[16088]), .B2(n4164), 
        .ZN(n20329) );
  MOAI22 U29235 ( .A1(n29007), .A2(n4163), .B1(ram[16089]), .B2(n4164), 
        .ZN(n20330) );
  MOAI22 U29236 ( .A1(n28772), .A2(n4163), .B1(ram[16090]), .B2(n4164), 
        .ZN(n20331) );
  MOAI22 U29237 ( .A1(n28537), .A2(n4163), .B1(ram[16091]), .B2(n4164), 
        .ZN(n20332) );
  MOAI22 U29238 ( .A1(n28302), .A2(n4163), .B1(ram[16092]), .B2(n4164), 
        .ZN(n20333) );
  MOAI22 U29239 ( .A1(n28067), .A2(n4163), .B1(ram[16093]), .B2(n4164), 
        .ZN(n20334) );
  MOAI22 U29240 ( .A1(n27832), .A2(n4163), .B1(ram[16094]), .B2(n4164), 
        .ZN(n20335) );
  MOAI22 U29241 ( .A1(n27597), .A2(n4163), .B1(ram[16095]), .B2(n4164), 
        .ZN(n20336) );
  MOAI22 U29242 ( .A1(n29242), .A2(n4165), .B1(ram[16096]), .B2(n4166), 
        .ZN(n20337) );
  MOAI22 U29243 ( .A1(n29007), .A2(n4165), .B1(ram[16097]), .B2(n4166), 
        .ZN(n20338) );
  MOAI22 U29244 ( .A1(n28772), .A2(n4165), .B1(ram[16098]), .B2(n4166), 
        .ZN(n20339) );
  MOAI22 U29245 ( .A1(n28537), .A2(n4165), .B1(ram[16099]), .B2(n4166), 
        .ZN(n20340) );
  MOAI22 U29246 ( .A1(n28302), .A2(n4165), .B1(ram[16100]), .B2(n4166), 
        .ZN(n20341) );
  MOAI22 U29247 ( .A1(n28067), .A2(n4165), .B1(ram[16101]), .B2(n4166), 
        .ZN(n20342) );
  MOAI22 U29248 ( .A1(n27832), .A2(n4165), .B1(ram[16102]), .B2(n4166), 
        .ZN(n20343) );
  MOAI22 U29249 ( .A1(n27597), .A2(n4165), .B1(ram[16103]), .B2(n4166), 
        .ZN(n20344) );
  MOAI22 U29250 ( .A1(n29242), .A2(n4167), .B1(ram[16104]), .B2(n4168), 
        .ZN(n20345) );
  MOAI22 U29251 ( .A1(n29007), .A2(n4167), .B1(ram[16105]), .B2(n4168), 
        .ZN(n20346) );
  MOAI22 U29252 ( .A1(n28772), .A2(n4167), .B1(ram[16106]), .B2(n4168), 
        .ZN(n20347) );
  MOAI22 U29253 ( .A1(n28537), .A2(n4167), .B1(ram[16107]), .B2(n4168), 
        .ZN(n20348) );
  MOAI22 U29254 ( .A1(n28302), .A2(n4167), .B1(ram[16108]), .B2(n4168), 
        .ZN(n20349) );
  MOAI22 U29255 ( .A1(n28067), .A2(n4167), .B1(ram[16109]), .B2(n4168), 
        .ZN(n20350) );
  MOAI22 U29256 ( .A1(n27832), .A2(n4167), .B1(ram[16110]), .B2(n4168), 
        .ZN(n20351) );
  MOAI22 U29257 ( .A1(n27597), .A2(n4167), .B1(ram[16111]), .B2(n4168), 
        .ZN(n20352) );
  MOAI22 U29258 ( .A1(n29242), .A2(n4169), .B1(ram[16112]), .B2(n4170), 
        .ZN(n20353) );
  MOAI22 U29259 ( .A1(n29007), .A2(n4169), .B1(ram[16113]), .B2(n4170), 
        .ZN(n20354) );
  MOAI22 U29260 ( .A1(n28772), .A2(n4169), .B1(ram[16114]), .B2(n4170), 
        .ZN(n20355) );
  MOAI22 U29261 ( .A1(n28537), .A2(n4169), .B1(ram[16115]), .B2(n4170), 
        .ZN(n20356) );
  MOAI22 U29262 ( .A1(n28302), .A2(n4169), .B1(ram[16116]), .B2(n4170), 
        .ZN(n20357) );
  MOAI22 U29263 ( .A1(n28067), .A2(n4169), .B1(ram[16117]), .B2(n4170), 
        .ZN(n20358) );
  MOAI22 U29264 ( .A1(n27832), .A2(n4169), .B1(ram[16118]), .B2(n4170), 
        .ZN(n20359) );
  MOAI22 U29265 ( .A1(n27597), .A2(n4169), .B1(ram[16119]), .B2(n4170), 
        .ZN(n20360) );
  MOAI22 U29266 ( .A1(n29243), .A2(n4171), .B1(ram[16120]), .B2(n4172), 
        .ZN(n20361) );
  MOAI22 U29267 ( .A1(n29008), .A2(n4171), .B1(ram[16121]), .B2(n4172), 
        .ZN(n20362) );
  MOAI22 U29268 ( .A1(n28773), .A2(n4171), .B1(ram[16122]), .B2(n4172), 
        .ZN(n20363) );
  MOAI22 U29269 ( .A1(n28538), .A2(n4171), .B1(ram[16123]), .B2(n4172), 
        .ZN(n20364) );
  MOAI22 U29270 ( .A1(n28303), .A2(n4171), .B1(ram[16124]), .B2(n4172), 
        .ZN(n20365) );
  MOAI22 U29271 ( .A1(n28068), .A2(n4171), .B1(ram[16125]), .B2(n4172), 
        .ZN(n20366) );
  MOAI22 U29272 ( .A1(n27833), .A2(n4171), .B1(ram[16126]), .B2(n4172), 
        .ZN(n20367) );
  MOAI22 U29273 ( .A1(n27598), .A2(n4171), .B1(ram[16127]), .B2(n4172), 
        .ZN(n20368) );
  MOAI22 U29274 ( .A1(n29243), .A2(n4173), .B1(ram[16128]), .B2(n4174), 
        .ZN(n20369) );
  MOAI22 U29275 ( .A1(n29008), .A2(n4173), .B1(ram[16129]), .B2(n4174), 
        .ZN(n20370) );
  MOAI22 U29276 ( .A1(n28773), .A2(n4173), .B1(ram[16130]), .B2(n4174), 
        .ZN(n20371) );
  MOAI22 U29277 ( .A1(n28538), .A2(n4173), .B1(ram[16131]), .B2(n4174), 
        .ZN(n20372) );
  MOAI22 U29278 ( .A1(n28303), .A2(n4173), .B1(ram[16132]), .B2(n4174), 
        .ZN(n20373) );
  MOAI22 U29279 ( .A1(n28068), .A2(n4173), .B1(ram[16133]), .B2(n4174), 
        .ZN(n20374) );
  MOAI22 U29280 ( .A1(n27833), .A2(n4173), .B1(ram[16134]), .B2(n4174), 
        .ZN(n20375) );
  MOAI22 U29281 ( .A1(n27598), .A2(n4173), .B1(ram[16135]), .B2(n4174), 
        .ZN(n20376) );
  MOAI22 U29282 ( .A1(n29243), .A2(n4176), .B1(ram[16136]), .B2(n4177), 
        .ZN(n20377) );
  MOAI22 U29283 ( .A1(n29008), .A2(n4176), .B1(ram[16137]), .B2(n4177), 
        .ZN(n20378) );
  MOAI22 U29284 ( .A1(n28773), .A2(n4176), .B1(ram[16138]), .B2(n4177), 
        .ZN(n20379) );
  MOAI22 U29285 ( .A1(n28538), .A2(n4176), .B1(ram[16139]), .B2(n4177), 
        .ZN(n20380) );
  MOAI22 U29286 ( .A1(n28303), .A2(n4176), .B1(ram[16140]), .B2(n4177), 
        .ZN(n20381) );
  MOAI22 U29287 ( .A1(n28068), .A2(n4176), .B1(ram[16141]), .B2(n4177), 
        .ZN(n20382) );
  MOAI22 U29288 ( .A1(n27833), .A2(n4176), .B1(ram[16142]), .B2(n4177), 
        .ZN(n20383) );
  MOAI22 U29289 ( .A1(n27598), .A2(n4176), .B1(ram[16143]), .B2(n4177), 
        .ZN(n20384) );
  MOAI22 U29290 ( .A1(n29243), .A2(n4178), .B1(ram[16144]), .B2(n4179), 
        .ZN(n20385) );
  MOAI22 U29291 ( .A1(n29008), .A2(n4178), .B1(ram[16145]), .B2(n4179), 
        .ZN(n20386) );
  MOAI22 U29292 ( .A1(n28773), .A2(n4178), .B1(ram[16146]), .B2(n4179), 
        .ZN(n20387) );
  MOAI22 U29293 ( .A1(n28538), .A2(n4178), .B1(ram[16147]), .B2(n4179), 
        .ZN(n20388) );
  MOAI22 U29294 ( .A1(n28303), .A2(n4178), .B1(ram[16148]), .B2(n4179), 
        .ZN(n20389) );
  MOAI22 U29295 ( .A1(n28068), .A2(n4178), .B1(ram[16149]), .B2(n4179), 
        .ZN(n20390) );
  MOAI22 U29296 ( .A1(n27833), .A2(n4178), .B1(ram[16150]), .B2(n4179), 
        .ZN(n20391) );
  MOAI22 U29297 ( .A1(n27598), .A2(n4178), .B1(ram[16151]), .B2(n4179), 
        .ZN(n20392) );
  MOAI22 U29298 ( .A1(n29243), .A2(n4180), .B1(ram[16152]), .B2(n4181), 
        .ZN(n20393) );
  MOAI22 U29299 ( .A1(n29008), .A2(n4180), .B1(ram[16153]), .B2(n4181), 
        .ZN(n20394) );
  MOAI22 U29300 ( .A1(n28773), .A2(n4180), .B1(ram[16154]), .B2(n4181), 
        .ZN(n20395) );
  MOAI22 U29301 ( .A1(n28538), .A2(n4180), .B1(ram[16155]), .B2(n4181), 
        .ZN(n20396) );
  MOAI22 U29302 ( .A1(n28303), .A2(n4180), .B1(ram[16156]), .B2(n4181), 
        .ZN(n20397) );
  MOAI22 U29303 ( .A1(n28068), .A2(n4180), .B1(ram[16157]), .B2(n4181), 
        .ZN(n20398) );
  MOAI22 U29304 ( .A1(n27833), .A2(n4180), .B1(ram[16158]), .B2(n4181), 
        .ZN(n20399) );
  MOAI22 U29305 ( .A1(n27598), .A2(n4180), .B1(ram[16159]), .B2(n4181), 
        .ZN(n20400) );
  MOAI22 U29306 ( .A1(n29243), .A2(n4182), .B1(ram[16160]), .B2(n4183), 
        .ZN(n20401) );
  MOAI22 U29307 ( .A1(n29008), .A2(n4182), .B1(ram[16161]), .B2(n4183), 
        .ZN(n20402) );
  MOAI22 U29308 ( .A1(n28773), .A2(n4182), .B1(ram[16162]), .B2(n4183), 
        .ZN(n20403) );
  MOAI22 U29309 ( .A1(n28538), .A2(n4182), .B1(ram[16163]), .B2(n4183), 
        .ZN(n20404) );
  MOAI22 U29310 ( .A1(n28303), .A2(n4182), .B1(ram[16164]), .B2(n4183), 
        .ZN(n20405) );
  MOAI22 U29311 ( .A1(n28068), .A2(n4182), .B1(ram[16165]), .B2(n4183), 
        .ZN(n20406) );
  MOAI22 U29312 ( .A1(n27833), .A2(n4182), .B1(ram[16166]), .B2(n4183), 
        .ZN(n20407) );
  MOAI22 U29313 ( .A1(n27598), .A2(n4182), .B1(ram[16167]), .B2(n4183), 
        .ZN(n20408) );
  MOAI22 U29314 ( .A1(n29243), .A2(n4184), .B1(ram[16168]), .B2(n4185), 
        .ZN(n20409) );
  MOAI22 U29315 ( .A1(n29008), .A2(n4184), .B1(ram[16169]), .B2(n4185), 
        .ZN(n20410) );
  MOAI22 U29316 ( .A1(n28773), .A2(n4184), .B1(ram[16170]), .B2(n4185), 
        .ZN(n20411) );
  MOAI22 U29317 ( .A1(n28538), .A2(n4184), .B1(ram[16171]), .B2(n4185), 
        .ZN(n20412) );
  MOAI22 U29318 ( .A1(n28303), .A2(n4184), .B1(ram[16172]), .B2(n4185), 
        .ZN(n20413) );
  MOAI22 U29319 ( .A1(n28068), .A2(n4184), .B1(ram[16173]), .B2(n4185), 
        .ZN(n20414) );
  MOAI22 U29320 ( .A1(n27833), .A2(n4184), .B1(ram[16174]), .B2(n4185), 
        .ZN(n20415) );
  MOAI22 U29321 ( .A1(n27598), .A2(n4184), .B1(ram[16175]), .B2(n4185), 
        .ZN(n20416) );
  MOAI22 U29322 ( .A1(n29243), .A2(n4186), .B1(ram[16176]), .B2(n4187), 
        .ZN(n20417) );
  MOAI22 U29323 ( .A1(n29008), .A2(n4186), .B1(ram[16177]), .B2(n4187), 
        .ZN(n20418) );
  MOAI22 U29324 ( .A1(n28773), .A2(n4186), .B1(ram[16178]), .B2(n4187), 
        .ZN(n20419) );
  MOAI22 U29325 ( .A1(n28538), .A2(n4186), .B1(ram[16179]), .B2(n4187), 
        .ZN(n20420) );
  MOAI22 U29326 ( .A1(n28303), .A2(n4186), .B1(ram[16180]), .B2(n4187), 
        .ZN(n20421) );
  MOAI22 U29327 ( .A1(n28068), .A2(n4186), .B1(ram[16181]), .B2(n4187), 
        .ZN(n20422) );
  MOAI22 U29328 ( .A1(n27833), .A2(n4186), .B1(ram[16182]), .B2(n4187), 
        .ZN(n20423) );
  MOAI22 U29329 ( .A1(n27598), .A2(n4186), .B1(ram[16183]), .B2(n4187), 
        .ZN(n20424) );
  MOAI22 U29330 ( .A1(n29243), .A2(n4188), .B1(ram[16184]), .B2(n4189), 
        .ZN(n20425) );
  MOAI22 U29331 ( .A1(n29008), .A2(n4188), .B1(ram[16185]), .B2(n4189), 
        .ZN(n20426) );
  MOAI22 U29332 ( .A1(n28773), .A2(n4188), .B1(ram[16186]), .B2(n4189), 
        .ZN(n20427) );
  MOAI22 U29333 ( .A1(n28538), .A2(n4188), .B1(ram[16187]), .B2(n4189), 
        .ZN(n20428) );
  MOAI22 U29334 ( .A1(n28303), .A2(n4188), .B1(ram[16188]), .B2(n4189), 
        .ZN(n20429) );
  MOAI22 U29335 ( .A1(n28068), .A2(n4188), .B1(ram[16189]), .B2(n4189), 
        .ZN(n20430) );
  MOAI22 U29336 ( .A1(n27833), .A2(n4188), .B1(ram[16190]), .B2(n4189), 
        .ZN(n20431) );
  MOAI22 U29337 ( .A1(n27598), .A2(n4188), .B1(ram[16191]), .B2(n4189), 
        .ZN(n20432) );
  MOAI22 U29338 ( .A1(n29243), .A2(n4190), .B1(ram[16192]), .B2(n4191), 
        .ZN(n20433) );
  MOAI22 U29339 ( .A1(n29008), .A2(n4190), .B1(ram[16193]), .B2(n4191), 
        .ZN(n20434) );
  MOAI22 U29340 ( .A1(n28773), .A2(n4190), .B1(ram[16194]), .B2(n4191), 
        .ZN(n20435) );
  MOAI22 U29341 ( .A1(n28538), .A2(n4190), .B1(ram[16195]), .B2(n4191), 
        .ZN(n20436) );
  MOAI22 U29342 ( .A1(n28303), .A2(n4190), .B1(ram[16196]), .B2(n4191), 
        .ZN(n20437) );
  MOAI22 U29343 ( .A1(n28068), .A2(n4190), .B1(ram[16197]), .B2(n4191), 
        .ZN(n20438) );
  MOAI22 U29344 ( .A1(n27833), .A2(n4190), .B1(ram[16198]), .B2(n4191), 
        .ZN(n20439) );
  MOAI22 U29345 ( .A1(n27598), .A2(n4190), .B1(ram[16199]), .B2(n4191), 
        .ZN(n20440) );
  MOAI22 U29346 ( .A1(n29243), .A2(n4193), .B1(ram[16200]), .B2(n4194), 
        .ZN(n20441) );
  MOAI22 U29347 ( .A1(n29008), .A2(n4193), .B1(ram[16201]), .B2(n4194), 
        .ZN(n20442) );
  MOAI22 U29348 ( .A1(n28773), .A2(n4193), .B1(ram[16202]), .B2(n4194), 
        .ZN(n20443) );
  MOAI22 U29349 ( .A1(n28538), .A2(n4193), .B1(ram[16203]), .B2(n4194), 
        .ZN(n20444) );
  MOAI22 U29350 ( .A1(n28303), .A2(n4193), .B1(ram[16204]), .B2(n4194), 
        .ZN(n20445) );
  MOAI22 U29351 ( .A1(n28068), .A2(n4193), .B1(ram[16205]), .B2(n4194), 
        .ZN(n20446) );
  MOAI22 U29352 ( .A1(n27833), .A2(n4193), .B1(ram[16206]), .B2(n4194), 
        .ZN(n20447) );
  MOAI22 U29353 ( .A1(n27598), .A2(n4193), .B1(ram[16207]), .B2(n4194), 
        .ZN(n20448) );
  MOAI22 U29354 ( .A1(n29243), .A2(n4195), .B1(ram[16208]), .B2(n4196), 
        .ZN(n20449) );
  MOAI22 U29355 ( .A1(n29008), .A2(n4195), .B1(ram[16209]), .B2(n4196), 
        .ZN(n20450) );
  MOAI22 U29356 ( .A1(n28773), .A2(n4195), .B1(ram[16210]), .B2(n4196), 
        .ZN(n20451) );
  MOAI22 U29357 ( .A1(n28538), .A2(n4195), .B1(ram[16211]), .B2(n4196), 
        .ZN(n20452) );
  MOAI22 U29358 ( .A1(n28303), .A2(n4195), .B1(ram[16212]), .B2(n4196), 
        .ZN(n20453) );
  MOAI22 U29359 ( .A1(n28068), .A2(n4195), .B1(ram[16213]), .B2(n4196), 
        .ZN(n20454) );
  MOAI22 U29360 ( .A1(n27833), .A2(n4195), .B1(ram[16214]), .B2(n4196), 
        .ZN(n20455) );
  MOAI22 U29361 ( .A1(n27598), .A2(n4195), .B1(ram[16215]), .B2(n4196), 
        .ZN(n20456) );
  MOAI22 U29362 ( .A1(n29243), .A2(n4197), .B1(ram[16216]), .B2(n4198), 
        .ZN(n20457) );
  MOAI22 U29363 ( .A1(n29008), .A2(n4197), .B1(ram[16217]), .B2(n4198), 
        .ZN(n20458) );
  MOAI22 U29364 ( .A1(n28773), .A2(n4197), .B1(ram[16218]), .B2(n4198), 
        .ZN(n20459) );
  MOAI22 U29365 ( .A1(n28538), .A2(n4197), .B1(ram[16219]), .B2(n4198), 
        .ZN(n20460) );
  MOAI22 U29366 ( .A1(n28303), .A2(n4197), .B1(ram[16220]), .B2(n4198), 
        .ZN(n20461) );
  MOAI22 U29367 ( .A1(n28068), .A2(n4197), .B1(ram[16221]), .B2(n4198), 
        .ZN(n20462) );
  MOAI22 U29368 ( .A1(n27833), .A2(n4197), .B1(ram[16222]), .B2(n4198), 
        .ZN(n20463) );
  MOAI22 U29369 ( .A1(n27598), .A2(n4197), .B1(ram[16223]), .B2(n4198), 
        .ZN(n20464) );
  MOAI22 U29370 ( .A1(n29244), .A2(n4199), .B1(ram[16224]), .B2(n4200), 
        .ZN(n20465) );
  MOAI22 U29371 ( .A1(n29009), .A2(n4199), .B1(ram[16225]), .B2(n4200), 
        .ZN(n20466) );
  MOAI22 U29372 ( .A1(n28774), .A2(n4199), .B1(ram[16226]), .B2(n4200), 
        .ZN(n20467) );
  MOAI22 U29373 ( .A1(n28539), .A2(n4199), .B1(ram[16227]), .B2(n4200), 
        .ZN(n20468) );
  MOAI22 U29374 ( .A1(n28304), .A2(n4199), .B1(ram[16228]), .B2(n4200), 
        .ZN(n20469) );
  MOAI22 U29375 ( .A1(n28069), .A2(n4199), .B1(ram[16229]), .B2(n4200), 
        .ZN(n20470) );
  MOAI22 U29376 ( .A1(n27834), .A2(n4199), .B1(ram[16230]), .B2(n4200), 
        .ZN(n20471) );
  MOAI22 U29377 ( .A1(n27599), .A2(n4199), .B1(ram[16231]), .B2(n4200), 
        .ZN(n20472) );
  MOAI22 U29378 ( .A1(n29244), .A2(n4201), .B1(ram[16232]), .B2(n4202), 
        .ZN(n20473) );
  MOAI22 U29379 ( .A1(n29009), .A2(n4201), .B1(ram[16233]), .B2(n4202), 
        .ZN(n20474) );
  MOAI22 U29380 ( .A1(n28774), .A2(n4201), .B1(ram[16234]), .B2(n4202), 
        .ZN(n20475) );
  MOAI22 U29381 ( .A1(n28539), .A2(n4201), .B1(ram[16235]), .B2(n4202), 
        .ZN(n20476) );
  MOAI22 U29382 ( .A1(n28304), .A2(n4201), .B1(ram[16236]), .B2(n4202), 
        .ZN(n20477) );
  MOAI22 U29383 ( .A1(n28069), .A2(n4201), .B1(ram[16237]), .B2(n4202), 
        .ZN(n20478) );
  MOAI22 U29384 ( .A1(n27834), .A2(n4201), .B1(ram[16238]), .B2(n4202), 
        .ZN(n20479) );
  MOAI22 U29385 ( .A1(n27599), .A2(n4201), .B1(ram[16239]), .B2(n4202), 
        .ZN(n20480) );
  MOAI22 U29386 ( .A1(n29244), .A2(n4203), .B1(ram[16240]), .B2(n4204), 
        .ZN(n20481) );
  MOAI22 U29387 ( .A1(n29009), .A2(n4203), .B1(ram[16241]), .B2(n4204), 
        .ZN(n20482) );
  MOAI22 U29388 ( .A1(n28774), .A2(n4203), .B1(ram[16242]), .B2(n4204), 
        .ZN(n20483) );
  MOAI22 U29389 ( .A1(n28539), .A2(n4203), .B1(ram[16243]), .B2(n4204), 
        .ZN(n20484) );
  MOAI22 U29390 ( .A1(n28304), .A2(n4203), .B1(ram[16244]), .B2(n4204), 
        .ZN(n20485) );
  MOAI22 U29391 ( .A1(n28069), .A2(n4203), .B1(ram[16245]), .B2(n4204), 
        .ZN(n20486) );
  MOAI22 U29392 ( .A1(n27834), .A2(n4203), .B1(ram[16246]), .B2(n4204), 
        .ZN(n20487) );
  MOAI22 U29393 ( .A1(n27599), .A2(n4203), .B1(ram[16247]), .B2(n4204), 
        .ZN(n20488) );
  MOAI22 U29394 ( .A1(n29244), .A2(n4205), .B1(ram[16248]), .B2(n4206), 
        .ZN(n20489) );
  MOAI22 U29395 ( .A1(n29009), .A2(n4205), .B1(ram[16249]), .B2(n4206), 
        .ZN(n20490) );
  MOAI22 U29396 ( .A1(n28774), .A2(n4205), .B1(ram[16250]), .B2(n4206), 
        .ZN(n20491) );
  MOAI22 U29397 ( .A1(n28539), .A2(n4205), .B1(ram[16251]), .B2(n4206), 
        .ZN(n20492) );
  MOAI22 U29398 ( .A1(n28304), .A2(n4205), .B1(ram[16252]), .B2(n4206), 
        .ZN(n20493) );
  MOAI22 U29399 ( .A1(n28069), .A2(n4205), .B1(ram[16253]), .B2(n4206), 
        .ZN(n20494) );
  MOAI22 U29400 ( .A1(n27834), .A2(n4205), .B1(ram[16254]), .B2(n4206), 
        .ZN(n20495) );
  MOAI22 U29401 ( .A1(n27599), .A2(n4205), .B1(ram[16255]), .B2(n4206), 
        .ZN(n20496) );
  MOAI22 U29402 ( .A1(n29244), .A2(n4207), .B1(ram[16256]), .B2(n4208), 
        .ZN(n20497) );
  MOAI22 U29403 ( .A1(n29009), .A2(n4207), .B1(ram[16257]), .B2(n4208), 
        .ZN(n20498) );
  MOAI22 U29404 ( .A1(n28774), .A2(n4207), .B1(ram[16258]), .B2(n4208), 
        .ZN(n20499) );
  MOAI22 U29405 ( .A1(n28539), .A2(n4207), .B1(ram[16259]), .B2(n4208), 
        .ZN(n20500) );
  MOAI22 U29406 ( .A1(n28304), .A2(n4207), .B1(ram[16260]), .B2(n4208), 
        .ZN(n20501) );
  MOAI22 U29407 ( .A1(n28069), .A2(n4207), .B1(ram[16261]), .B2(n4208), 
        .ZN(n20502) );
  MOAI22 U29408 ( .A1(n27834), .A2(n4207), .B1(ram[16262]), .B2(n4208), 
        .ZN(n20503) );
  MOAI22 U29409 ( .A1(n27599), .A2(n4207), .B1(ram[16263]), .B2(n4208), 
        .ZN(n20504) );
  MOAI22 U29410 ( .A1(n29244), .A2(n4210), .B1(ram[16264]), .B2(n4211), 
        .ZN(n20505) );
  MOAI22 U29411 ( .A1(n29009), .A2(n4210), .B1(ram[16265]), .B2(n4211), 
        .ZN(n20506) );
  MOAI22 U29412 ( .A1(n28774), .A2(n4210), .B1(ram[16266]), .B2(n4211), 
        .ZN(n20507) );
  MOAI22 U29413 ( .A1(n28539), .A2(n4210), .B1(ram[16267]), .B2(n4211), 
        .ZN(n20508) );
  MOAI22 U29414 ( .A1(n28304), .A2(n4210), .B1(ram[16268]), .B2(n4211), 
        .ZN(n20509) );
  MOAI22 U29415 ( .A1(n28069), .A2(n4210), .B1(ram[16269]), .B2(n4211), 
        .ZN(n20510) );
  MOAI22 U29416 ( .A1(n27834), .A2(n4210), .B1(ram[16270]), .B2(n4211), 
        .ZN(n20511) );
  MOAI22 U29417 ( .A1(n27599), .A2(n4210), .B1(ram[16271]), .B2(n4211), 
        .ZN(n20512) );
  MOAI22 U29418 ( .A1(n29244), .A2(n4212), .B1(ram[16272]), .B2(n4213), 
        .ZN(n20513) );
  MOAI22 U29419 ( .A1(n29009), .A2(n4212), .B1(ram[16273]), .B2(n4213), 
        .ZN(n20514) );
  MOAI22 U29420 ( .A1(n28774), .A2(n4212), .B1(ram[16274]), .B2(n4213), 
        .ZN(n20515) );
  MOAI22 U29421 ( .A1(n28539), .A2(n4212), .B1(ram[16275]), .B2(n4213), 
        .ZN(n20516) );
  MOAI22 U29422 ( .A1(n28304), .A2(n4212), .B1(ram[16276]), .B2(n4213), 
        .ZN(n20517) );
  MOAI22 U29423 ( .A1(n28069), .A2(n4212), .B1(ram[16277]), .B2(n4213), 
        .ZN(n20518) );
  MOAI22 U29424 ( .A1(n27834), .A2(n4212), .B1(ram[16278]), .B2(n4213), 
        .ZN(n20519) );
  MOAI22 U29425 ( .A1(n27599), .A2(n4212), .B1(ram[16279]), .B2(n4213), 
        .ZN(n20520) );
  MOAI22 U29426 ( .A1(n29244), .A2(n4214), .B1(ram[16280]), .B2(n4215), 
        .ZN(n20521) );
  MOAI22 U29427 ( .A1(n29009), .A2(n4214), .B1(ram[16281]), .B2(n4215), 
        .ZN(n20522) );
  MOAI22 U29428 ( .A1(n28774), .A2(n4214), .B1(ram[16282]), .B2(n4215), 
        .ZN(n20523) );
  MOAI22 U29429 ( .A1(n28539), .A2(n4214), .B1(ram[16283]), .B2(n4215), 
        .ZN(n20524) );
  MOAI22 U29430 ( .A1(n28304), .A2(n4214), .B1(ram[16284]), .B2(n4215), 
        .ZN(n20525) );
  MOAI22 U29431 ( .A1(n28069), .A2(n4214), .B1(ram[16285]), .B2(n4215), 
        .ZN(n20526) );
  MOAI22 U29432 ( .A1(n27834), .A2(n4214), .B1(ram[16286]), .B2(n4215), 
        .ZN(n20527) );
  MOAI22 U29433 ( .A1(n27599), .A2(n4214), .B1(ram[16287]), .B2(n4215), 
        .ZN(n20528) );
  MOAI22 U29434 ( .A1(n29244), .A2(n4216), .B1(ram[16288]), .B2(n4217), 
        .ZN(n20529) );
  MOAI22 U29435 ( .A1(n29009), .A2(n4216), .B1(ram[16289]), .B2(n4217), 
        .ZN(n20530) );
  MOAI22 U29436 ( .A1(n28774), .A2(n4216), .B1(ram[16290]), .B2(n4217), 
        .ZN(n20531) );
  MOAI22 U29437 ( .A1(n28539), .A2(n4216), .B1(ram[16291]), .B2(n4217), 
        .ZN(n20532) );
  MOAI22 U29438 ( .A1(n28304), .A2(n4216), .B1(ram[16292]), .B2(n4217), 
        .ZN(n20533) );
  MOAI22 U29439 ( .A1(n28069), .A2(n4216), .B1(ram[16293]), .B2(n4217), 
        .ZN(n20534) );
  MOAI22 U29440 ( .A1(n27834), .A2(n4216), .B1(ram[16294]), .B2(n4217), 
        .ZN(n20535) );
  MOAI22 U29441 ( .A1(n27599), .A2(n4216), .B1(ram[16295]), .B2(n4217), 
        .ZN(n20536) );
  MOAI22 U29442 ( .A1(n29244), .A2(n4218), .B1(ram[16296]), .B2(n4219), 
        .ZN(n20537) );
  MOAI22 U29443 ( .A1(n29009), .A2(n4218), .B1(ram[16297]), .B2(n4219), 
        .ZN(n20538) );
  MOAI22 U29444 ( .A1(n28774), .A2(n4218), .B1(ram[16298]), .B2(n4219), 
        .ZN(n20539) );
  MOAI22 U29445 ( .A1(n28539), .A2(n4218), .B1(ram[16299]), .B2(n4219), 
        .ZN(n20540) );
  MOAI22 U29446 ( .A1(n28304), .A2(n4218), .B1(ram[16300]), .B2(n4219), 
        .ZN(n20541) );
  MOAI22 U29447 ( .A1(n28069), .A2(n4218), .B1(ram[16301]), .B2(n4219), 
        .ZN(n20542) );
  MOAI22 U29448 ( .A1(n27834), .A2(n4218), .B1(ram[16302]), .B2(n4219), 
        .ZN(n20543) );
  MOAI22 U29449 ( .A1(n27599), .A2(n4218), .B1(ram[16303]), .B2(n4219), 
        .ZN(n20544) );
  MOAI22 U29450 ( .A1(n29244), .A2(n4220), .B1(ram[16304]), .B2(n4221), 
        .ZN(n20545) );
  MOAI22 U29451 ( .A1(n29009), .A2(n4220), .B1(ram[16305]), .B2(n4221), 
        .ZN(n20546) );
  MOAI22 U29452 ( .A1(n28774), .A2(n4220), .B1(ram[16306]), .B2(n4221), 
        .ZN(n20547) );
  MOAI22 U29453 ( .A1(n28539), .A2(n4220), .B1(ram[16307]), .B2(n4221), 
        .ZN(n20548) );
  MOAI22 U29454 ( .A1(n28304), .A2(n4220), .B1(ram[16308]), .B2(n4221), 
        .ZN(n20549) );
  MOAI22 U29455 ( .A1(n28069), .A2(n4220), .B1(ram[16309]), .B2(n4221), 
        .ZN(n20550) );
  MOAI22 U29456 ( .A1(n27834), .A2(n4220), .B1(ram[16310]), .B2(n4221), 
        .ZN(n20551) );
  MOAI22 U29457 ( .A1(n27599), .A2(n4220), .B1(ram[16311]), .B2(n4221), 
        .ZN(n20552) );
  MOAI22 U29458 ( .A1(n29244), .A2(n4222), .B1(ram[16312]), .B2(n4223), 
        .ZN(n20553) );
  MOAI22 U29459 ( .A1(n29009), .A2(n4222), .B1(ram[16313]), .B2(n4223), 
        .ZN(n20554) );
  MOAI22 U29460 ( .A1(n28774), .A2(n4222), .B1(ram[16314]), .B2(n4223), 
        .ZN(n20555) );
  MOAI22 U29461 ( .A1(n28539), .A2(n4222), .B1(ram[16315]), .B2(n4223), 
        .ZN(n20556) );
  MOAI22 U29462 ( .A1(n28304), .A2(n4222), .B1(ram[16316]), .B2(n4223), 
        .ZN(n20557) );
  MOAI22 U29463 ( .A1(n28069), .A2(n4222), .B1(ram[16317]), .B2(n4223), 
        .ZN(n20558) );
  MOAI22 U29464 ( .A1(n27834), .A2(n4222), .B1(ram[16318]), .B2(n4223), 
        .ZN(n20559) );
  MOAI22 U29465 ( .A1(n27599), .A2(n4222), .B1(ram[16319]), .B2(n4223), 
        .ZN(n20560) );
  MOAI22 U29466 ( .A1(n29244), .A2(n4224), .B1(ram[16320]), .B2(n4225), 
        .ZN(n20561) );
  MOAI22 U29467 ( .A1(n29009), .A2(n4224), .B1(ram[16321]), .B2(n4225), 
        .ZN(n20562) );
  MOAI22 U29468 ( .A1(n28774), .A2(n4224), .B1(ram[16322]), .B2(n4225), 
        .ZN(n20563) );
  MOAI22 U29469 ( .A1(n28539), .A2(n4224), .B1(ram[16323]), .B2(n4225), 
        .ZN(n20564) );
  MOAI22 U29470 ( .A1(n28304), .A2(n4224), .B1(ram[16324]), .B2(n4225), 
        .ZN(n20565) );
  MOAI22 U29471 ( .A1(n28069), .A2(n4224), .B1(ram[16325]), .B2(n4225), 
        .ZN(n20566) );
  MOAI22 U29472 ( .A1(n27834), .A2(n4224), .B1(ram[16326]), .B2(n4225), 
        .ZN(n20567) );
  MOAI22 U29473 ( .A1(n27599), .A2(n4224), .B1(ram[16327]), .B2(n4225), 
        .ZN(n20568) );
  MOAI22 U29474 ( .A1(n29245), .A2(n4227), .B1(ram[16328]), .B2(n4228), 
        .ZN(n20569) );
  MOAI22 U29475 ( .A1(n29010), .A2(n4227), .B1(ram[16329]), .B2(n4228), 
        .ZN(n20570) );
  MOAI22 U29476 ( .A1(n28775), .A2(n4227), .B1(ram[16330]), .B2(n4228), 
        .ZN(n20571) );
  MOAI22 U29477 ( .A1(n28540), .A2(n4227), .B1(ram[16331]), .B2(n4228), 
        .ZN(n20572) );
  MOAI22 U29478 ( .A1(n28305), .A2(n4227), .B1(ram[16332]), .B2(n4228), 
        .ZN(n20573) );
  MOAI22 U29479 ( .A1(n28070), .A2(n4227), .B1(ram[16333]), .B2(n4228), 
        .ZN(n20574) );
  MOAI22 U29480 ( .A1(n27835), .A2(n4227), .B1(ram[16334]), .B2(n4228), 
        .ZN(n20575) );
  MOAI22 U29481 ( .A1(n27600), .A2(n4227), .B1(ram[16335]), .B2(n4228), 
        .ZN(n20576) );
  MOAI22 U29482 ( .A1(n29245), .A2(n4229), .B1(ram[16336]), .B2(n4230), 
        .ZN(n20577) );
  MOAI22 U29483 ( .A1(n29010), .A2(n4229), .B1(ram[16337]), .B2(n4230), 
        .ZN(n20578) );
  MOAI22 U29484 ( .A1(n28775), .A2(n4229), .B1(ram[16338]), .B2(n4230), 
        .ZN(n20579) );
  MOAI22 U29485 ( .A1(n28540), .A2(n4229), .B1(ram[16339]), .B2(n4230), 
        .ZN(n20580) );
  MOAI22 U29486 ( .A1(n28305), .A2(n4229), .B1(ram[16340]), .B2(n4230), 
        .ZN(n20581) );
  MOAI22 U29487 ( .A1(n28070), .A2(n4229), .B1(ram[16341]), .B2(n4230), 
        .ZN(n20582) );
  MOAI22 U29488 ( .A1(n27835), .A2(n4229), .B1(ram[16342]), .B2(n4230), 
        .ZN(n20583) );
  MOAI22 U29489 ( .A1(n27600), .A2(n4229), .B1(ram[16343]), .B2(n4230), 
        .ZN(n20584) );
  MOAI22 U29490 ( .A1(n29245), .A2(n4231), .B1(ram[16344]), .B2(n4232), 
        .ZN(n20585) );
  MOAI22 U29491 ( .A1(n29010), .A2(n4231), .B1(ram[16345]), .B2(n4232), 
        .ZN(n20586) );
  MOAI22 U29492 ( .A1(n28775), .A2(n4231), .B1(ram[16346]), .B2(n4232), 
        .ZN(n20587) );
  MOAI22 U29493 ( .A1(n28540), .A2(n4231), .B1(ram[16347]), .B2(n4232), 
        .ZN(n20588) );
  MOAI22 U29494 ( .A1(n28305), .A2(n4231), .B1(ram[16348]), .B2(n4232), 
        .ZN(n20589) );
  MOAI22 U29495 ( .A1(n28070), .A2(n4231), .B1(ram[16349]), .B2(n4232), 
        .ZN(n20590) );
  MOAI22 U29496 ( .A1(n27835), .A2(n4231), .B1(ram[16350]), .B2(n4232), 
        .ZN(n20591) );
  MOAI22 U29497 ( .A1(n27600), .A2(n4231), .B1(ram[16351]), .B2(n4232), 
        .ZN(n20592) );
  MOAI22 U29498 ( .A1(n29245), .A2(n4233), .B1(ram[16352]), .B2(n4234), 
        .ZN(n20593) );
  MOAI22 U29499 ( .A1(n29010), .A2(n4233), .B1(ram[16353]), .B2(n4234), 
        .ZN(n20594) );
  MOAI22 U29500 ( .A1(n28775), .A2(n4233), .B1(ram[16354]), .B2(n4234), 
        .ZN(n20595) );
  MOAI22 U29501 ( .A1(n28540), .A2(n4233), .B1(ram[16355]), .B2(n4234), 
        .ZN(n20596) );
  MOAI22 U29502 ( .A1(n28305), .A2(n4233), .B1(ram[16356]), .B2(n4234), 
        .ZN(n20597) );
  MOAI22 U29503 ( .A1(n28070), .A2(n4233), .B1(ram[16357]), .B2(n4234), 
        .ZN(n20598) );
  MOAI22 U29504 ( .A1(n27835), .A2(n4233), .B1(ram[16358]), .B2(n4234), 
        .ZN(n20599) );
  MOAI22 U29505 ( .A1(n27600), .A2(n4233), .B1(ram[16359]), .B2(n4234), 
        .ZN(n20600) );
  MOAI22 U29506 ( .A1(n29245), .A2(n4235), .B1(ram[16360]), .B2(n4236), 
        .ZN(n20601) );
  MOAI22 U29507 ( .A1(n29010), .A2(n4235), .B1(ram[16361]), .B2(n4236), 
        .ZN(n20602) );
  MOAI22 U29508 ( .A1(n28775), .A2(n4235), .B1(ram[16362]), .B2(n4236), 
        .ZN(n20603) );
  MOAI22 U29509 ( .A1(n28540), .A2(n4235), .B1(ram[16363]), .B2(n4236), 
        .ZN(n20604) );
  MOAI22 U29510 ( .A1(n28305), .A2(n4235), .B1(ram[16364]), .B2(n4236), 
        .ZN(n20605) );
  MOAI22 U29511 ( .A1(n28070), .A2(n4235), .B1(ram[16365]), .B2(n4236), 
        .ZN(n20606) );
  MOAI22 U29512 ( .A1(n27835), .A2(n4235), .B1(ram[16366]), .B2(n4236), 
        .ZN(n20607) );
  MOAI22 U29513 ( .A1(n27600), .A2(n4235), .B1(ram[16367]), .B2(n4236), 
        .ZN(n20608) );
  MOAI22 U29514 ( .A1(n29245), .A2(n4237), .B1(ram[16368]), .B2(n4238), 
        .ZN(n20609) );
  MOAI22 U29515 ( .A1(n29010), .A2(n4237), .B1(ram[16369]), .B2(n4238), 
        .ZN(n20610) );
  MOAI22 U29516 ( .A1(n28775), .A2(n4237), .B1(ram[16370]), .B2(n4238), 
        .ZN(n20611) );
  MOAI22 U29517 ( .A1(n28540), .A2(n4237), .B1(ram[16371]), .B2(n4238), 
        .ZN(n20612) );
  MOAI22 U29518 ( .A1(n28305), .A2(n4237), .B1(ram[16372]), .B2(n4238), 
        .ZN(n20613) );
  MOAI22 U29519 ( .A1(n28070), .A2(n4237), .B1(ram[16373]), .B2(n4238), 
        .ZN(n20614) );
  MOAI22 U29520 ( .A1(n27835), .A2(n4237), .B1(ram[16374]), .B2(n4238), 
        .ZN(n20615) );
  MOAI22 U29521 ( .A1(n27600), .A2(n4237), .B1(ram[16375]), .B2(n4238), 
        .ZN(n20616) );
  BUF U29522 ( .I(raddr[5]), .Z(n29320) );
  BUF U29523 ( .I(raddr[4]), .Z(n29319) );
  INV U29524 ( .I(raddr[7]), .ZN(n26085) );
  INV U29525 ( .I(raddr[6]), .ZN(n26091) );
  NAND2 U29526 ( .A1(din[2]), .A2(n29493), .ZN(n17) );
  NAND2 U29527 ( .A1(din[5]), .A2(n29493), .ZN(n20) );
  NAND2 U29528 ( .A1(din[6]), .A2(n29493), .ZN(n21) );
  NAND2 U29529 ( .A1(din[0]), .A2(n29492), .ZN(n14) );
  NAND2 U29530 ( .A1(din[1]), .A2(n29492), .ZN(n16) );
  NAND2 U29531 ( .A1(din[3]), .A2(n29492), .ZN(n18) );
  NAND2 U29532 ( .A1(din[4]), .A2(n29492), .ZN(n19) );
  NAND2 U29533 ( .A1(din[7]), .A2(n29492), .ZN(n22) );
  MOAI22 U29534 ( .A1(n29127), .A2(n1123), .B1(ram[4088]), .B2(n1124), 
        .ZN(n8329) );
  MOAI22 U29535 ( .A1(n28892), .A2(n1123), .B1(ram[4089]), .B2(n1124), 
        .ZN(n8330) );
  MOAI22 U29536 ( .A1(n28657), .A2(n1123), .B1(ram[4090]), .B2(n1124), 
        .ZN(n8331) );
  MOAI22 U29537 ( .A1(n28422), .A2(n1123), .B1(ram[4091]), .B2(n1124), 
        .ZN(n8332) );
  MOAI22 U29538 ( .A1(n28187), .A2(n1123), .B1(ram[4092]), .B2(n1124), 
        .ZN(n8333) );
  MOAI22 U29539 ( .A1(n27952), .A2(n1123), .B1(ram[4093]), .B2(n1124), 
        .ZN(n8334) );
  MOAI22 U29540 ( .A1(n27717), .A2(n1123), .B1(ram[4094]), .B2(n1124), 
        .ZN(n8335) );
  MOAI22 U29541 ( .A1(n27482), .A2(n1123), .B1(ram[4095]), .B2(n1124), 
        .ZN(n8336) );
  MOAI22 U29542 ( .A1(n29166), .A2(n2157), .B1(ram[8184]), .B2(n2158), 
        .ZN(n12425) );
  MOAI22 U29543 ( .A1(n28931), .A2(n2157), .B1(ram[8185]), .B2(n2158), 
        .ZN(n12426) );
  MOAI22 U29544 ( .A1(n28696), .A2(n2157), .B1(ram[8186]), .B2(n2158), 
        .ZN(n12427) );
  MOAI22 U29545 ( .A1(n28461), .A2(n2157), .B1(ram[8187]), .B2(n2158), 
        .ZN(n12428) );
  MOAI22 U29546 ( .A1(n28226), .A2(n2157), .B1(ram[8188]), .B2(n2158), 
        .ZN(n12429) );
  MOAI22 U29547 ( .A1(n27991), .A2(n2157), .B1(ram[8189]), .B2(n2158), 
        .ZN(n12430) );
  MOAI22 U29548 ( .A1(n27756), .A2(n2157), .B1(ram[8190]), .B2(n2158), 
        .ZN(n12431) );
  MOAI22 U29549 ( .A1(n27521), .A2(n2157), .B1(ram[8191]), .B2(n2158), 
        .ZN(n12432) );
  MOAI22 U29550 ( .A1(n29206), .A2(n3190), .B1(ram[12280]), .B2(n3191), 
        .ZN(n16521) );
  MOAI22 U29551 ( .A1(n28971), .A2(n3190), .B1(ram[12281]), .B2(n3191), 
        .ZN(n16522) );
  MOAI22 U29552 ( .A1(n28736), .A2(n3190), .B1(ram[12282]), .B2(n3191), 
        .ZN(n16523) );
  MOAI22 U29553 ( .A1(n28501), .A2(n3190), .B1(ram[12283]), .B2(n3191), 
        .ZN(n16524) );
  MOAI22 U29554 ( .A1(n28266), .A2(n3190), .B1(ram[12284]), .B2(n3191), 
        .ZN(n16525) );
  MOAI22 U29555 ( .A1(n28031), .A2(n3190), .B1(ram[12285]), .B2(n3191), 
        .ZN(n16526) );
  MOAI22 U29556 ( .A1(n27796), .A2(n3190), .B1(ram[12286]), .B2(n3191), 
        .ZN(n16527) );
  MOAI22 U29557 ( .A1(n27561), .A2(n3190), .B1(ram[12287]), .B2(n3191), 
        .ZN(n16528) );
  MOAI22 U29558 ( .A1(n29245), .A2(n4239), .B1(ram[16376]), .B2(n4240), 
        .ZN(n20617) );
  MOAI22 U29559 ( .A1(n29010), .A2(n4239), .B1(ram[16377]), .B2(n4240), 
        .ZN(n20618) );
  MOAI22 U29560 ( .A1(n28775), .A2(n4239), .B1(ram[16378]), .B2(n4240), 
        .ZN(n20619) );
  MOAI22 U29561 ( .A1(n28540), .A2(n4239), .B1(ram[16379]), .B2(n4240), 
        .ZN(n20620) );
  MOAI22 U29562 ( .A1(n28305), .A2(n4239), .B1(ram[16380]), .B2(n4240), 
        .ZN(n20621) );
  MOAI22 U29563 ( .A1(n28070), .A2(n4239), .B1(ram[16381]), .B2(n4240), 
        .ZN(n20622) );
  MOAI22 U29564 ( .A1(n27835), .A2(n4239), .B1(ram[16382]), .B2(n4240), 
        .ZN(n20623) );
  MOAI22 U29565 ( .A1(n27600), .A2(n4239), .B1(ram[16383]), .B2(n4240), 
        .ZN(n20624) );
  BUF U29566 ( .I(raddr[8]), .Z(n29321) );
  MUX21 U29567 ( .I0(n20778), .I1(n20693), .S(n29321), .Z(n20783) );
  MUX21 U29568 ( .I0(n21120), .I1(n21035), .S(n29321), .Z(n21125) );
  MUX21 U29569 ( .I0(n21291), .I1(n21206), .S(n29321), .Z(n21296) );
  MUX21 U29570 ( .I0(n21462), .I1(n21377), .S(n29321), .Z(n21467) );
  MUX21 U29571 ( .I0(n21804), .I1(n21719), .S(n29321), .Z(n21809) );
  MUX21 U29572 ( .I0(n21975), .I1(n21890), .S(n29321), .Z(n21980) );
  MUX21 U29573 ( .I0(n22146), .I1(n22061), .S(n29321), .Z(n22151) );
  MUX21 U29574 ( .I0(n22488), .I1(n22403), .S(n29321), .Z(n22493) );
  MUX21 U29575 ( .I0(n22659), .I1(n22574), .S(raddr[8]), .Z(n22664) );
  MUX21 U29576 ( .I0(n22830), .I1(n22745), .S(n29321), .Z(n22835) );
  MUX21 U29577 ( .I0(n23172), .I1(n23087), .S(raddr[8]), .Z(n23177) );
  MUX21 U29578 ( .I0(n23343), .I1(n23258), .S(raddr[8]), .Z(n23348) );
  MUX21 U29579 ( .I0(n23514), .I1(n23429), .S(n29321), .Z(n23519) );
  MUX21 U29580 ( .I0(n23856), .I1(n23771), .S(raddr[8]), .Z(n23861) );
  MUX21 U29581 ( .I0(n24027), .I1(n23942), .S(raddr[8]), .Z(n24032) );
  MUX21 U29582 ( .I0(n24198), .I1(n24113), .S(n29321), .Z(n24203) );
  MUX21 U29583 ( .I0(n24540), .I1(n24455), .S(raddr[8]), .Z(n24545) );
  MUX21 U29584 ( .I0(n24711), .I1(n24626), .S(n29321), .Z(n24716) );
  MUX21 U29585 ( .I0(n24882), .I1(n24797), .S(n29321), .Z(n24887) );
  MUX21 U29586 ( .I0(n25224), .I1(n25139), .S(raddr[8]), .Z(n25229) );
  MUX21 U29587 ( .I0(n25395), .I1(n25310), .S(raddr[8]), .Z(n25400) );
  MUX21 U29588 ( .I0(n25566), .I1(n25481), .S(n29321), .Z(n25571) );
  MUX21 U29589 ( .I0(n25908), .I1(n25823), .S(n29321), .Z(n25913) );
  MUX21 U29590 ( .I0(n26079), .I1(n25994), .S(n29321), .Z(n26084) );
  INV U29591 ( .I(waddr[0]), .ZN(n29582) );
  INV U29592 ( .I(waddr[1]), .ZN(n29583) );
  INV U29593 ( .I(waddr[2]), .ZN(n29584) );
  INV U29594 ( .I(waddr[3]), .ZN(n29585) );
  INV U29595 ( .I(waddr[4]), .ZN(n29586) );
  INV U29596 ( .I(waddr[5]), .ZN(n29587) );
  INV U29597 ( .I(waddr[6]), .ZN(n29588) );
  INV U29598 ( .I(waddr[7]), .ZN(n29589) );
  INV U29599 ( .I(waddr[8]), .ZN(n29590) );
  INV U29600 ( .I(waddr[9]), .ZN(n29591) );
  INV U29601 ( .I(waddr[10]), .ZN(n29592) );
endmodule


module fifo_shift_ram ( clk, reset_n, ram_re, push, din, sel, dout );
  input [10:0] push;
  input [7:0] din;
  input [3:0] sel;
  output [7:0] dout;
  input clk, reset_n, ram_re;
  wire   N119, N120, N121, N122, N123, N124, N125, N126, N127, N128, N129,
         N142, N143, N144, N145, N146, N147, N148, N149, N150, N151, N152,
         N165, N166, N167, N168, N169, N170, N171, N172, N173, N174, N175,
         N188, N189, N190, N191, N192, N193, N194, N195, N196, N197, N198,
         N211, N212, N213, N214, N215, N216, N217, N218, N219, N220, N221,
         N234, N235, N236, N237, N238, N239, N240, N241, N242, N243, N244,
         N257, N258, N259, N260, N261, N262, N263, N264, N265, N266, N267,
         N280, N281, N282, N283, N284, N285, N286, N287, N288, N289, N290,
         N303, N304, N305, N306, N307, N308, N309, N310, N311, N312, N313,
         N326, N327, N328, N329, N330, N331, N332, N333, N334, N335, N336,
         N349, N350, N351, N352, N353, N354, N355, N356, N357, N358, N359,
         N539, N540, N541, N542, N543, N544, N545, N546, N547, N548, N549,
         N562, N563, N564, N565, N566, N567, N568, N569, N570, N571, N572,
         N585, N586, N587, N588, N589, N590, N591, N592, N593, N594, N595,
         N608, N609, N610, N611, N612, N613, N614, N615, N616, N617, N618,
         N631, N632, N633, N634, N635, N636, N637, N638, N639, N640, N641,
         N654, N655, N656, N657, N658, N659, N660, N661, N662, N663, N664,
         N677, N678, N679, N680, N681, N682, N683, N684, N685, N686, N687,
         N700, N701, N702, N703, N704, N705, N706, N707, N708, N709, N710,
         N723, N724, N725, N726, N727, N728, N729, N730, N731, N732, N733,
         N746, N747, N748, N749, N750, N751, N752, N753, N754, N755, N756,
         N769, N770, N771, N772, N773, N774, N775, N776, N777, N778, N779,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82,
         n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96,
         n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n296, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679;
  wire   [120:0] waddr;
  wire   [10:0] addra;
  wire   [120:0] raddr;
  wire   [10:0] addrb;

  DFF_RST waddr_reg_1__0_ ( .D(n632), .CP(clk), .CDN(n21), .Q(waddr[110])
         );
  DFF_RST waddr_reg_1__1_ ( .D(n631), .CP(clk), .CDN(n21), .Q(waddr[111])
         );
  DFF_RST waddr_reg_1__2_ ( .D(n630), .CP(clk), .CDN(n21), .Q(waddr[112])
         );
  DFF_RST waddr_reg_1__3_ ( .D(n629), .CP(clk), .CDN(n21), .Q(waddr[113])
         );
  DFF_RST waddr_reg_1__4_ ( .D(n628), .CP(clk), .CDN(n21), .Q(waddr[114])
         );
  DFF_RST waddr_reg_1__5_ ( .D(n627), .CP(clk), .CDN(n21), .Q(waddr[115])
         );
  DFF_RST waddr_reg_1__6_ ( .D(n626), .CP(clk), .CDN(n21), .Q(waddr[116])
         );
  DFF_RST waddr_reg_1__7_ ( .D(n625), .CP(clk), .CDN(n21), .Q(waddr[117])
         );
  DFF_RST waddr_reg_1__8_ ( .D(n624), .CP(clk), .CDN(n21), .Q(waddr[118])
         );
  DFF_RST waddr_reg_1__9_ ( .D(n623), .CP(clk), .CDN(n21), .Q(waddr[119])
         );
  DFF_RST waddr_reg_1__10_ ( .D(n622), .CP(clk), .CDN(n21), .Q(waddr[120])
         );
  DFF_RST waddr_reg_2__0_ ( .D(n621), .CP(clk), .CDN(n21), .Q(waddr[99]) );
  DFF_RST waddr_reg_2__1_ ( .D(n620), .CP(clk), .CDN(n21), .Q(waddr[100])
         );
  DFF_RST waddr_reg_2__2_ ( .D(n619), .CP(clk), .CDN(n22), .Q(waddr[101])
         );
  DFF_RST waddr_reg_2__3_ ( .D(n618), .CP(clk), .CDN(n22), .Q(waddr[102])
         );
  DFF_RST waddr_reg_2__4_ ( .D(n617), .CP(clk), .CDN(n22), .Q(waddr[103])
         );
  DFF_RST waddr_reg_2__5_ ( .D(n616), .CP(clk), .CDN(n22), .Q(waddr[104])
         );
  DFF_RST waddr_reg_2__7_ ( .D(n614), .CP(clk), .CDN(n22), .Q(waddr[106])
         );
  DFF_RST waddr_reg_2__8_ ( .D(n613), .CP(clk), .CDN(n22), .Q(waddr[107])
         );
  DFF_RST waddr_reg_2__9_ ( .D(n612), .CP(clk), .CDN(n22), .Q(waddr[108])
         );
  DFF_RST waddr_reg_2__10_ ( .D(n611), .CP(clk), .CDN(n22), .Q(waddr[109])
         );
  DFF_RST waddr_reg_3__0_ ( .D(n610), .CP(clk), .CDN(n22), .Q(waddr[88]) );
  DFF_RST waddr_reg_3__1_ ( .D(n609), .CP(clk), .CDN(n22), .Q(waddr[89]) );
  DFF_RST waddr_reg_3__2_ ( .D(n608), .CP(clk), .CDN(n22), .Q(waddr[90]) );
  DFF_RST waddr_reg_3__3_ ( .D(n607), .CP(clk), .CDN(n22), .Q(waddr[91]) );
  DFF_RST waddr_reg_3__4_ ( .D(n606), .CP(clk), .CDN(n22), .Q(waddr[92]) );
  DFF_RST waddr_reg_3__5_ ( .D(n605), .CP(clk), .CDN(n23), .Q(waddr[93]) );
  DFF_RST waddr_reg_3__6_ ( .D(n604), .CP(clk), .CDN(n23), .Q(waddr[94]) );
  DFF_RST waddr_reg_3__8_ ( .D(n602), .CP(clk), .CDN(n23), .Q(waddr[96]) );
  DFF_RST waddr_reg_3__9_ ( .D(n601), .CP(clk), .CDN(n23), .Q(waddr[97]) );
  DFF_RST waddr_reg_3__10_ ( .D(n600), .CP(clk), .CDN(n23), .Q(waddr[98])
         );
  DFF_RST waddr_reg_4__0_ ( .D(n599), .CP(clk), .CDN(n23), .Q(waddr[77]) );
  DFF_RST waddr_reg_4__1_ ( .D(n598), .CP(clk), .CDN(n23), .Q(waddr[78]) );
  DFF_RST waddr_reg_4__2_ ( .D(n597), .CP(clk), .CDN(n23), .Q(waddr[79]) );
  DFF_RST waddr_reg_4__3_ ( .D(n596), .CP(clk), .CDN(n23), .Q(waddr[80]) );
  DFF_RST waddr_reg_4__4_ ( .D(n595), .CP(clk), .CDN(n23), .Q(waddr[81]) );
  DFF_RST waddr_reg_4__5_ ( .D(n594), .CP(clk), .CDN(n23), .Q(waddr[82]) );
  DFF_RST waddr_reg_4__6_ ( .D(n593), .CP(clk), .CDN(n23), .Q(waddr[83]) );
  DFF_RST waddr_reg_4__7_ ( .D(n592), .CP(clk), .CDN(n23), .Q(waddr[84]) );
  DFF_RST waddr_reg_4__9_ ( .D(n590), .CP(clk), .CDN(n24), .Q(waddr[86]) );
  DFF_RST waddr_reg_4__10_ ( .D(n589), .CP(clk), .CDN(n24), .Q(waddr[87])
         );
  DFF_RST waddr_reg_5__0_ ( .D(n588), .CP(clk), .CDN(n24), .Q(waddr[66]) );
  DFF_RST waddr_reg_5__1_ ( .D(n587), .CP(clk), .CDN(n24), .Q(waddr[67]) );
  DFF_RST waddr_reg_5__2_ ( .D(n586), .CP(clk), .CDN(n24), .Q(waddr[68]) );
  DFF_RST waddr_reg_5__3_ ( .D(n585), .CP(clk), .CDN(n24), .Q(waddr[69]) );
  DFF_RST waddr_reg_5__4_ ( .D(n584), .CP(clk), .CDN(n24), .Q(waddr[70]) );
  DFF_RST waddr_reg_5__5_ ( .D(n583), .CP(clk), .CDN(n24), .Q(waddr[71]) );
  DFF_RST waddr_reg_5__6_ ( .D(n582), .CP(clk), .CDN(n24), .Q(waddr[72]) );
  DFF_RST waddr_reg_5__9_ ( .D(n579), .CP(clk), .CDN(n24), .Q(waddr[75]) );
  DFF_RST waddr_reg_5__10_ ( .D(n578), .CP(clk), .CDN(n24), .Q(waddr[76])
         );
  DFF_RST waddr_reg_6__0_ ( .D(n577), .CP(clk), .CDN(n24), .Q(waddr[55]) );
  DFF_RST waddr_reg_6__1_ ( .D(n576), .CP(clk), .CDN(n24), .Q(waddr[56]) );
  DFF_RST waddr_reg_6__2_ ( .D(n575), .CP(clk), .CDN(n25), .Q(waddr[57]) );
  DFF_RST waddr_reg_6__3_ ( .D(n574), .CP(clk), .CDN(n25), .Q(waddr[58]) );
  DFF_RST waddr_reg_6__4_ ( .D(n573), .CP(clk), .CDN(n25), .Q(waddr[59]) );
  DFF_RST waddr_reg_6__5_ ( .D(n572), .CP(clk), .CDN(n25), .Q(waddr[60]) );
  DFF_RST waddr_reg_6__6_ ( .D(n571), .CP(clk), .CDN(n25), .Q(waddr[61]) );
  DFF_RST waddr_reg_6__7_ ( .D(n570), .CP(clk), .CDN(n25), .Q(waddr[62]) );
  DFF_RST waddr_reg_6__8_ ( .D(n569), .CP(clk), .CDN(n25), .Q(waddr[63]) );
  DFF_RST waddr_reg_6__10_ ( .D(n567), .CP(clk), .CDN(n25), .Q(waddr[65])
         );
  DFF_RST waddr_reg_7__0_ ( .D(n566), .CP(clk), .CDN(n25), .Q(waddr[44]) );
  DFF_RST waddr_reg_7__1_ ( .D(n565), .CP(clk), .CDN(n25), .Q(waddr[45]) );
  DFF_RST waddr_reg_7__2_ ( .D(n564), .CP(clk), .CDN(n25), .Q(waddr[46]) );
  DFF_RST waddr_reg_7__3_ ( .D(n563), .CP(clk), .CDN(n25), .Q(waddr[47]) );
  DFF_RST waddr_reg_7__4_ ( .D(n562), .CP(clk), .CDN(n25), .Q(waddr[48]) );
  DFF_RST waddr_reg_7__5_ ( .D(n561), .CP(clk), .CDN(n26), .Q(waddr[49]) );
  DFF_RST waddr_reg_7__6_ ( .D(n560), .CP(clk), .CDN(n26), .Q(waddr[50]) );
  DFF_RST waddr_reg_7__8_ ( .D(n558), .CP(clk), .CDN(n26), .Q(waddr[52]) );
  DFF_RST waddr_reg_7__10_ ( .D(n556), .CP(clk), .CDN(n26), .Q(waddr[54])
         );
  DFF_RST waddr_reg_8__0_ ( .D(n555), .CP(clk), .CDN(n26), .Q(waddr[33]) );
  DFF_RST waddr_reg_8__1_ ( .D(n554), .CP(clk), .CDN(n26), .Q(waddr[34]) );
  DFF_RST waddr_reg_8__2_ ( .D(n553), .CP(clk), .CDN(n26), .Q(waddr[35]) );
  DFF_RST waddr_reg_8__3_ ( .D(n552), .CP(clk), .CDN(n26), .Q(waddr[36]) );
  DFF_RST waddr_reg_8__4_ ( .D(n551), .CP(clk), .CDN(n26), .Q(waddr[37]) );
  DFF_RST waddr_reg_8__5_ ( .D(n550), .CP(clk), .CDN(n26), .Q(waddr[38]) );
  DFF_RST waddr_reg_8__6_ ( .D(n549), .CP(clk), .CDN(n26), .Q(waddr[39]) );
  DFF_RST waddr_reg_8__7_ ( .D(n548), .CP(clk), .CDN(n26), .Q(waddr[40]) );
  DFF_RST waddr_reg_8__10_ ( .D(n545), .CP(clk), .CDN(n26), .Q(waddr[43])
         );
  DFF_RST waddr_reg_9__0_ ( .D(n544), .CP(clk), .CDN(n27), .Q(waddr[22]) );
  DFF_RST waddr_reg_9__1_ ( .D(n543), .CP(clk), .CDN(n27), .Q(waddr[23]) );
  DFF_RST waddr_reg_9__2_ ( .D(n542), .CP(clk), .CDN(n27), .Q(waddr[24]) );
  DFF_RST waddr_reg_9__3_ ( .D(n541), .CP(clk), .CDN(n27), .Q(waddr[25]) );
  DFF_RST waddr_reg_9__4_ ( .D(n540), .CP(clk), .CDN(n27), .Q(waddr[26]) );
  DFF_RST waddr_reg_9__5_ ( .D(n539), .CP(clk), .CDN(n27), .Q(waddr[27]) );
  DFF_RST waddr_reg_9__6_ ( .D(n538), .CP(clk), .CDN(n27), .Q(waddr[28]) );
  DFF_RST waddr_reg_9__7_ ( .D(n537), .CP(clk), .CDN(n27), .Q(waddr[29]) );
  DFF_RST waddr_reg_9__8_ ( .D(n536), .CP(clk), .CDN(n27), .Q(waddr[30]) );
  DFF_RST waddr_reg_9__9_ ( .D(n535), .CP(clk), .CDN(n27), .Q(waddr[31]) );
  DFF_RST waddr_reg_10__0_ ( .D(n533), .CP(clk), .CDN(n27), .Q(waddr[11])
         );
  DFF_RST waddr_reg_10__1_ ( .D(n532), .CP(clk), .CDN(n27), .Q(waddr[12])
         );
  DFF_RST waddr_reg_10__2_ ( .D(n531), .CP(clk), .CDN(n27), .Q(waddr[13])
         );
  DFF_RST waddr_reg_10__3_ ( .D(n530), .CP(clk), .CDN(n28), .Q(waddr[14])
         );
  DFF_RST waddr_reg_10__4_ ( .D(n529), .CP(clk), .CDN(n28), .Q(waddr[15])
         );
  DFF_RST waddr_reg_10__5_ ( .D(n528), .CP(clk), .CDN(n28), .Q(waddr[16])
         );
  DFF_RST waddr_reg_10__6_ ( .D(n527), .CP(clk), .CDN(n28), .Q(waddr[17])
         );
  DFF_RST waddr_reg_10__7_ ( .D(n526), .CP(clk), .CDN(n28), .Q(waddr[18])
         );
  DFF_RST waddr_reg_10__9_ ( .D(n524), .CP(clk), .CDN(n28), .Q(waddr[20])
         );
  DFF_RST waddr_reg_11__0_ ( .D(n522), .CP(clk), .CDN(n28), .Q(waddr[0]) );
  DFF_RST waddr_reg_11__1_ ( .D(n521), .CP(clk), .CDN(n28), .Q(waddr[1]) );
  DFF_RST waddr_reg_11__2_ ( .D(n520), .CP(clk), .CDN(n28), .Q(waddr[2]) );
  DFF_RST waddr_reg_11__3_ ( .D(n519), .CP(clk), .CDN(n28), .Q(waddr[3]) );
  DFF_RST waddr_reg_11__4_ ( .D(n518), .CP(clk), .CDN(n28), .Q(waddr[4]) );
  DFF_RST waddr_reg_11__5_ ( .D(n517), .CP(clk), .CDN(n28), .Q(waddr[5]) );
  DFF_RST waddr_reg_11__6_ ( .D(n516), .CP(clk), .CDN(n28), .Q(waddr[6]) );
  DFF_RST waddr_reg_11__7_ ( .D(n515), .CP(clk), .CDN(n29), .Q(waddr[7]) );
  DFF_RST waddr_reg_11__8_ ( .D(n514), .CP(clk), .CDN(n29), .Q(waddr[8]) );
  DFF_RST raddr_reg_1__0_ ( .D(n511), .CP(clk), .CDN(n29), .Q(raddr[110])
         );
  DFF_RST raddr_reg_1__1_ ( .D(n510), .CP(clk), .CDN(n29), .Q(raddr[111])
         );
  DFF_RST raddr_reg_1__2_ ( .D(n509), .CP(clk), .CDN(n29), .Q(raddr[112])
         );
  DFF_RST raddr_reg_1__3_ ( .D(n508), .CP(clk), .CDN(n29), .Q(raddr[113])
         );
  DFF_RST raddr_reg_1__4_ ( .D(n507), .CP(clk), .CDN(n29), .Q(raddr[114])
         );
  DFF_RST raddr_reg_1__5_ ( .D(n506), .CP(clk), .CDN(n29), .Q(raddr[115])
         );
  DFF_RST raddr_reg_1__6_ ( .D(n505), .CP(clk), .CDN(n29), .Q(raddr[116])
         );
  DFF_RST raddr_reg_1__7_ ( .D(n504), .CP(clk), .CDN(n29), .Q(raddr[117])
         );
  DFF_RST raddr_reg_1__8_ ( .D(n503), .CP(clk), .CDN(n29), .Q(raddr[118])
         );
  DFF_RST raddr_reg_1__9_ ( .D(n502), .CP(clk), .CDN(n29), .Q(raddr[119])
         );
  DFF_RST raddr_reg_1__10_ ( .D(n501), .CP(clk), .CDN(n29), .Q(raddr[120])
         );
  DFF_RST raddr_reg_2__0_ ( .D(n500), .CP(clk), .CDN(n30), .Q(raddr[99]) );
  DFF_RST raddr_reg_2__1_ ( .D(n499), .CP(clk), .CDN(n30), .Q(raddr[100])
         );
  DFF_RST raddr_reg_2__2_ ( .D(n498), .CP(clk), .CDN(n30), .Q(raddr[101])
         );
  DFF_RST raddr_reg_2__3_ ( .D(n497), .CP(clk), .CDN(n30), .Q(raddr[102])
         );
  DFF_RST raddr_reg_2__4_ ( .D(n496), .CP(clk), .CDN(n30), .Q(raddr[103])
         );
  DFF_RST raddr_reg_2__5_ ( .D(n495), .CP(clk), .CDN(n30), .Q(raddr[104])
         );
  DFF_RST raddr_reg_2__7_ ( .D(n493), .CP(clk), .CDN(n30), .Q(raddr[106])
         );
  DFF_RST raddr_reg_2__8_ ( .D(n492), .CP(clk), .CDN(n30), .Q(raddr[107])
         );
  DFF_RST raddr_reg_2__9_ ( .D(n491), .CP(clk), .CDN(n30), .Q(raddr[108])
         );
  DFF_RST raddr_reg_2__10_ ( .D(n490), .CP(clk), .CDN(n30), .Q(raddr[109])
         );
  DFF_RST raddr_reg_3__0_ ( .D(n489), .CP(clk), .CDN(n30), .Q(raddr[88]) );
  DFF_RST raddr_reg_3__1_ ( .D(n488), .CP(clk), .CDN(n30), .Q(raddr[89]) );
  DFF_RST raddr_reg_3__2_ ( .D(n487), .CP(clk), .CDN(n30), .Q(raddr[90]) );
  DFF_RST raddr_reg_3__3_ ( .D(n486), .CP(clk), .CDN(n31), .Q(raddr[91]) );
  DFF_RST raddr_reg_3__4_ ( .D(n485), .CP(clk), .CDN(n31), .Q(raddr[92]) );
  DFF_RST raddr_reg_3__5_ ( .D(n484), .CP(clk), .CDN(n31), .Q(raddr[93]) );
  DFF_RST raddr_reg_3__6_ ( .D(n483), .CP(clk), .CDN(n31), .Q(raddr[94]) );
  DFF_RST raddr_reg_3__8_ ( .D(n481), .CP(clk), .CDN(n31), .Q(raddr[96]) );
  DFF_RST raddr_reg_3__9_ ( .D(n480), .CP(clk), .CDN(n31), .Q(raddr[97]) );
  DFF_RST raddr_reg_3__10_ ( .D(n479), .CP(clk), .CDN(n31), .Q(raddr[98])
         );
  DFF_RST raddr_reg_4__0_ ( .D(n478), .CP(clk), .CDN(n31), .Q(raddr[77]) );
  DFF_RST raddr_reg_4__1_ ( .D(n477), .CP(clk), .CDN(n31), .Q(raddr[78]) );
  DFF_RST raddr_reg_4__2_ ( .D(n476), .CP(clk), .CDN(n31), .Q(raddr[79]) );
  DFF_RST raddr_reg_4__3_ ( .D(n475), .CP(clk), .CDN(n31), .Q(raddr[80]) );
  DFF_RST raddr_reg_4__4_ ( .D(n474), .CP(clk), .CDN(n31), .Q(raddr[81]) );
  DFF_RST raddr_reg_4__5_ ( .D(n473), .CP(clk), .CDN(n31), .Q(raddr[82]) );
  DFF_RST raddr_reg_4__6_ ( .D(n472), .CP(clk), .CDN(n32), .Q(raddr[83]) );
  DFF_RST raddr_reg_4__7_ ( .D(n471), .CP(clk), .CDN(n32), .Q(raddr[84]) );
  DFF_RST raddr_reg_4__9_ ( .D(n469), .CP(clk), .CDN(n32), .Q(raddr[86]) );
  DFF_RST raddr_reg_4__10_ ( .D(n468), .CP(clk), .CDN(n32), .Q(raddr[87])
         );
  DFF_RST raddr_reg_5__0_ ( .D(n467), .CP(clk), .CDN(n32), .Q(raddr[66]) );
  DFF_RST raddr_reg_5__1_ ( .D(n466), .CP(clk), .CDN(n32), .Q(raddr[67]) );
  DFF_RST raddr_reg_5__2_ ( .D(n465), .CP(clk), .CDN(n32), .Q(raddr[68]) );
  DFF_RST raddr_reg_5__3_ ( .D(n464), .CP(clk), .CDN(n32), .Q(raddr[69]) );
  DFF_RST raddr_reg_5__4_ ( .D(n463), .CP(clk), .CDN(n32), .Q(raddr[70]) );
  DFF_RST raddr_reg_5__5_ ( .D(n462), .CP(clk), .CDN(n32), .Q(raddr[71]) );
  DFF_RST raddr_reg_5__6_ ( .D(n461), .CP(clk), .CDN(n32), .Q(raddr[72]) );
  DFF_RST raddr_reg_5__9_ ( .D(n458), .CP(clk), .CDN(n32), .Q(raddr[75]) );
  DFF_RST raddr_reg_5__10_ ( .D(n457), .CP(clk), .CDN(n32), .Q(raddr[76])
         );
  DFF_RST raddr_reg_6__0_ ( .D(n456), .CP(clk), .CDN(n33), .Q(raddr[55]) );
  DFF_RST raddr_reg_6__1_ ( .D(n455), .CP(clk), .CDN(n33), .Q(raddr[56]) );
  DFF_RST raddr_reg_6__2_ ( .D(n454), .CP(clk), .CDN(n33), .Q(raddr[57]) );
  DFF_RST raddr_reg_6__3_ ( .D(n453), .CP(clk), .CDN(n33), .Q(raddr[58]) );
  DFF_RST raddr_reg_6__4_ ( .D(n452), .CP(clk), .CDN(n33), .Q(raddr[59]) );
  DFF_RST raddr_reg_6__5_ ( .D(n451), .CP(clk), .CDN(n33), .Q(raddr[60]) );
  DFF_RST raddr_reg_6__6_ ( .D(n450), .CP(clk), .CDN(n33), .Q(raddr[61]) );
  DFF_RST raddr_reg_6__7_ ( .D(n449), .CP(clk), .CDN(n33), .Q(raddr[62]) );
  DFF_RST raddr_reg_6__8_ ( .D(n448), .CP(clk), .CDN(n33), .Q(raddr[63]) );
  DFF_RST raddr_reg_6__10_ ( .D(n446), .CP(clk), .CDN(n33), .Q(raddr[65])
         );
  DFF_RST raddr_reg_7__0_ ( .D(n445), .CP(clk), .CDN(n33), .Q(raddr[44]) );
  DFF_RST raddr_reg_7__1_ ( .D(n444), .CP(clk), .CDN(n33), .Q(raddr[45]) );
  DFF_RST raddr_reg_7__2_ ( .D(n443), .CP(clk), .CDN(n33), .Q(raddr[46]) );
  DFF_RST raddr_reg_7__3_ ( .D(n442), .CP(clk), .CDN(n34), .Q(raddr[47]) );
  DFF_RST raddr_reg_7__4_ ( .D(n441), .CP(clk), .CDN(n34), .Q(raddr[48]) );
  DFF_RST raddr_reg_7__5_ ( .D(n440), .CP(clk), .CDN(n34), .Q(raddr[49]) );
  DFF_RST raddr_reg_7__6_ ( .D(n439), .CP(clk), .CDN(n34), .Q(raddr[50]) );
  DFF_RST raddr_reg_7__8_ ( .D(n437), .CP(clk), .CDN(n34), .Q(raddr[52]) );
  DFF_RST raddr_reg_7__10_ ( .D(n435), .CP(clk), .CDN(n34), .Q(raddr[54])
         );
  DFF_RST raddr_reg_8__0_ ( .D(n434), .CP(clk), .CDN(n34), .Q(raddr[33]) );
  DFF_RST raddr_reg_8__1_ ( .D(n433), .CP(clk), .CDN(n34), .Q(raddr[34]) );
  DFF_RST raddr_reg_8__2_ ( .D(n432), .CP(clk), .CDN(n34), .Q(raddr[35]) );
  DFF_RST raddr_reg_8__3_ ( .D(n431), .CP(clk), .CDN(n34), .Q(raddr[36]) );
  DFF_RST raddr_reg_8__4_ ( .D(n430), .CP(clk), .CDN(n34), .Q(raddr[37]) );
  DFF_RST raddr_reg_8__5_ ( .D(n429), .CP(clk), .CDN(n34), .Q(raddr[38]) );
  DFF_RST raddr_reg_8__6_ ( .D(n428), .CP(clk), .CDN(n34), .Q(raddr[39]) );
  DFF_RST raddr_reg_8__7_ ( .D(n427), .CP(clk), .CDN(n35), .Q(raddr[40]) );
  DFF_RST raddr_reg_8__10_ ( .D(n424), .CP(clk), .CDN(n35), .Q(raddr[43])
         );
  DFF_RST raddr_reg_9__0_ ( .D(n423), .CP(clk), .CDN(n35), .Q(raddr[22]) );
  DFF_RST raddr_reg_9__1_ ( .D(n422), .CP(clk), .CDN(n35), .Q(raddr[23]) );
  DFF_RST raddr_reg_9__2_ ( .D(n421), .CP(clk), .CDN(n35), .Q(raddr[24]) );
  DFF_RST raddr_reg_9__3_ ( .D(n420), .CP(clk), .CDN(n35), .Q(raddr[25]) );
  DFF_RST raddr_reg_9__4_ ( .D(n419), .CP(clk), .CDN(n35), .Q(raddr[26]) );
  DFF_RST raddr_reg_9__5_ ( .D(n418), .CP(clk), .CDN(n35), .Q(raddr[27]) );
  DFF_RST raddr_reg_9__6_ ( .D(n417), .CP(clk), .CDN(n35), .Q(raddr[28]) );
  DFF_RST raddr_reg_9__7_ ( .D(n416), .CP(clk), .CDN(n35), .Q(raddr[29]) );
  DFF_RST raddr_reg_9__8_ ( .D(n415), .CP(clk), .CDN(n35), .Q(raddr[30]) );
  DFF_RST raddr_reg_9__9_ ( .D(n414), .CP(clk), .CDN(n35), .Q(raddr[31]) );
  DFF_RST raddr_reg_10__0_ ( .D(n412), .CP(clk), .CDN(n35), .Q(raddr[11])
         );
  DFF_RST raddr_reg_10__1_ ( .D(n411), .CP(clk), .CDN(n36), .Q(raddr[12])
         );
  DFF_RST raddr_reg_10__2_ ( .D(n410), .CP(clk), .CDN(n36), .Q(raddr[13])
         );
  DFF_RST raddr_reg_10__3_ ( .D(n409), .CP(clk), .CDN(n36), .Q(raddr[14])
         );
  DFF_RST raddr_reg_10__4_ ( .D(n408), .CP(clk), .CDN(n36), .Q(raddr[15])
         );
  DFF_RST raddr_reg_10__5_ ( .D(n407), .CP(clk), .CDN(n36), .Q(raddr[16])
         );
  DFF_RST raddr_reg_10__6_ ( .D(n406), .CP(clk), .CDN(n36), .Q(raddr[17])
         );
  DFF_RST raddr_reg_10__7_ ( .D(n405), .CP(clk), .CDN(n36), .Q(raddr[18])
         );
  DFF_RST raddr_reg_10__9_ ( .D(n403), .CP(clk), .CDN(n36), .Q(raddr[20])
         );
  DFF_RST raddr_reg_11__0_ ( .D(n401), .CP(clk), .CDN(n36), .Q(raddr[0]) );
  DFF_RST raddr_reg_11__1_ ( .D(n400), .CP(clk), .CDN(n36), .Q(raddr[1]) );
  DFF_RST raddr_reg_11__2_ ( .D(n399), .CP(clk), .CDN(n36), .Q(raddr[2]) );
  DFF_RST raddr_reg_11__3_ ( .D(n398), .CP(clk), .CDN(n36), .Q(raddr[3]) );
  DFF_RST raddr_reg_11__4_ ( .D(n397), .CP(clk), .CDN(n36), .Q(raddr[4]) );
  DFF_RST raddr_reg_11__5_ ( .D(n396), .CP(clk), .CDN(n37), .Q(raddr[5]) );
  DFF_RST raddr_reg_11__6_ ( .D(n395), .CP(clk), .CDN(n37), .Q(raddr[6]) );
  DFF_RST raddr_reg_11__7_ ( .D(n394), .CP(clk), .CDN(n37), .Q(raddr[7]) );
  DFF_RST raddr_reg_11__8_ ( .D(n393), .CP(clk), .CDN(n37), .Q(raddr[8]) );
  ram2p_2kx8 ram_block ( .wclk(clk), .we(n20), .re(ram_re), .rclk(clk), .din(
        din), .waddr(addra), .raddr(addrb), .dout(dout) );
  fifo_shift_ram_DW01_inc_0 add_203 ( .A(raddr[10:0]), .SUM({N779, N778, N777, 
        N776, N775, N774, N773, N772, N771, N770, N769}) );
  fifo_shift_ram_DW01_inc_1 add_198 ( .A(raddr[21:11]), .SUM({N756, N755, N754, 
        N753, N752, N751, N750, N749, N748, N747, N746}) );
  fifo_shift_ram_DW01_inc_2 add_193 ( .A(raddr[32:22]), .SUM({N733, N732, N731, 
        N730, N729, N728, N727, N726, N725, N724, N723}) );
  fifo_shift_ram_DW01_inc_3 add_188 ( .A(raddr[43:33]), .SUM({N710, N709, N708, 
        N707, N706, N705, N704, N703, N702, N701, N700}) );
  fifo_shift_ram_DW01_inc_4 add_183 ( .A(raddr[54:44]), .SUM({N687, N686, N685, 
        N684, N683, N682, N681, N680, N679, N678, N677}) );
  fifo_shift_ram_DW01_inc_5 add_178 ( .A(raddr[65:55]), .SUM({N664, N663, N662, 
        N661, N660, N659, N658, N657, N656, N655, N654}) );
  fifo_shift_ram_DW01_inc_6 add_173 ( .A(raddr[76:66]), .SUM({N641, N640, N639, 
        N638, N637, N636, N635, N634, N633, N632, N631}) );
  fifo_shift_ram_DW01_inc_7 add_168 ( .A(raddr[87:77]), .SUM({N618, N617, N616, 
        N615, N614, N613, N612, N611, N610, N609, N608}) );
  fifo_shift_ram_DW01_inc_8 add_163 ( .A(raddr[98:88]), .SUM({N595, N594, N593, 
        N592, N591, N590, N589, N588, N587, N586, N585}) );
  fifo_shift_ram_DW01_inc_9 add_158 ( .A(raddr[109:99]), .SUM({N572, N571, 
        N570, N569, N568, N567, N566, N565, N564, N563, N562}) );
  fifo_shift_ram_DW01_inc_10 add_153 ( .A(raddr[120:110]), .SUM({N549, N548, 
        N547, N546, N545, N544, N543, N542, N541, N540, N539}) );
  fifo_shift_ram_DW01_inc_11 add_123 ( .A(waddr[10:0]), .SUM({N359, N358, N357, 
        N356, N355, N354, N353, N352, N351, N350, N349}) );
  fifo_shift_ram_DW01_inc_12 add_118 ( .A(waddr[21:11]), .SUM({N336, N335, 
        N334, N333, N332, N331, N330, N329, N328, N327, N326}) );
  fifo_shift_ram_DW01_inc_13 add_113 ( .A(waddr[32:22]), .SUM({N313, N312, 
        N311, N310, N309, N308, N307, N306, N305, N304, N303}) );
  fifo_shift_ram_DW01_inc_14 add_108 ( .A(waddr[43:33]), .SUM({N290, N289, 
        N288, N287, N286, N285, N284, N283, N282, N281, N280}) );
  fifo_shift_ram_DW01_inc_15 add_103 ( .A(waddr[54:44]), .SUM({N267, N266, 
        N265, N264, N263, N262, N261, N260, N259, N258, N257}) );
  fifo_shift_ram_DW01_inc_16 add_98 ( .A(waddr[65:55]), .SUM({N244, N243, N242, 
        N241, N240, N239, N238, N237, N236, N235, N234}) );
  fifo_shift_ram_DW01_inc_17 add_93 ( .A(waddr[76:66]), .SUM({N221, N220, N219, 
        N218, N217, N216, N215, N214, N213, N212, N211}) );
  fifo_shift_ram_DW01_inc_18 add_88 ( .A(waddr[87:77]), .SUM({N198, N197, N196, 
        N195, N194, N193, N192, N191, N190, N189, N188}) );
  fifo_shift_ram_DW01_inc_19 add_83 ( .A(waddr[98:88]), .SUM({N175, N174, N173, 
        N172, N171, N170, N169, N168, N167, N166, N165}) );
  fifo_shift_ram_DW01_inc_20 add_78 ( .A(waddr[109:99]), .SUM({N152, N151, 
        N150, N149, N148, N147, N146, N145, N144, N143, N142}) );
  fifo_shift_ram_DW01_inc_21 add_73 ( .A(waddr[120:110]), .SUM({N129, N128, 
        N127, N126, N125, N124, N123, N122, N121, N120, N119}) );
  DFF_SET raddr_reg_9__10_ ( .D(n413), .CP(clk), .SDN(n37), .Q(raddr[32])
         );
  DFF_SET raddr_reg_10__10_ ( .D(n402), .CP(clk), .SDN(n37), .Q(raddr[21])
         );
  DFF_SET raddr_reg_11__10_ ( .D(n391), .CP(clk), .SDN(n37), .Q(raddr[10])
         );
  DFF_SET waddr_reg_9__10_ ( .D(n534), .CP(clk), .SDN(n38), .Q(waddr[32])
         );
  DFF_SET waddr_reg_10__10_ ( .D(n523), .CP(clk), .SDN(n38), .Q(waddr[21])
         );
  DFF_SET waddr_reg_3__7_ ( .D(n603), .CP(clk), .SDN(n39), .Q(waddr[95]) );
  DFF_SET waddr_reg_6__9_ ( .D(n568), .CP(clk), .SDN(n38), .Q(waddr[64]) );
  DFF_SET raddr_reg_3__7_ ( .D(n482), .CP(clk), .SDN(n38), .Q(raddr[95]) );
  DFF_SET raddr_reg_6__9_ ( .D(n447), .CP(clk), .SDN(n37), .Q(raddr[64]) );
  DFF_SET waddr_reg_2__6_ ( .D(n615), .CP(clk), .SDN(n39), .Q(waddr[105])
         );
  DFF_SET raddr_reg_2__6_ ( .D(n494), .CP(clk), .SDN(n38), .Q(raddr[105])
         );
  DFF_SET waddr_reg_5__8_ ( .D(n580), .CP(clk), .SDN(n39), .Q(waddr[74]) );
  DFF_SET waddr_reg_8__9_ ( .D(n546), .CP(clk), .SDN(n38), .Q(waddr[42]) );
  DFF_SET waddr_reg_11__9_ ( .D(n513), .CP(clk), .SDN(n38), .Q(waddr[9]) );
  DFF_SET raddr_reg_5__8_ ( .D(n459), .CP(clk), .SDN(n38), .Q(raddr[74]) );
  DFF_SET raddr_reg_8__9_ ( .D(n425), .CP(clk), .SDN(n37), .Q(raddr[42]) );
  DFF_SET raddr_reg_11__9_ ( .D(n392), .CP(clk), .SDN(n37), .Q(raddr[9]) );
  DFF_SET waddr_reg_11__10_ ( .D(n512), .CP(clk), .SDN(n38), .Q(waddr[10])
         );
  DFF_SET waddr_reg_5__7_ ( .D(n581), .CP(clk), .SDN(n39), .Q(waddr[73]) );
  DFF_SET waddr_reg_8__8_ ( .D(n547), .CP(clk), .SDN(n38), .Q(waddr[41]) );
  DFF_SET raddr_reg_5__7_ ( .D(n460), .CP(clk), .SDN(n38), .Q(raddr[73]) );
  DFF_SET raddr_reg_8__8_ ( .D(n426), .CP(clk), .SDN(n37), .Q(raddr[41]) );
  DFF_SET waddr_reg_4__8_ ( .D(n591), .CP(clk), .SDN(n39), .Q(waddr[85]) );
  DFF_SET waddr_reg_7__9_ ( .D(n557), .CP(clk), .SDN(n38), .Q(waddr[53]) );
  DFF_SET waddr_reg_10__8_ ( .D(n525), .CP(clk), .SDN(n38), .Q(waddr[19])
         );
  DFF_SET raddr_reg_4__8_ ( .D(n470), .CP(clk), .SDN(n38), .Q(raddr[85]) );
  DFF_SET raddr_reg_7__9_ ( .D(n436), .CP(clk), .SDN(n37), .Q(raddr[53]) );
  DFF_SET raddr_reg_10__8_ ( .D(n404), .CP(clk), .SDN(n37), .Q(raddr[19])
         );
  DFF_SET waddr_reg_7__7_ ( .D(n559), .CP(clk), .SDN(n38), .Q(waddr[51]) );
  DFF_SET raddr_reg_7__7_ ( .D(n438), .CP(clk), .SDN(n37), .Q(raddr[51]) );
  I_NAND4 U3 ( .A1(n2), .B1(n297), .B2(n298), .B3(n299), .ZN(addrb[9]) );
  AND4 U4 ( .A1(n387), .A2(n388), .A3(n389), .A4(n390), .Z(n1) );
  INV U5 ( .I(n1), .ZN(n20) );
  AO22 U6 ( .A1(raddr[108]), .A2(n3), .B1(raddr[119]), .B2(n5), .Z(n2) );
  NAND4 U7 ( .A1(n372), .A2(n373), .A3(n374), .A4(n375), .ZN(addra[1]) );
  NAND4 U8 ( .A1(n380), .A2(n381), .A3(n382), .A4(n383), .ZN(addra[0]) );
  NAND4 U9 ( .A1(n368), .A2(n369), .A3(n370), .A4(n371), .ZN(addra[2]) );
  NAND4 U10 ( .A1(n352), .A2(n353), .A3(n354), .A4(n355), .ZN(addra[6]) );
  NAND4 U11 ( .A1(n364), .A2(n365), .A3(n366), .A4(n367), .ZN(addra[3]) );
  NAND4 U12 ( .A1(n348), .A2(n349), .A3(n350), .A4(n351), .ZN(addra[7]) );
  NAND4 U13 ( .A1(n360), .A2(n361), .A3(n362), .A4(n363), .ZN(addra[4]) );
  NAND4 U14 ( .A1(n344), .A2(n345), .A3(n346), .A4(n347), .ZN(addra[8]) );
  NAND4 U15 ( .A1(n356), .A2(n357), .A3(n358), .A4(n359), .ZN(addra[5]) );
  BUF U16 ( .I(n41), .Z(n36) );
  BUF U17 ( .I(n41), .Z(n35) );
  BUF U18 ( .I(n41), .Z(n34) );
  BUF U19 ( .I(n42), .Z(n33) );
  BUF U20 ( .I(n42), .Z(n32) );
  BUF U21 ( .I(n42), .Z(n31) );
  BUF U22 ( .I(n43), .Z(n30) );
  BUF U23 ( .I(n43), .Z(n29) );
  BUF U24 ( .I(n43), .Z(n28) );
  BUF U25 ( .I(n44), .Z(n27) );
  BUF U26 ( .I(n44), .Z(n26) );
  BUF U27 ( .I(n44), .Z(n25) );
  BUF U28 ( .I(n45), .Z(n24) );
  BUF U29 ( .I(n45), .Z(n23) );
  BUF U30 ( .I(n45), .Z(n22) );
  AND2 U31 ( .A1(n386), .A2(n384), .Z(n289) );
  AND2 U32 ( .A1(n386), .A2(n384), .Z(n3) );
  AND2 U33 ( .A1(n386), .A2(n384), .Z(n4) );
  INV U34 ( .I(n143), .ZN(n676) );
  INV U35 ( .I(n151), .ZN(n675) );
  INV U36 ( .I(n159), .ZN(n674) );
  INV U37 ( .I(n180), .ZN(n671) );
  INV U38 ( .I(n173), .ZN(n672) );
  INV U39 ( .I(n202), .ZN(n668) );
  INV U40 ( .I(n188), .ZN(n670) );
  INV U41 ( .I(n195), .ZN(n669) );
  INV U42 ( .I(n135), .ZN(n677) );
  INV U43 ( .I(n165), .ZN(n673) );
  BUF U44 ( .I(n46), .Z(n21) );
  BUF U45 ( .I(n47), .Z(n46) );
  BUF U46 ( .I(n40), .Z(n38) );
  BUF U47 ( .I(n40), .Z(n37) );
  BUF U48 ( .I(n48), .Z(n41) );
  BUF U49 ( .I(n48), .Z(n42) );
  BUF U50 ( .I(n48), .Z(n43) );
  BUF U51 ( .I(n47), .Z(n44) );
  BUF U52 ( .I(n47), .Z(n45) );
  BUF U53 ( .I(n40), .Z(n39) );
  NOR2 U54 ( .A1(sel[2]), .A2(sel[1]), .ZN(n384) );
  I_NOR2 U55 ( .A1(sel[3]), .B1(n384), .ZN(n222) );
  AND3 U56 ( .A1(n385), .A2(sel[2]), .A3(sel[1]), .Z(n253) );
  AND3 U57 ( .A1(n386), .A2(sel[1]), .A3(sel[2]), .Z(n245) );
  NOR2 U58 ( .A1(n679), .A2(sel[3]), .ZN(n386) );
  BUF U59 ( .I(n275), .Z(n9) );
  I_NOR3 U60 ( .A1(n386), .B1(sel[2]), .B2(n678), .ZN(n275) );
  BUF U61 ( .I(n282), .Z(n7) );
  I_NOR3 U62 ( .A1(n385), .B1(n678), .B2(sel[2]), .ZN(n282) );
  I_NOR2 U63 ( .A1(sel[3]), .B1(n384), .ZN(n12) );
  AND3 U64 ( .A1(n385), .A2(sel[2]), .A3(sel[1]), .Z(n10) );
  AND3 U65 ( .A1(n386), .A2(n678), .A3(sel[2]), .Z(n260) );
  AND3 U66 ( .A1(sel[3]), .A2(n679), .A3(n384), .Z(n237) );
  AND3 U67 ( .A1(sel[3]), .A2(n679), .A3(n384), .Z(n11) );
  AND3 U68 ( .A1(n385), .A2(sel[2]), .A3(n678), .Z(n268) );
  AND3 U69 ( .A1(n385), .A2(sel[2]), .A3(n678), .Z(n8) );
  AND2 U70 ( .A1(n385), .A2(n384), .Z(n6) );
  AND2 U71 ( .A1(n385), .A2(n384), .Z(n5) );
  AND2 U72 ( .A1(n385), .A2(n384), .Z(n295) );
  NAND2 U73 ( .A1(n13), .A2(n20), .ZN(n143) );
  NAND2 U74 ( .A1(n4), .A2(n20), .ZN(n202) );
  NAND2 U75 ( .A1(n245), .A2(n20), .ZN(n159) );
  NAND2 U76 ( .A1(n9), .A2(n20), .ZN(n188) );
  NAND2 U77 ( .A1(n7), .A2(n20), .ZN(n195) );
  NAND2 U78 ( .A1(n8), .A2(n20), .ZN(n180) );
  NAND2 U79 ( .A1(n260), .A2(n20), .ZN(n173) );
  NAND2 U80 ( .A1(n11), .A2(n20), .ZN(n151) );
  NAND2 U81 ( .A1(n222), .A2(n20), .ZN(n18) );
  NAND2 U82 ( .A1(n12), .A2(n20), .ZN(n135) );
  NAND2 U83 ( .A1(n12), .A2(n20), .ZN(n19) );
  NAND2 U84 ( .A1(n253), .A2(n20), .ZN(n16) );
  NAND2 U85 ( .A1(n10), .A2(n20), .ZN(n165) );
  NAND2 U86 ( .A1(n10), .A2(n20), .ZN(n17) );
  AND2 U87 ( .A1(n6), .A2(n20), .Z(n15) );
  AND2 U88 ( .A1(n295), .A2(n20), .Z(n209) );
  AND2 U89 ( .A1(n6), .A2(n20), .Z(n14) );
  BUF U90 ( .I(reset_n), .Z(n48) );
  BUF U91 ( .I(reset_n), .Z(n47) );
  BUF U92 ( .I(n49), .Z(n40) );
  BUF U93 ( .I(reset_n), .Z(n49) );
  AND3 U94 ( .A1(n384), .A2(sel[3]), .A3(sel[0]), .Z(n230) );
  AND3 U95 ( .A1(n384), .A2(sel[3]), .A3(sel[0]), .Z(n13) );
  NOR2 U96 ( .A1(sel[3]), .A2(sel[0]), .ZN(n385) );
  NOR3 U97 ( .A1(push[1]), .A2(push[3]), .A3(push[2]), .ZN(n388) );
  NOR3 U98 ( .A1(push[7]), .A2(push[9]), .A3(push[8]), .ZN(n390) );
  NOR3 U99 ( .A1(push[4]), .A2(push[6]), .A3(push[5]), .ZN(n389) );
  NOR2 U100 ( .A1(push[10]), .A2(push[0]), .ZN(n387) );
  NOR2 U101 ( .A1(n202), .A2(n205), .ZN(n203) );
  NOR2 U102 ( .A1(n202), .A2(n285), .ZN(n283) );
  NOR2 U103 ( .A1(n143), .A2(n144), .ZN(n145) );
  NOR2 U104 ( .A1(n143), .A2(n224), .ZN(n225) );
  NOR2 U105 ( .A1(n188), .A2(n191), .ZN(n189) );
  NOR2 U106 ( .A1(n195), .A2(n198), .ZN(n196) );
  NOR2 U107 ( .A1(n188), .A2(n271), .ZN(n269) );
  NOR2 U108 ( .A1(n195), .A2(n278), .ZN(n276) );
  NOR2 U109 ( .A1(n173), .A2(n176), .ZN(n174) );
  NOR2 U110 ( .A1(n173), .A2(n256), .ZN(n254) );
  NOR2 U111 ( .A1(n159), .A2(n160), .ZN(n157) );
  NOR2 U112 ( .A1(n159), .A2(n240), .ZN(n238) );
  NOR2 U113 ( .A1(n18), .A2(n216), .ZN(n218) );
  NOR2 U114 ( .A1(n19), .A2(n136), .ZN(n138) );
  NOR2 U115 ( .A1(n16), .A2(n248), .ZN(n246) );
  NOR2 U116 ( .A1(n17), .A2(n168), .ZN(n166) );
  NOR2 U117 ( .A1(n180), .A2(n183), .ZN(n181) );
  NOR2 U118 ( .A1(n180), .A2(n263), .ZN(n261) );
  AND2 U119 ( .A1(n152), .A2(n675), .Z(n153) );
  AND2 U120 ( .A1(n232), .A2(n675), .Z(n233) );
  MOAI22 U121 ( .A1(n209), .A2(n119), .B1(N548), .B2(n210), .ZN(n502) );
  MOAI22 U122 ( .A1(n15), .A2(n118), .B1(N547), .B2(n210), .ZN(n503) );
  MOAI22 U123 ( .A1(n209), .A2(n58), .B1(N127), .B2(n290), .ZN(n624) );
  MOAI22 U124 ( .A1(n15), .A2(n57), .B1(N126), .B2(n290), .ZN(n625) );
  MOAI22 U125 ( .A1(n14), .A2(n117), .B1(N546), .B2(n210), .ZN(n504) );
  MOAI22 U126 ( .A1(n14), .A2(n59), .B1(N128), .B2(n290), .ZN(n623) );
  MOAI22 U127 ( .A1(n675), .A2(n657), .B1(N732), .B2(n153), .ZN(n414) );
  MOAI22 U128 ( .A1(n675), .A2(n656), .B1(N731), .B2(n153), .ZN(n415) );
  MOAI22 U129 ( .A1(n675), .A2(n655), .B1(N729), .B2(n153), .ZN(n417) );
  MOAI22 U130 ( .A1(n675), .A2(n654), .B1(N726), .B2(n153), .ZN(n420) );
  MOAI22 U131 ( .A1(n675), .A2(n99), .B1(N312), .B2(n233), .ZN(n535) );
  MOAI22 U132 ( .A1(n675), .A2(n98), .B1(N311), .B2(n233), .ZN(n536) );
  MOAI22 U133 ( .A1(n675), .A2(n97), .B1(N309), .B2(n233), .ZN(n538) );
  MOAI22 U134 ( .A1(n675), .A2(n96), .B1(N306), .B2(n233), .ZN(n541) );
  MOAI22 U135 ( .A1(n676), .A2(n662), .B1(N751), .B2(n145), .ZN(n407) );
  MOAI22 U136 ( .A1(n676), .A2(n661), .B1(N749), .B2(n145), .ZN(n409) );
  MOAI22 U137 ( .A1(n676), .A2(n660), .B1(N748), .B2(n145), .ZN(n410) );
  MOAI22 U138 ( .A1(n676), .A2(n659), .B1(N747), .B2(n145), .ZN(n411) );
  MOAI22 U139 ( .A1(n676), .A2(n104), .B1(N331), .B2(n225), .ZN(n528) );
  MOAI22 U140 ( .A1(n676), .A2(n103), .B1(N329), .B2(n225), .ZN(n530) );
  MOAI22 U141 ( .A1(n676), .A2(n102), .B1(N328), .B2(n225), .ZN(n531) );
  MOAI22 U142 ( .A1(n676), .A2(n101), .B1(N327), .B2(n225), .ZN(n532) );
  MOAI22 U143 ( .A1(n674), .A2(n652), .B1(N707), .B2(n157), .ZN(n427) );
  MOAI22 U144 ( .A1(n674), .A2(n651), .B1(N703), .B2(n157), .ZN(n431) );
  MOAI22 U145 ( .A1(n674), .A2(n650), .B1(N702), .B2(n157), .ZN(n432) );
  MOAI22 U146 ( .A1(n674), .A2(n649), .B1(N701), .B2(n157), .ZN(n433) );
  MOAI22 U147 ( .A1(n672), .A2(n644), .B1(N662), .B2(n174), .ZN(n448) );
  MOAI22 U148 ( .A1(n672), .A2(n643), .B1(N661), .B2(n174), .ZN(n449) );
  MOAI22 U149 ( .A1(n672), .A2(n642), .B1(N659), .B2(n174), .ZN(n451) );
  MOAI22 U150 ( .A1(n672), .A2(n641), .B1(N658), .B2(n174), .ZN(n452) );
  MOAI22 U151 ( .A1(n672), .A2(n640), .B1(N656), .B2(n174), .ZN(n454) );
  MOAI22 U152 ( .A1(n674), .A2(n94), .B1(N287), .B2(n238), .ZN(n548) );
  MOAI22 U153 ( .A1(n674), .A2(n93), .B1(N283), .B2(n238), .ZN(n552) );
  MOAI22 U154 ( .A1(n674), .A2(n92), .B1(N282), .B2(n238), .ZN(n553) );
  MOAI22 U155 ( .A1(n674), .A2(n91), .B1(N281), .B2(n238), .ZN(n554) );
  MOAI22 U156 ( .A1(n672), .A2(n86), .B1(N242), .B2(n254), .ZN(n569) );
  MOAI22 U157 ( .A1(n672), .A2(n85), .B1(N241), .B2(n254), .ZN(n570) );
  MOAI22 U158 ( .A1(n672), .A2(n84), .B1(N239), .B2(n254), .ZN(n572) );
  MOAI22 U159 ( .A1(n672), .A2(n83), .B1(N238), .B2(n254), .ZN(n573) );
  MOAI22 U160 ( .A1(n672), .A2(n82), .B1(N236), .B2(n254), .ZN(n575) );
  MOAI22 U161 ( .A1(n671), .A2(n638), .B1(N640), .B2(n181), .ZN(n458) );
  MOAI22 U162 ( .A1(n671), .A2(n637), .B1(N637), .B2(n181), .ZN(n461) );
  MOAI22 U163 ( .A1(n671), .A2(n636), .B1(N636), .B2(n181), .ZN(n462) );
  MOAI22 U164 ( .A1(n671), .A2(n635), .B1(N635), .B2(n181), .ZN(n463) );
  MOAI22 U165 ( .A1(n671), .A2(n634), .B1(N634), .B2(n181), .ZN(n464) );
  MOAI22 U166 ( .A1(n671), .A2(n633), .B1(N633), .B2(n181), .ZN(n465) );
  MOAI22 U167 ( .A1(n671), .A2(n80), .B1(N220), .B2(n261), .ZN(n579) );
  MOAI22 U168 ( .A1(n671), .A2(n79), .B1(N217), .B2(n261), .ZN(n582) );
  MOAI22 U169 ( .A1(n671), .A2(n78), .B1(N216), .B2(n261), .ZN(n583) );
  MOAI22 U170 ( .A1(n671), .A2(n77), .B1(N215), .B2(n261), .ZN(n584) );
  MOAI22 U171 ( .A1(n671), .A2(n76), .B1(N214), .B2(n261), .ZN(n585) );
  MOAI22 U172 ( .A1(n671), .A2(n75), .B1(N213), .B2(n261), .ZN(n586) );
  MOAI22 U173 ( .A1(n670), .A2(n296), .B1(N617), .B2(n189), .ZN(n469) );
  MOAI22 U174 ( .A1(n670), .A2(n133), .B1(N615), .B2(n189), .ZN(n471) );
  MOAI22 U175 ( .A1(n670), .A2(n132), .B1(N613), .B2(n189), .ZN(n473) );
  MOAI22 U176 ( .A1(n670), .A2(n131), .B1(N609), .B2(n189), .ZN(n477) );
  MOAI22 U177 ( .A1(n669), .A2(n129), .B1(N594), .B2(n196), .ZN(n480) );
  MOAI22 U178 ( .A1(n669), .A2(n128), .B1(N593), .B2(n196), .ZN(n481) );
  MOAI22 U179 ( .A1(n669), .A2(n127), .B1(N591), .B2(n196), .ZN(n483) );
  MOAI22 U180 ( .A1(n669), .A2(n126), .B1(N589), .B2(n196), .ZN(n485) );
  MOAI22 U181 ( .A1(n669), .A2(n125), .B1(N586), .B2(n196), .ZN(n488) );
  MOAI22 U182 ( .A1(n670), .A2(n74), .B1(N197), .B2(n269), .ZN(n590) );
  MOAI22 U183 ( .A1(n670), .A2(n73), .B1(N195), .B2(n269), .ZN(n592) );
  MOAI22 U184 ( .A1(n670), .A2(n72), .B1(N193), .B2(n269), .ZN(n594) );
  MOAI22 U185 ( .A1(n670), .A2(n71), .B1(N189), .B2(n269), .ZN(n598) );
  MOAI22 U186 ( .A1(n669), .A2(n69), .B1(N174), .B2(n276), .ZN(n601) );
  MOAI22 U187 ( .A1(n669), .A2(n68), .B1(N173), .B2(n276), .ZN(n602) );
  MOAI22 U188 ( .A1(n669), .A2(n67), .B1(N171), .B2(n276), .ZN(n604) );
  MOAI22 U189 ( .A1(n669), .A2(n66), .B1(N169), .B2(n276), .ZN(n606) );
  MOAI22 U190 ( .A1(n669), .A2(n65), .B1(N166), .B2(n276), .ZN(n609) );
  MOAI22 U191 ( .A1(n677), .A2(n667), .B1(N774), .B2(n138), .ZN(n396) );
  MOAI22 U192 ( .A1(n677), .A2(n666), .B1(N773), .B2(n138), .ZN(n397) );
  MOAI22 U193 ( .A1(n677), .A2(n665), .B1(N772), .B2(n138), .ZN(n398) );
  MOAI22 U194 ( .A1(n673), .A2(n648), .B1(N683), .B2(n166), .ZN(n439) );
  MOAI22 U195 ( .A1(n673), .A2(n647), .B1(N682), .B2(n166), .ZN(n440) );
  MOAI22 U196 ( .A1(n673), .A2(n646), .B1(N681), .B2(n166), .ZN(n441) );
  MOAI22 U197 ( .A1(n668), .A2(n124), .B1(N571), .B2(n203), .ZN(n491) );
  MOAI22 U198 ( .A1(n668), .A2(n123), .B1(N570), .B2(n203), .ZN(n492) );
  MOAI22 U199 ( .A1(n668), .A2(n122), .B1(N569), .B2(n203), .ZN(n493) );
  MOAI22 U200 ( .A1(n677), .A2(n109), .B1(N354), .B2(n218), .ZN(n517) );
  MOAI22 U201 ( .A1(n677), .A2(n108), .B1(N353), .B2(n218), .ZN(n518) );
  MOAI22 U202 ( .A1(n677), .A2(n107), .B1(N352), .B2(n218), .ZN(n519) );
  MOAI22 U203 ( .A1(n673), .A2(n90), .B1(N263), .B2(n246), .ZN(n560) );
  MOAI22 U204 ( .A1(n673), .A2(n89), .B1(N262), .B2(n246), .ZN(n561) );
  MOAI22 U205 ( .A1(n673), .A2(n88), .B1(N261), .B2(n246), .ZN(n562) );
  MOAI22 U206 ( .A1(n668), .A2(n64), .B1(N151), .B2(n283), .ZN(n612) );
  MOAI22 U207 ( .A1(n668), .A2(n63), .B1(N150), .B2(n283), .ZN(n613) );
  MOAI22 U208 ( .A1(n668), .A2(n62), .B1(N149), .B2(n283), .ZN(n614) );
  NAND3 U209 ( .A1(n118), .A2(n119), .A3(n117), .ZN(n214) );
  NAND3 U210 ( .A1(n58), .A2(n59), .A3(n57), .ZN(n294) );
  NAND4 U211 ( .A1(n336), .A2(n337), .A3(n338), .A4(n339), .ZN(addrb[0]) );
  AOI22 U212 ( .A1(raddr[99]), .A2(n289), .B1(raddr[110]), .B2(n295), 
        .ZN(n336) );
  AOI222 U213 ( .A1(raddr[55]), .A2(n260), .B1(raddr[33]), .B2(n245), 
        .C1(raddr[44]), .C2(n253), .ZN(n338) );
  AOI222 U214 ( .A1(raddr[88]), .A2(n7), .B1(raddr[66]), .B2(n268), .C1(
        raddr[77]), .C2(n9), .ZN(n337) );
  NAND4 U215 ( .A1(n328), .A2(n329), .A3(n330), .A4(n331), .ZN(addrb[1]) );
  AOI22 U216 ( .A1(raddr[100]), .A2(n4), .B1(raddr[111]), .B2(n6), .ZN(
        n328) );
  AOI222 U217 ( .A1(raddr[56]), .A2(n260), .B1(raddr[34]), .B2(n245), 
        .C1(raddr[45]), .C2(n253), .ZN(n330) );
  AOI222 U218 ( .A1(raddr[89]), .A2(n7), .B1(raddr[67]), .B2(n268), .C1(
        raddr[78]), .C2(n9), .ZN(n329) );
  AOI222 U219 ( .A1(raddr[22]), .A2(n237), .B1(raddr[0]), .B2(n222), .C1(
        raddr[11]), .C2(n230), .ZN(n339) );
  AOI222 U220 ( .A1(raddr[23]), .A2(n237), .B1(raddr[1]), .B2(n222), .C1(
        raddr[12]), .C2(n230), .ZN(n331) );
  AOI222 U221 ( .A1(raddr[25]), .A2(n237), .B1(raddr[3]), .B2(n222), .C1(
        raddr[14]), .C2(n230), .ZN(n323) );
  AOI222 U222 ( .A1(raddr[24]), .A2(n11), .B1(raddr[2]), .B2(n12), .C1(
        raddr[13]), .C2(n13), .ZN(n327) );
  AOI222 U223 ( .A1(raddr[91]), .A2(n7), .B1(raddr[69]), .B2(n268), .C1(
        raddr[80]), .C2(n9), .ZN(n321) );
  AOI222 U224 ( .A1(raddr[90]), .A2(n7), .B1(raddr[68]), .B2(n8), .C1(
        raddr[79]), .C2(n9), .ZN(n325) );
  NAND4 U225 ( .A1(n320), .A2(n321), .A3(n322), .A4(n323), .ZN(addrb[3]) );
  AOI22 U226 ( .A1(raddr[102]), .A2(n3), .B1(raddr[113]), .B2(n5), .ZN(
        n320) );
  AOI222 U227 ( .A1(raddr[58]), .A2(n260), .B1(raddr[36]), .B2(n245), 
        .C1(raddr[47]), .C2(n253), .ZN(n322) );
  NAND4 U228 ( .A1(n324), .A2(n325), .A3(n326), .A4(n327), .ZN(addrb[2]) );
  AOI22 U229 ( .A1(raddr[101]), .A2(n289), .B1(raddr[112]), .B2(n295), 
        .ZN(n324) );
  AOI222 U230 ( .A1(raddr[57]), .A2(n260), .B1(raddr[35]), .B2(n245), 
        .C1(raddr[46]), .C2(n10), .ZN(n326) );
  AOI22 U231 ( .A1(waddr[105]), .A2(n4), .B1(waddr[116]), .B2(n6), .ZN(
        n352) );
  AOI222 U232 ( .A1(waddr[61]), .A2(n260), .B1(waddr[39]), .B2(n245), 
        .C1(waddr[50]), .C2(n253), .ZN(n354) );
  AOI222 U233 ( .A1(waddr[94]), .A2(n7), .B1(waddr[72]), .B2(n268), .C1(
        waddr[83]), .C2(n9), .ZN(n353) );
  AOI22 U234 ( .A1(waddr[102]), .A2(n4), .B1(waddr[113]), .B2(n6), .ZN(
        n364) );
  AOI222 U235 ( .A1(waddr[58]), .A2(n260), .B1(waddr[36]), .B2(n245), 
        .C1(waddr[47]), .C2(n10), .ZN(n366) );
  AOI222 U236 ( .A1(waddr[91]), .A2(n7), .B1(waddr[69]), .B2(n8), .C1(
        waddr[80]), .C2(n9), .ZN(n365) );
  AOI22 U237 ( .A1(waddr[99]), .A2(n3), .B1(waddr[110]), .B2(n5), .ZN(
        n380) );
  AOI222 U238 ( .A1(waddr[55]), .A2(n260), .B1(waddr[33]), .B2(n245), 
        .C1(waddr[44]), .C2(n253), .ZN(n382) );
  AOI222 U239 ( .A1(waddr[88]), .A2(n7), .B1(waddr[66]), .B2(n268), .C1(
        waddr[77]), .C2(n9), .ZN(n381) );
  AOI22 U240 ( .A1(waddr[106]), .A2(n289), .B1(waddr[117]), .B2(n295), 
        .ZN(n348) );
  AOI222 U241 ( .A1(waddr[62]), .A2(n260), .B1(waddr[40]), .B2(n245), 
        .C1(waddr[51]), .C2(n10), .ZN(n350) );
  AOI222 U242 ( .A1(waddr[95]), .A2(n7), .B1(waddr[73]), .B2(n8), .C1(
        waddr[84]), .C2(n9), .ZN(n349) );
  AOI22 U243 ( .A1(waddr[103]), .A2(n289), .B1(waddr[114]), .B2(n295), 
        .ZN(n360) );
  AOI222 U244 ( .A1(waddr[59]), .A2(n260), .B1(waddr[37]), .B2(n245), 
        .C1(waddr[48]), .C2(n253), .ZN(n362) );
  AOI222 U245 ( .A1(waddr[92]), .A2(n7), .B1(waddr[70]), .B2(n268), .C1(
        waddr[81]), .C2(n9), .ZN(n361) );
  AOI22 U246 ( .A1(waddr[100]), .A2(n289), .B1(waddr[111]), .B2(n295), 
        .ZN(n372) );
  AOI222 U247 ( .A1(waddr[56]), .A2(n260), .B1(waddr[34]), .B2(n245), 
        .C1(waddr[45]), .C2(n10), .ZN(n374) );
  AOI222 U248 ( .A1(waddr[89]), .A2(n7), .B1(waddr[67]), .B2(n8), .C1(
        waddr[78]), .C2(n9), .ZN(n373) );
  AOI22 U249 ( .A1(waddr[107]), .A2(n3), .B1(waddr[118]), .B2(n5), .ZN(
        n344) );
  AOI222 U250 ( .A1(waddr[63]), .A2(n260), .B1(waddr[41]), .B2(n245), 
        .C1(waddr[52]), .C2(n253), .ZN(n346) );
  AOI222 U251 ( .A1(waddr[96]), .A2(n7), .B1(waddr[74]), .B2(n268), .C1(
        waddr[85]), .C2(n9), .ZN(n345) );
  AOI22 U252 ( .A1(waddr[104]), .A2(n3), .B1(waddr[115]), .B2(n5), .ZN(
        n356) );
  AOI222 U253 ( .A1(waddr[60]), .A2(n260), .B1(waddr[38]), .B2(n245), 
        .C1(waddr[49]), .C2(n10), .ZN(n358) );
  AOI222 U254 ( .A1(waddr[93]), .A2(n7), .B1(waddr[71]), .B2(n8), .C1(
        waddr[82]), .C2(n9), .ZN(n357) );
  AOI22 U255 ( .A1(waddr[101]), .A2(n3), .B1(waddr[112]), .B2(n5), .ZN(
        n368) );
  AOI222 U256 ( .A1(waddr[57]), .A2(n260), .B1(waddr[35]), .B2(n245), 
        .C1(waddr[46]), .C2(n253), .ZN(n370) );
  AOI222 U257 ( .A1(waddr[90]), .A2(n7), .B1(waddr[68]), .B2(n268), .C1(
        waddr[79]), .C2(n9), .ZN(n369) );
  AOI222 U258 ( .A1(raddr[27]), .A2(n237), .B1(raddr[5]), .B2(n222), .C1(
        raddr[16]), .C2(n230), .ZN(n315) );
  AOI222 U259 ( .A1(waddr[30]), .A2(n237), .B1(waddr[8]), .B2(n222), .C1(
        waddr[19]), .C2(n230), .ZN(n347) );
  AOI222 U260 ( .A1(waddr[28]), .A2(n237), .B1(waddr[6]), .B2(n222), .C1(
        waddr[17]), .C2(n230), .ZN(n355) );
  AOI222 U261 ( .A1(waddr[26]), .A2(n237), .B1(waddr[4]), .B2(n222), .C1(
        waddr[15]), .C2(n230), .ZN(n363) );
  AOI222 U262 ( .A1(waddr[24]), .A2(n237), .B1(waddr[2]), .B2(n222), .C1(
        waddr[13]), .C2(n230), .ZN(n371) );
  AOI222 U263 ( .A1(waddr[22]), .A2(n237), .B1(waddr[0]), .B2(n222), .C1(
        waddr[11]), .C2(n230), .ZN(n383) );
  AOI222 U264 ( .A1(raddr[29]), .A2(n237), .B1(raddr[7]), .B2(n222), .C1(
        raddr[18]), .C2(n230), .ZN(n307) );
  AOI222 U265 ( .A1(raddr[26]), .A2(n11), .B1(raddr[4]), .B2(n12), .C1(
        raddr[15]), .C2(n13), .ZN(n319) );
  AOI222 U266 ( .A1(waddr[29]), .A2(n11), .B1(waddr[7]), .B2(n12), .C1(
        waddr[18]), .C2(n13), .ZN(n351) );
  AOI222 U267 ( .A1(waddr[27]), .A2(n11), .B1(waddr[5]), .B2(n12), .C1(
        waddr[16]), .C2(n13), .ZN(n359) );
  AOI222 U268 ( .A1(waddr[25]), .A2(n11), .B1(waddr[3]), .B2(n12), .C1(
        waddr[14]), .C2(n13), .ZN(n367) );
  AOI222 U269 ( .A1(waddr[23]), .A2(n11), .B1(waddr[1]), .B2(n12), .C1(
        waddr[12]), .C2(n13), .ZN(n375) );
  AOI222 U270 ( .A1(raddr[28]), .A2(n11), .B1(raddr[6]), .B2(n12), .C1(
        raddr[17]), .C2(n13), .ZN(n311) );
  AOI222 U271 ( .A1(raddr[62]), .A2(n260), .B1(raddr[40]), .B2(n245), 
        .C1(raddr[51]), .C2(n253), .ZN(n306) );
  AOI222 U272 ( .A1(raddr[93]), .A2(n7), .B1(raddr[71]), .B2(n268), .C1(
        raddr[82]), .C2(n9), .ZN(n313) );
  AOI222 U273 ( .A1(raddr[92]), .A2(n7), .B1(raddr[70]), .B2(n8), .C1(
        raddr[81]), .C2(n9), .ZN(n317) );
  AOI222 U274 ( .A1(raddr[95]), .A2(n7), .B1(raddr[73]), .B2(n268), .C1(
        raddr[84]), .C2(n9), .ZN(n305) );
  AOI222 U275 ( .A1(raddr[94]), .A2(n7), .B1(raddr[72]), .B2(n8), .C1(
        raddr[83]), .C2(n9), .ZN(n309) );
  NAND4 U276 ( .A1(n312), .A2(n313), .A3(n314), .A4(n315), .ZN(addrb[5]) );
  AOI22 U277 ( .A1(raddr[104]), .A2(n289), .B1(raddr[115]), .B2(n295), 
        .ZN(n312) );
  AOI222 U278 ( .A1(raddr[60]), .A2(n260), .B1(raddr[38]), .B2(n245), 
        .C1(raddr[49]), .C2(n253), .ZN(n314) );
  NAND4 U279 ( .A1(n316), .A2(n317), .A3(n318), .A4(n319), .ZN(addrb[4]) );
  AOI22 U280 ( .A1(raddr[103]), .A2(n4), .B1(raddr[114]), .B2(n6), .ZN(
        n316) );
  AOI222 U281 ( .A1(raddr[59]), .A2(n260), .B1(raddr[37]), .B2(n245), 
        .C1(raddr[48]), .C2(n10), .ZN(n318) );
  NAND4 U282 ( .A1(n304), .A2(n305), .A3(n306), .A4(n307), .ZN(addrb[7]) );
  AOI22 U283 ( .A1(raddr[106]), .A2(n4), .B1(raddr[117]), .B2(n6), .ZN(
        n304) );
  NAND4 U284 ( .A1(n308), .A2(n309), .A3(n310), .A4(n311), .ZN(addrb[6]) );
  AOI22 U285 ( .A1(raddr[105]), .A2(n3), .B1(raddr[116]), .B2(n5), .ZN(
        n308) );
  AOI222 U286 ( .A1(raddr[64]), .A2(n260), .B1(raddr[42]), .B2(n245), 
        .C1(raddr[53]), .C2(n253), .ZN(n298) );
  AOI222 U287 ( .A1(raddr[97]), .A2(n7), .B1(raddr[75]), .B2(n268), .C1(
        raddr[86]), .C2(n9), .ZN(n297) );
  NAND4 U288 ( .A1(n332), .A2(n333), .A3(n334), .A4(n335), .ZN(addrb[10])
         );
  AOI22 U289 ( .A1(raddr[109]), .A2(n3), .B1(raddr[120]), .B2(n5), .ZN(
        n332) );
  AOI222 U290 ( .A1(raddr[65]), .A2(n260), .B1(raddr[43]), .B2(n245), 
        .C1(raddr[54]), .C2(n10), .ZN(n334) );
  AOI222 U291 ( .A1(raddr[98]), .A2(n7), .B1(raddr[76]), .B2(n8), .C1(
        raddr[87]), .C2(n9), .ZN(n333) );
  NAND4 U292 ( .A1(n340), .A2(n341), .A3(n342), .A4(n343), .ZN(addra[9]) );
  AOI22 U293 ( .A1(waddr[108]), .A2(n4), .B1(waddr[119]), .B2(n6), .ZN(
        n340) );
  AOI222 U294 ( .A1(waddr[64]), .A2(n260), .B1(waddr[42]), .B2(n245), 
        .C1(waddr[53]), .C2(n10), .ZN(n342) );
  AOI222 U295 ( .A1(waddr[97]), .A2(n7), .B1(waddr[75]), .B2(n8), .C1(
        waddr[86]), .C2(n9), .ZN(n341) );
  NAND4 U296 ( .A1(n376), .A2(n377), .A3(n378), .A4(n379), .ZN(addra[10])
         );
  AOI22 U297 ( .A1(waddr[109]), .A2(n289), .B1(waddr[120]), .B2(n6), .ZN(
        n376) );
  AOI222 U298 ( .A1(waddr[65]), .A2(n260), .B1(waddr[43]), .B2(n245), 
        .C1(waddr[54]), .C2(n253), .ZN(n378) );
  AOI222 U299 ( .A1(waddr[98]), .A2(n7), .B1(waddr[76]), .B2(n268), .C1(
        waddr[87]), .C2(n9), .ZN(n377) );
  AOI222 U300 ( .A1(waddr[32]), .A2(n237), .B1(waddr[10]), .B2(n222), 
        .C1(waddr[21]), .C2(n230), .ZN(n379) );
  AOI222 U301 ( .A1(raddr[31]), .A2(n237), .B1(raddr[9]), .B2(n222), .C1(
        raddr[20]), .C2(n230), .ZN(n299) );
  AOI222 U302 ( .A1(waddr[31]), .A2(n11), .B1(waddr[9]), .B2(n12), .C1(
        waddr[20]), .C2(n13), .ZN(n343) );
  AOI222 U303 ( .A1(raddr[30]), .A2(n11), .B1(raddr[8]), .B2(n12), .C1(
        raddr[19]), .C2(n13), .ZN(n303) );
  AOI222 U304 ( .A1(raddr[32]), .A2(n11), .B1(raddr[10]), .B2(n12), .C1(
        raddr[21]), .C2(n13), .ZN(n335) );
  AOI222 U305 ( .A1(raddr[61]), .A2(n260), .B1(raddr[39]), .B2(n245), 
        .C1(raddr[50]), .C2(n10), .ZN(n310) );
  AOI222 U306 ( .A1(raddr[63]), .A2(n260), .B1(raddr[41]), .B2(n245), 
        .C1(raddr[52]), .C2(n10), .ZN(n302) );
  AOI222 U307 ( .A1(raddr[96]), .A2(n7), .B1(raddr[74]), .B2(n8), .C1(
        raddr[85]), .C2(n9), .ZN(n301) );
  NAND4 U308 ( .A1(n300), .A2(n301), .A3(n302), .A4(n303), .ZN(addrb[8]) );
  AOI22 U309 ( .A1(raddr[107]), .A2(n289), .B1(raddr[118]), .B2(n295), 
        .ZN(n300) );
  MOAI22 U310 ( .A1(n146), .A2(n143), .B1(n143), .B2(raddr[19]), .ZN(n404) );
  NOR2 U311 ( .A1(n144), .A2(N754), .ZN(n146) );
  MOAI22 U312 ( .A1(n226), .A2(n143), .B1(n143), .B2(waddr[19]), .ZN(n525) );
  NOR2 U313 ( .A1(n224), .A2(N334), .ZN(n226) );
  MOAI22 U314 ( .A1(n204), .A2(n202), .B1(n202), .B2(raddr[105]), .ZN(
        n494) );
  NOR2 U315 ( .A1(n205), .A2(N568), .ZN(n204) );
  MOAI22 U316 ( .A1(n284), .A2(n202), .B1(n202), .B2(waddr[105]), .ZN(
        n615) );
  NOR2 U317 ( .A1(n285), .A2(N148), .ZN(n284) );
  MOAI22 U318 ( .A1(n158), .A2(n159), .B1(n159), .B2(raddr[42]), .ZN(n425) );
  NOR2 U319 ( .A1(n160), .A2(N709), .ZN(n158) );
  MOAI22 U320 ( .A1(n161), .A2(n159), .B1(n159), .B2(raddr[41]), .ZN(n426) );
  NOR2 U321 ( .A1(n160), .A2(N708), .ZN(n161) );
  MOAI22 U322 ( .A1(n239), .A2(n159), .B1(n159), .B2(waddr[42]), .ZN(n546) );
  NOR2 U323 ( .A1(n240), .A2(N289), .ZN(n239) );
  MOAI22 U324 ( .A1(n241), .A2(n159), .B1(n159), .B2(waddr[41]), .ZN(n547) );
  NOR2 U325 ( .A1(n240), .A2(N288), .ZN(n241) );
  MOAI22 U326 ( .A1(n190), .A2(n188), .B1(n188), .B2(raddr[85]), .ZN(n470) );
  NOR2 U327 ( .A1(n191), .A2(N616), .ZN(n190) );
  MOAI22 U328 ( .A1(n197), .A2(n195), .B1(n195), .B2(raddr[95]), .ZN(n482) );
  NOR2 U329 ( .A1(n198), .A2(N592), .ZN(n197) );
  MOAI22 U330 ( .A1(n270), .A2(n188), .B1(n188), .B2(waddr[85]), .ZN(n591) );
  NOR2 U331 ( .A1(n271), .A2(N196), .ZN(n270) );
  MOAI22 U332 ( .A1(n277), .A2(n195), .B1(n195), .B2(waddr[95]), .ZN(n603) );
  NOR2 U333 ( .A1(n278), .A2(N172), .ZN(n277) );
  MOAI22 U334 ( .A1(n182), .A2(n180), .B1(n180), .B2(raddr[74]), .ZN(n459) );
  NOR2 U335 ( .A1(n183), .A2(N639), .ZN(n182) );
  MOAI22 U336 ( .A1(n184), .A2(n180), .B1(n180), .B2(raddr[73]), .ZN(n460) );
  NOR2 U337 ( .A1(n183), .A2(N638), .ZN(n184) );
  MOAI22 U338 ( .A1(n262), .A2(n180), .B1(n180), .B2(waddr[74]), .ZN(n580) );
  NOR2 U339 ( .A1(n263), .A2(N219), .ZN(n262) );
  MOAI22 U340 ( .A1(n264), .A2(n180), .B1(n180), .B2(waddr[73]), .ZN(n581) );
  NOR2 U341 ( .A1(n263), .A2(N218), .ZN(n264) );
  MOAI22 U342 ( .A1(n175), .A2(n173), .B1(n173), .B2(raddr[64]), .ZN(n447) );
  NOR2 U343 ( .A1(n176), .A2(N663), .ZN(n175) );
  MOAI22 U344 ( .A1(n255), .A2(n173), .B1(n173), .B2(waddr[64]), .ZN(n568) );
  NOR2 U345 ( .A1(n256), .A2(N243), .ZN(n255) );
  MOAI22 U346 ( .A1(n134), .A2(n18), .B1(n19), .B2(raddr[10]), .ZN(n391)
         );
  NOR2 U347 ( .A1(n136), .A2(N779), .ZN(n134) );
  MOAI22 U348 ( .A1(n215), .A2(n19), .B1(n135), .B2(waddr[10]), .ZN(n512)
         );
  NOR2 U349 ( .A1(n216), .A2(N359), .ZN(n215) );
  MOAI22 U350 ( .A1(n137), .A2(n18), .B1(n18), .B2(raddr[9]), .ZN(n392)
         );
  NOR2 U351 ( .A1(n136), .A2(N778), .ZN(n137) );
  MOAI22 U352 ( .A1(n167), .A2(n16), .B1(n17), .B2(raddr[53]), .ZN(n436)
         );
  NOR2 U353 ( .A1(n168), .A2(N686), .ZN(n167) );
  MOAI22 U354 ( .A1(n169), .A2(n16), .B1(n16), .B2(raddr[51]), .ZN(n438)
         );
  NOR2 U355 ( .A1(n168), .A2(N684), .ZN(n169) );
  MOAI22 U356 ( .A1(n217), .A2(n18), .B1(n19), .B2(waddr[9]), .ZN(n513)
         );
  NOR2 U357 ( .A1(n216), .A2(N358), .ZN(n217) );
  MOAI22 U358 ( .A1(n247), .A2(n17), .B1(n165), .B2(waddr[53]), .ZN(n557)
         );
  NOR2 U359 ( .A1(n248), .A2(N266), .ZN(n247) );
  MOAI22 U360 ( .A1(n249), .A2(n16), .B1(n17), .B2(waddr[51]), .ZN(n559)
         );
  NOR2 U361 ( .A1(n248), .A2(N264), .ZN(n249) );
  MOAI22 U362 ( .A1(n209), .A2(n116), .B1(N545), .B2(n210), .ZN(n505) );
  MOAI22 U363 ( .A1(n15), .A2(n115), .B1(N544), .B2(n210), .ZN(n506) );
  MOAI22 U364 ( .A1(n209), .A2(n113), .B1(N542), .B2(n210), .ZN(n508) );
  MOAI22 U365 ( .A1(n15), .A2(n112), .B1(N541), .B2(n210), .ZN(n509) );
  MOAI22 U366 ( .A1(n209), .A2(n110), .B1(N539), .B2(n210), .ZN(n511) );
  MOAI22 U367 ( .A1(n15), .A2(n60), .B1(N129), .B2(n290), .ZN(n622) );
  MOAI22 U368 ( .A1(n209), .A2(n55), .B1(N124), .B2(n290), .ZN(n627) );
  MOAI22 U369 ( .A1(n15), .A2(n54), .B1(N123), .B2(n290), .ZN(n628) );
  MOAI22 U370 ( .A1(n209), .A2(n52), .B1(N121), .B2(n290), .ZN(n630) );
  MOAI22 U371 ( .A1(n15), .A2(n51), .B1(N120), .B2(n290), .ZN(n631) );
  MOAI22 U372 ( .A1(n14), .A2(n120), .B1(N549), .B2(n210), .ZN(n501) );
  MOAI22 U373 ( .A1(n14), .A2(n114), .B1(N543), .B2(n210), .ZN(n507) );
  MOAI22 U374 ( .A1(n14), .A2(n111), .B1(N540), .B2(n210), .ZN(n510) );
  MOAI22 U375 ( .A1(n14), .A2(n56), .B1(N125), .B2(n290), .ZN(n626) );
  MOAI22 U376 ( .A1(n14), .A2(n53), .B1(N122), .B2(n290), .ZN(n629) );
  MOAI22 U377 ( .A1(n14), .A2(n50), .B1(N119), .B2(n290), .ZN(n632) );
  OAI22 U378 ( .A1(n676), .A2(n663), .B1(n142), .B2(n143), .ZN(n402) );
  NOR2 U379 ( .A1(n144), .A2(N756), .ZN(n142) );
  OAI22 U380 ( .A1(n676), .A2(n105), .B1(n223), .B2(n143), .ZN(n523) );
  NOR2 U381 ( .A1(n224), .A2(N336), .ZN(n223) );
  MOAI22 U382 ( .A1(n674), .A2(n653), .B1(N710), .B2(n157), .ZN(n424) );
  MOAI22 U383 ( .A1(n672), .A2(n639), .B1(N654), .B2(n174), .ZN(n456) );
  MOAI22 U384 ( .A1(n674), .A2(n95), .B1(N290), .B2(n238), .ZN(n545) );
  MOAI22 U385 ( .A1(n672), .A2(n81), .B1(N234), .B2(n254), .ZN(n577) );
  MOAI22 U386 ( .A1(n670), .A2(n130), .B1(N608), .B2(n189), .ZN(n478) );
  MOAI22 U387 ( .A1(n670), .A2(n70), .B1(N188), .B2(n269), .ZN(n599) );
  MOAI22 U388 ( .A1(n677), .A2(n664), .B1(N769), .B2(n138), .ZN(n401) );
  MOAI22 U389 ( .A1(n673), .A2(n645), .B1(N677), .B2(n166), .ZN(n445) );
  MOAI22 U390 ( .A1(n668), .A2(n121), .B1(N562), .B2(n203), .ZN(n500) );
  MOAI22 U391 ( .A1(n677), .A2(n106), .B1(N349), .B2(n218), .ZN(n522) );
  MOAI22 U392 ( .A1(n673), .A2(n87), .B1(N257), .B2(n246), .ZN(n566) );
  MOAI22 U393 ( .A1(n668), .A2(n61), .B1(N142), .B2(n283), .ZN(n621) );
  OAI22 U394 ( .A1(n675), .A2(n658), .B1(n150), .B2(n151), .ZN(n413) );
  I_NOR2 U395 ( .A1(n152), .B1(N733), .ZN(n150) );
  OAI22 U396 ( .A1(n675), .A2(n100), .B1(n231), .B2(n151), .ZN(n534) );
  I_NOR2 U397 ( .A1(n232), .B1(N313), .ZN(n231) );
  AND2 U398 ( .A1(n209), .A2(n211), .Z(n210) );
  NAND4 U399 ( .A1(raddr[114]), .A2(n110), .A3(n212), .A4(n213), .ZN(n211)
         );
  NOR3 U400 ( .A1(raddr[120]), .A2(raddr[112]), .A3(raddr[111]), .ZN(n212)
         );
  NOR4 U401 ( .A1(n214), .A2(raddr[113]), .A3(raddr[116]), .A4(raddr[115]), 
        .ZN(n213) );
  AND2 U402 ( .A1(n15), .A2(n291), .Z(n290) );
  NAND4 U403 ( .A1(waddr[114]), .A2(n50), .A3(n292), .A4(n293), .ZN(n291)
         );
  NOR3 U404 ( .A1(waddr[120]), .A2(waddr[112]), .A3(waddr[111]), .ZN(n292)
         );
  NOR4 U405 ( .A1(n294), .A2(waddr[113]), .A3(waddr[116]), .A4(waddr[115]), 
        .ZN(n293) );
  AO22 U406 ( .A1(n151), .A2(raddr[22]), .B1(N723), .B2(n153), .Z(n423)
         );
  AO22 U407 ( .A1(n195), .A2(raddr[88]), .B1(N585), .B2(n196), .Z(n489)
         );
  AO22 U408 ( .A1(n151), .A2(waddr[22]), .B1(N303), .B2(n233), .Z(n544)
         );
  AO22 U409 ( .A1(n195), .A2(waddr[88]), .B1(N165), .B2(n276), .Z(n610)
         );
  AO22 U410 ( .A1(n180), .A2(raddr[66]), .B1(N631), .B2(n181), .Z(n467)
         );
  AO22 U411 ( .A1(n180), .A2(waddr[66]), .B1(N211), .B2(n261), .Z(n588)
         );
  AO22 U412 ( .A1(n143), .A2(raddr[17]), .B1(N752), .B2(n145), .Z(n406)
         );
  AO22 U413 ( .A1(n16), .A2(raddr[47]), .B1(N680), .B2(n166), .Z(n442) );
  AO22 U414 ( .A1(n188), .A2(raddr[80]), .B1(N611), .B2(n189), .Z(n475)
         );
  AO22 U415 ( .A1(n143), .A2(waddr[17]), .B1(N332), .B2(n225), .Z(n527)
         );
  AO22 U416 ( .A1(n17), .A2(waddr[47]), .B1(N260), .B2(n246), .Z(n563) );
  AO22 U417 ( .A1(n188), .A2(waddr[80]), .B1(N191), .B2(n269), .Z(n596)
         );
  AO22 U418 ( .A1(n143), .A2(raddr[11]), .B1(N746), .B2(n145), .Z(n412)
         );
  AO22 U419 ( .A1(n143), .A2(waddr[11]), .B1(N326), .B2(n225), .Z(n533)
         );
  AO22 U420 ( .A1(n18), .A2(raddr[6]), .B1(N775), .B2(n138), .Z(n395) );
  AO22 U421 ( .A1(n151), .A2(raddr[24]), .B1(N725), .B2(n153), .Z(n421)
         );
  AO22 U422 ( .A1(n159), .A2(raddr[38]), .B1(N705), .B2(n157), .Z(n429)
         );
  AO22 U423 ( .A1(n173), .A2(raddr[56]), .B1(N655), .B2(n174), .Z(n455)
         );
  AO22 U424 ( .A1(n195), .A2(raddr[90]), .B1(N587), .B2(n196), .Z(n487)
         );
  AO22 U425 ( .A1(n202), .A2(raddr[102]), .B1(N565), .B2(n203), .Z(n497)
         );
  AO22 U426 ( .A1(n19), .A2(waddr[6]), .B1(N355), .B2(n218), .Z(n516) );
  AO22 U427 ( .A1(n151), .A2(waddr[24]), .B1(N305), .B2(n233), .Z(n542)
         );
  AO22 U428 ( .A1(n159), .A2(waddr[38]), .B1(N285), .B2(n238), .Z(n550)
         );
  AO22 U429 ( .A1(n173), .A2(waddr[56]), .B1(N235), .B2(n254), .Z(n576)
         );
  AO22 U430 ( .A1(n195), .A2(waddr[90]), .B1(N167), .B2(n276), .Z(n608)
         );
  AO22 U431 ( .A1(n202), .A2(waddr[102]), .B1(N145), .B2(n283), .Z(n618)
         );
  AO22 U432 ( .A1(n159), .A2(raddr[33]), .B1(N700), .B2(n157), .Z(n434)
         );
  AO22 U433 ( .A1(n159), .A2(waddr[33]), .B1(N280), .B2(n238), .Z(n555)
         );
  AO22 U434 ( .A1(n143), .A2(raddr[20]), .B1(N755), .B2(n145), .Z(n403)
         );
  AO22 U435 ( .A1(n17), .A2(raddr[52]), .B1(N685), .B2(n166), .Z(n437) );
  AO22 U436 ( .A1(n188), .A2(raddr[81]), .B1(N612), .B2(n189), .Z(n474)
         );
  AO22 U437 ( .A1(n143), .A2(waddr[20]), .B1(N335), .B2(n225), .Z(n524)
         );
  AO22 U438 ( .A1(n165), .A2(waddr[52]), .B1(N265), .B2(n246), .Z(n558)
         );
  AO22 U439 ( .A1(n188), .A2(waddr[81]), .B1(N192), .B2(n269), .Z(n595)
         );
  AO22 U440 ( .A1(n135), .A2(raddr[8]), .B1(N777), .B2(n138), .Z(n393) );
  AO22 U441 ( .A1(n143), .A2(raddr[15]), .B1(N750), .B2(n145), .Z(n408)
         );
  AO22 U442 ( .A1(n151), .A2(raddr[27]), .B1(N728), .B2(n153), .Z(n418)
         );
  AO22 U443 ( .A1(n159), .A2(raddr[39]), .B1(N706), .B2(n157), .Z(n428)
         );
  AO22 U444 ( .A1(n173), .A2(raddr[58]), .B1(N657), .B2(n174), .Z(n453)
         );
  AO22 U445 ( .A1(n180), .A2(raddr[67]), .B1(N632), .B2(n181), .Z(n466)
         );
  AO22 U446 ( .A1(n188), .A2(raddr[79]), .B1(N610), .B2(n189), .Z(n476)
         );
  AO22 U447 ( .A1(n195), .A2(raddr[91]), .B1(N588), .B2(n196), .Z(n486)
         );
  AO22 U448 ( .A1(n202), .A2(raddr[103]), .B1(N566), .B2(n203), .Z(n496)
         );
  AO22 U449 ( .A1(n18), .A2(waddr[8]), .B1(N357), .B2(n218), .Z(n514) );
  AO22 U450 ( .A1(n143), .A2(waddr[15]), .B1(N330), .B2(n225), .Z(n529)
         );
  AO22 U451 ( .A1(n151), .A2(waddr[27]), .B1(N308), .B2(n233), .Z(n539)
         );
  AO22 U452 ( .A1(n159), .A2(waddr[39]), .B1(N286), .B2(n238), .Z(n549)
         );
  AO22 U453 ( .A1(n173), .A2(waddr[58]), .B1(N237), .B2(n254), .Z(n574)
         );
  AO22 U454 ( .A1(n180), .A2(waddr[67]), .B1(N212), .B2(n261), .Z(n587)
         );
  AO22 U455 ( .A1(n188), .A2(waddr[79]), .B1(N190), .B2(n269), .Z(n597)
         );
  AO22 U456 ( .A1(n195), .A2(waddr[91]), .B1(N168), .B2(n276), .Z(n607)
         );
  AO22 U457 ( .A1(n202), .A2(waddr[103]), .B1(N146), .B2(n283), .Z(n617)
         );
  AO22 U458 ( .A1(n202), .A2(raddr[100]), .B1(N563), .B2(n203), .Z(n499)
         );
  AO22 U459 ( .A1(n202), .A2(waddr[100]), .B1(N143), .B2(n283), .Z(n620)
         );
  AO22 U460 ( .A1(n135), .A2(raddr[2]), .B1(N771), .B2(n138), .Z(n399) );
  AO22 U461 ( .A1(n151), .A2(raddr[23]), .B1(N724), .B2(n153), .Z(n422)
         );
  AO22 U462 ( .A1(n159), .A2(raddr[37]), .B1(N704), .B2(n157), .Z(n430)
         );
  AO22 U463 ( .A1(n202), .A2(raddr[101]), .B1(N564), .B2(n203), .Z(n498)
         );
  AO22 U464 ( .A1(n18), .A2(waddr[2]), .B1(N351), .B2(n218), .Z(n520) );
  AO22 U465 ( .A1(n151), .A2(waddr[23]), .B1(N304), .B2(n233), .Z(n543)
         );
  AO22 U466 ( .A1(n159), .A2(waddr[37]), .B1(N284), .B2(n238), .Z(n551)
         );
  AO22 U467 ( .A1(n202), .A2(waddr[101]), .B1(N144), .B2(n283), .Z(n619)
         );
  AO22 U468 ( .A1(n165), .A2(raddr[46]), .B1(N679), .B2(n166), .Z(n443)
         );
  AO22 U469 ( .A1(n16), .A2(waddr[46]), .B1(N259), .B2(n246), .Z(n564) );
  AO22 U470 ( .A1(n17), .A2(raddr[45]), .B1(N678), .B2(n166), .Z(n444) );
  AO22 U471 ( .A1(n165), .A2(waddr[45]), .B1(N258), .B2(n246), .Z(n565)
         );
  AO22 U472 ( .A1(n180), .A2(raddr[76]), .B1(N641), .B2(n181), .Z(n457)
         );
  AO22 U473 ( .A1(n180), .A2(waddr[76]), .B1(N221), .B2(n261), .Z(n578)
         );
  AO22 U474 ( .A1(n202), .A2(raddr[109]), .B1(N572), .B2(n203), .Z(n490)
         );
  AO22 U475 ( .A1(n202), .A2(waddr[109]), .B1(N152), .B2(n283), .Z(n611)
         );
  AO22 U476 ( .A1(n19), .A2(raddr[1]), .B1(N770), .B2(n138), .Z(n400) );
  AO22 U477 ( .A1(n135), .A2(waddr[1]), .B1(N350), .B2(n218), .Z(n521) );
  AO22 U478 ( .A1(n151), .A2(raddr[29]), .B1(N730), .B2(n153), .Z(n416)
         );
  AO22 U479 ( .A1(n151), .A2(raddr[26]), .B1(N727), .B2(n153), .Z(n419)
         );
  AO22 U480 ( .A1(n151), .A2(waddr[29]), .B1(N310), .B2(n233), .Z(n537)
         );
  AO22 U481 ( .A1(n151), .A2(waddr[26]), .B1(N307), .B2(n233), .Z(n540)
         );
  AO22 U482 ( .A1(n188), .A2(raddr[87]), .B1(N618), .B2(n189), .Z(n468)
         );
  AO22 U483 ( .A1(n188), .A2(waddr[87]), .B1(N198), .B2(n269), .Z(n589)
         );
  AO22 U484 ( .A1(n165), .A2(raddr[54]), .B1(N687), .B2(n166), .Z(n435)
         );
  AO22 U485 ( .A1(n16), .A2(waddr[54]), .B1(N267), .B2(n246), .Z(n556) );
  AO22 U486 ( .A1(n173), .A2(raddr[65]), .B1(N664), .B2(n174), .Z(n446)
         );
  AO22 U487 ( .A1(n195), .A2(raddr[98]), .B1(N595), .B2(n196), .Z(n479)
         );
  AO22 U488 ( .A1(n173), .A2(waddr[65]), .B1(N244), .B2(n254), .Z(n567)
         );
  AO22 U489 ( .A1(n195), .A2(waddr[98]), .B1(N175), .B2(n276), .Z(n600)
         );
  AO22 U490 ( .A1(n143), .A2(raddr[18]), .B1(N753), .B2(n145), .Z(n405)
         );
  AO22 U491 ( .A1(n188), .A2(raddr[83]), .B1(N614), .B2(n189), .Z(n472)
         );
  AO22 U492 ( .A1(n143), .A2(waddr[18]), .B1(N333), .B2(n225), .Z(n526)
         );
  AO22 U493 ( .A1(n188), .A2(waddr[83]), .B1(N194), .B2(n269), .Z(n593)
         );
  AO22 U494 ( .A1(n19), .A2(raddr[7]), .B1(N776), .B2(n138), .Z(n394) );
  AO22 U495 ( .A1(n173), .A2(raddr[61]), .B1(N660), .B2(n174), .Z(n450)
         );
  AO22 U496 ( .A1(n195), .A2(raddr[93]), .B1(N590), .B2(n196), .Z(n484)
         );
  AO22 U497 ( .A1(n202), .A2(raddr[104]), .B1(N567), .B2(n203), .Z(n495)
         );
  AO22 U498 ( .A1(n135), .A2(waddr[7]), .B1(N356), .B2(n218), .Z(n515) );
  AO22 U499 ( .A1(n173), .A2(waddr[61]), .B1(N240), .B2(n254), .Z(n571)
         );
  AO22 U500 ( .A1(n195), .A2(waddr[93]), .B1(N170), .B2(n276), .Z(n605)
         );
  AO22 U501 ( .A1(n202), .A2(waddr[104]), .B1(N147), .B2(n283), .Z(n616)
         );
  NAND4 U502 ( .A1(raddr[29]), .A2(raddr[26]), .A3(n154), .A4(n155), .ZN(
        n152) );
  NOR3 U503 ( .A1(n654), .A2(raddr[22]), .A3(n658), .ZN(n154) );
  NOR4 U504 ( .A1(n156), .A2(raddr[23]), .A3(raddr[27]), .A4(raddr[24]), 
        .ZN(n155) );
  NAND3 U505 ( .A1(n656), .A2(n657), .A3(n655), .ZN(n156) );
  NAND4 U506 ( .A1(waddr[29]), .A2(waddr[26]), .A3(n234), .A4(n235), .ZN(
        n232) );
  NOR3 U507 ( .A1(n96), .A2(waddr[22]), .A3(n100), .ZN(n234) );
  NOR4 U508 ( .A1(n236), .A2(waddr[23]), .A3(waddr[27]), .A4(waddr[24]), 
        .ZN(n235) );
  NAND3 U509 ( .A1(n98), .A2(n99), .A3(n97), .ZN(n236) );
  AND4 U510 ( .A1(raddr[64]), .A2(raddr[61]), .A3(n177), .A4(n178), .Z(
        n176) );
  NOR3 U511 ( .A1(n642), .A2(n639), .A3(n640), .ZN(n177) );
  NOR4 U512 ( .A1(n179), .A2(raddr[65]), .A3(raddr[58]), .A4(raddr[56]), 
        .ZN(n178) );
  NAND3 U513 ( .A1(n643), .A2(n644), .A3(n641), .ZN(n179) );
  AND4 U514 ( .A1(waddr[64]), .A2(waddr[61]), .A3(n257), .A4(n258), .Z(
        n256) );
  NOR3 U515 ( .A1(n84), .A2(n81), .A3(n82), .ZN(n257) );
  NOR4 U516 ( .A1(n259), .A2(waddr[65]), .A3(waddr[58]), .A4(waddr[56]), 
        .ZN(n258) );
  NAND3 U517 ( .A1(n85), .A2(n86), .A3(n83), .ZN(n259) );
  AND4 U518 ( .A1(raddr[53]), .A2(raddr[51]), .A3(n170), .A4(n171), .Z(
        n168) );
  NOR3 U519 ( .A1(n648), .A2(n646), .A3(n647), .ZN(n170) );
  NOR4 U520 ( .A1(n172), .A2(raddr[54]), .A3(raddr[52]), .A4(raddr[47]), 
        .ZN(n171) );
  NAND3 U521 ( .A1(raddr[45]), .A2(n645), .A3(raddr[46]), .ZN(n172) );
  AND4 U522 ( .A1(raddr[74]), .A2(raddr[73]), .A3(n185), .A4(n186), .Z(
        n183) );
  NOR3 U523 ( .A1(n637), .A2(n633), .A3(n635), .ZN(n185) );
  NOR4 U524 ( .A1(n187), .A2(raddr[66]), .A3(raddr[67]), .A4(raddr[76]), 
        .ZN(n186) );
  NAND3 U525 ( .A1(n636), .A2(n638), .A3(n634), .ZN(n187) );
  AND4 U526 ( .A1(waddr[53]), .A2(waddr[51]), .A3(n250), .A4(n251), .Z(
        n248) );
  NOR3 U527 ( .A1(n90), .A2(n88), .A3(n89), .ZN(n250) );
  NOR4 U528 ( .A1(n252), .A2(waddr[54]), .A3(waddr[52]), .A4(waddr[47]), 
        .ZN(n251) );
  NAND3 U529 ( .A1(waddr[45]), .A2(n87), .A3(waddr[46]), .ZN(n252) );
  AND4 U530 ( .A1(waddr[74]), .A2(waddr[73]), .A3(n265), .A4(n266), .Z(
        n263) );
  NOR3 U531 ( .A1(n79), .A2(n75), .A3(n77), .ZN(n265) );
  NOR4 U532 ( .A1(n267), .A2(waddr[66]), .A3(waddr[67]), .A4(waddr[76]), 
        .ZN(n266) );
  NAND3 U533 ( .A1(n78), .A2(n80), .A3(n76), .ZN(n267) );
  AND4 U534 ( .A1(raddr[9]), .A2(raddr[7]), .A3(n139), .A4(n140), .Z(n136)
         );
  NOR3 U535 ( .A1(n667), .A2(n665), .A3(n666), .ZN(n139) );
  NOR4 U536 ( .A1(n141), .A2(raddr[2]), .A3(raddr[8]), .A4(raddr[6]), .ZN(
        n140) );
  NAND3 U537 ( .A1(raddr[10]), .A2(n664), .A3(raddr[1]), .ZN(n141) );
  AND4 U538 ( .A1(raddr[19]), .A2(raddr[18]), .A3(n147), .A4(n148), .Z(
        n144) );
  NOR3 U539 ( .A1(n662), .A2(n663), .A3(n661), .ZN(n147) );
  NOR4 U540 ( .A1(n149), .A2(raddr[15]), .A3(raddr[20]), .A4(raddr[17]), 
        .ZN(n148) );
  NAND3 U541 ( .A1(n659), .A2(n660), .A3(raddr[11]), .ZN(n149) );
  AND4 U542 ( .A1(waddr[9]), .A2(waddr[7]), .A3(n219), .A4(n220), .Z(n216)
         );
  NOR3 U543 ( .A1(n109), .A2(n107), .A3(n108), .ZN(n219) );
  NOR4 U544 ( .A1(n221), .A2(waddr[2]), .A3(waddr[8]), .A4(waddr[6]), .ZN(
        n220) );
  NAND3 U545 ( .A1(waddr[10]), .A2(n106), .A3(waddr[1]), .ZN(n221) );
  AND4 U546 ( .A1(waddr[19]), .A2(waddr[18]), .A3(n227), .A4(n228), .Z(
        n224) );
  NOR3 U547 ( .A1(n104), .A2(n105), .A3(n103), .ZN(n227) );
  NOR4 U548 ( .A1(n229), .A2(waddr[15]), .A3(waddr[20]), .A4(waddr[17]), 
        .ZN(n228) );
  NAND3 U549 ( .A1(n101), .A2(n102), .A3(waddr[11]), .ZN(n229) );
  AND4 U550 ( .A1(raddr[85]), .A2(raddr[83]), .A3(n192), .A4(n193), .Z(
        n191) );
  NOR3 U551 ( .A1(n131), .A2(raddr[87]), .A3(n130), .ZN(n192) );
  NOR4 U552 ( .A1(n194), .A2(raddr[79]), .A3(raddr[81]), .A4(raddr[80]), 
        .ZN(n193) );
  NAND3 U553 ( .A1(n133), .A2(n296), .A3(n132), .ZN(n194) );
  AND4 U554 ( .A1(raddr[95]), .A2(raddr[93]), .A3(n199), .A4(n200), .Z(
        n198) );
  NOR3 U555 ( .A1(n126), .A2(raddr[88]), .A3(n125), .ZN(n199) );
  NOR4 U556 ( .A1(n201), .A2(raddr[98]), .A3(raddr[91]), .A4(raddr[90]), 
        .ZN(n200) );
  NAND3 U557 ( .A1(n128), .A2(n129), .A3(n127), .ZN(n201) );
  AND4 U558 ( .A1(raddr[105]), .A2(raddr[104]), .A3(n206), .A4(n207), .Z(
        n205) );
  NOR3 U559 ( .A1(n121), .A2(raddr[100]), .A3(raddr[109]), .ZN(n206) );
  NOR4 U560 ( .A1(n208), .A2(raddr[101]), .A3(raddr[103]), .A4(raddr[102]), .ZN(n207) );
  NAND3 U561 ( .A1(n123), .A2(n124), .A3(n122), .ZN(n208) );
  AND4 U562 ( .A1(waddr[85]), .A2(waddr[83]), .A3(n272), .A4(n273), .Z(n271) );
  NOR3 U563 ( .A1(n71), .A2(waddr[87]), .A3(n70), .ZN(n272) );
  NOR4 U564 ( .A1(n274), .A2(waddr[79]), .A3(waddr[81]), .A4(waddr[80]), .ZN(n273) );
  NAND3 U565 ( .A1(n73), .A2(n74), .A3(n72), .ZN(n274) );
  AND4 U566 ( .A1(waddr[95]), .A2(waddr[93]), .A3(n279), .A4(n280), .Z(n278) );
  NOR3 U567 ( .A1(n66), .A2(waddr[88]), .A3(n65), .ZN(n279) );
  NOR4 U568 ( .A1(n281), .A2(waddr[98]), .A3(waddr[91]), .A4(waddr[90]), .ZN(n280) );
  NAND3 U569 ( .A1(n68), .A2(n69), .A3(n67), .ZN(n281) );
  AND4 U570 ( .A1(waddr[105]), .A2(waddr[104]), .A3(n286), .A4(n287), .Z(n285) );
  NOR3 U571 ( .A1(n61), .A2(waddr[100]), .A3(waddr[109]), .ZN(n286) );
  NOR4 U572 ( .A1(n288), .A2(waddr[101]), .A3(waddr[103]), .A4(waddr[102]), .ZN(n287) );
  NAND3 U573 ( .A1(n63), .A2(n64), .A3(n62), .ZN(n288) );
  AND4 U574 ( .A1(raddr[42]), .A2(raddr[41]), .A3(n162), .A4(n163), .Z(n160) );
  NOR3 U575 ( .A1(n652), .A2(n649), .A3(n650), .ZN(n162) );
  NOR4 U576 ( .A1(n164), .A2(raddr[37]), .A3(raddr[39]), .A4(raddr[38]), .ZN(n163) );
  NAND3 U577 ( .A1(n653), .A2(n651), .A3(raddr[33]), .ZN(n164) );
  AND4 U578 ( .A1(waddr[42]), .A2(waddr[41]), .A3(n242), .A4(n243), .Z(n240) );
  NOR3 U579 ( .A1(n94), .A2(n91), .A3(n92), .ZN(n242) );
  NOR4 U580 ( .A1(n244), .A2(waddr[37]), .A3(waddr[39]), .A4(waddr[38]), .ZN(n243) );
  NAND3 U581 ( .A1(n95), .A2(n93), .A3(waddr[33]), .ZN(n244) );
  INV U582 ( .I(waddr[110]), .ZN(n50) );
  INV U583 ( .I(waddr[111]), .ZN(n51) );
  INV U584 ( .I(waddr[112]), .ZN(n52) );
  INV U585 ( .I(waddr[113]), .ZN(n53) );
  INV U586 ( .I(waddr[114]), .ZN(n54) );
  INV U587 ( .I(waddr[115]), .ZN(n55) );
  INV U588 ( .I(waddr[116]), .ZN(n56) );
  INV U589 ( .I(waddr[117]), .ZN(n57) );
  INV U590 ( .I(waddr[118]), .ZN(n58) );
  INV U591 ( .I(waddr[119]), .ZN(n59) );
  INV U592 ( .I(waddr[120]), .ZN(n60) );
  INV U593 ( .I(waddr[99]), .ZN(n61) );
  INV U594 ( .I(waddr[106]), .ZN(n62) );
  INV U595 ( .I(waddr[107]), .ZN(n63) );
  INV U596 ( .I(waddr[108]), .ZN(n64) );
  INV U597 ( .I(waddr[89]), .ZN(n65) );
  INV U598 ( .I(waddr[92]), .ZN(n66) );
  INV U599 ( .I(waddr[94]), .ZN(n67) );
  INV U600 ( .I(waddr[96]), .ZN(n68) );
  INV U601 ( .I(waddr[97]), .ZN(n69) );
  INV U602 ( .I(waddr[77]), .ZN(n70) );
  INV U603 ( .I(waddr[78]), .ZN(n71) );
  INV U604 ( .I(waddr[82]), .ZN(n72) );
  INV U605 ( .I(waddr[84]), .ZN(n73) );
  INV U606 ( .I(waddr[86]), .ZN(n74) );
  INV U607 ( .I(waddr[68]), .ZN(n75) );
  INV U608 ( .I(waddr[69]), .ZN(n76) );
  INV U609 ( .I(waddr[70]), .ZN(n77) );
  INV U610 ( .I(waddr[71]), .ZN(n78) );
  INV U611 ( .I(waddr[72]), .ZN(n79) );
  INV U612 ( .I(waddr[75]), .ZN(n80) );
  INV U613 ( .I(waddr[55]), .ZN(n81) );
  INV U614 ( .I(waddr[57]), .ZN(n82) );
  INV U615 ( .I(waddr[59]), .ZN(n83) );
  INV U616 ( .I(waddr[60]), .ZN(n84) );
  INV U617 ( .I(waddr[62]), .ZN(n85) );
  INV U618 ( .I(waddr[63]), .ZN(n86) );
  INV U619 ( .I(waddr[44]), .ZN(n87) );
  INV U620 ( .I(waddr[48]), .ZN(n88) );
  INV U621 ( .I(waddr[49]), .ZN(n89) );
  INV U622 ( .I(waddr[50]), .ZN(n90) );
  INV U623 ( .I(waddr[34]), .ZN(n91) );
  INV U624 ( .I(waddr[35]), .ZN(n92) );
  INV U625 ( .I(waddr[36]), .ZN(n93) );
  INV U626 ( .I(waddr[40]), .ZN(n94) );
  INV U627 ( .I(waddr[43]), .ZN(n95) );
  INV U628 ( .I(waddr[25]), .ZN(n96) );
  INV U629 ( .I(waddr[28]), .ZN(n97) );
  INV U630 ( .I(waddr[30]), .ZN(n98) );
  INV U631 ( .I(waddr[31]), .ZN(n99) );
  INV U632 ( .I(waddr[32]), .ZN(n100) );
  INV U633 ( .I(waddr[12]), .ZN(n101) );
  INV U634 ( .I(waddr[13]), .ZN(n102) );
  INV U635 ( .I(waddr[14]), .ZN(n103) );
  INV U636 ( .I(waddr[16]), .ZN(n104) );
  INV U637 ( .I(waddr[21]), .ZN(n105) );
  INV U638 ( .I(waddr[0]), .ZN(n106) );
  INV U639 ( .I(waddr[3]), .ZN(n107) );
  INV U640 ( .I(waddr[4]), .ZN(n108) );
  INV U641 ( .I(waddr[5]), .ZN(n109) );
  INV U642 ( .I(raddr[110]), .ZN(n110) );
  INV U643 ( .I(raddr[111]), .ZN(n111) );
  INV U644 ( .I(raddr[112]), .ZN(n112) );
  INV U645 ( .I(raddr[113]), .ZN(n113) );
  INV U646 ( .I(raddr[114]), .ZN(n114) );
  INV U647 ( .I(raddr[115]), .ZN(n115) );
  INV U648 ( .I(raddr[116]), .ZN(n116) );
  INV U649 ( .I(raddr[117]), .ZN(n117) );
  INV U650 ( .I(raddr[118]), .ZN(n118) );
  INV U651 ( .I(raddr[119]), .ZN(n119) );
  INV U652 ( .I(raddr[120]), .ZN(n120) );
  INV U653 ( .I(raddr[99]), .ZN(n121) );
  INV U654 ( .I(raddr[106]), .ZN(n122) );
  INV U655 ( .I(raddr[107]), .ZN(n123) );
  INV U656 ( .I(raddr[108]), .ZN(n124) );
  INV U657 ( .I(raddr[89]), .ZN(n125) );
  INV U658 ( .I(raddr[92]), .ZN(n126) );
  INV U659 ( .I(raddr[94]), .ZN(n127) );
  INV U660 ( .I(raddr[96]), .ZN(n128) );
  INV U661 ( .I(raddr[97]), .ZN(n129) );
  INV U662 ( .I(raddr[77]), .ZN(n130) );
  INV U663 ( .I(raddr[78]), .ZN(n131) );
  INV U664 ( .I(raddr[82]), .ZN(n132) );
  INV U665 ( .I(raddr[84]), .ZN(n133) );
  INV U666 ( .I(raddr[86]), .ZN(n296) );
  INV U667 ( .I(raddr[68]), .ZN(n633) );
  INV U668 ( .I(raddr[69]), .ZN(n634) );
  INV U669 ( .I(raddr[70]), .ZN(n635) );
  INV U670 ( .I(raddr[71]), .ZN(n636) );
  INV U671 ( .I(raddr[72]), .ZN(n637) );
  INV U672 ( .I(raddr[75]), .ZN(n638) );
  INV U673 ( .I(raddr[55]), .ZN(n639) );
  INV U674 ( .I(raddr[57]), .ZN(n640) );
  INV U675 ( .I(raddr[59]), .ZN(n641) );
  INV U676 ( .I(raddr[60]), .ZN(n642) );
  INV U677 ( .I(raddr[62]), .ZN(n643) );
  INV U678 ( .I(raddr[63]), .ZN(n644) );
  INV U679 ( .I(raddr[44]), .ZN(n645) );
  INV U680 ( .I(raddr[48]), .ZN(n646) );
  INV U681 ( .I(raddr[49]), .ZN(n647) );
  INV U682 ( .I(raddr[50]), .ZN(n648) );
  INV U683 ( .I(raddr[34]), .ZN(n649) );
  INV U684 ( .I(raddr[35]), .ZN(n650) );
  INV U685 ( .I(raddr[36]), .ZN(n651) );
  INV U686 ( .I(raddr[40]), .ZN(n652) );
  INV U687 ( .I(raddr[43]), .ZN(n653) );
  INV U688 ( .I(raddr[25]), .ZN(n654) );
  INV U689 ( .I(raddr[28]), .ZN(n655) );
  INV U690 ( .I(raddr[30]), .ZN(n656) );
  INV U691 ( .I(raddr[31]), .ZN(n657) );
  INV U692 ( .I(raddr[32]), .ZN(n658) );
  INV U693 ( .I(raddr[12]), .ZN(n659) );
  INV U694 ( .I(raddr[13]), .ZN(n660) );
  INV U695 ( .I(raddr[14]), .ZN(n661) );
  INV U696 ( .I(raddr[16]), .ZN(n662) );
  INV U697 ( .I(raddr[21]), .ZN(n663) );
  INV U698 ( .I(raddr[0]), .ZN(n664) );
  INV U699 ( .I(raddr[3]), .ZN(n665) );
  INV U700 ( .I(raddr[4]), .ZN(n666) );
  INV U701 ( .I(raddr[5]), .ZN(n667) );
  INV U702 ( .I(sel[1]), .ZN(n678) );
  INV U703 ( .I(sel[0]), .ZN(n679) );
endmodule


module count_WIDTH8 ( clk, rst_n, ld_n, up_dn, cen, din, tc, zero, cnt_out );
  input [7:0] din;
  output [7:0] cnt_out;
  input clk, rst_n, ld_n, up_dn, cen;
  output tc, zero;
  wire   N11, N12, N13, N14, N15, N16, N17, N18, N19, N20, N21, N22, N23, N24,
         N25, N26, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n34, n1, n2, n35, n36, n37, n38, n39, n40;

  DFF_RST cnt_out_reg_0_ ( .D(n34), .CP(clk), .CDN(rst_n), .Q(cnt_out[0]));
  DFF_RST cnt_out_reg_7_ ( .D(n27), .CP(clk), .CDN(rst_n), .Q(cnt_out[7]));
  DFF_RST cnt_out_reg_1_ ( .D(n33), .CP(clk), .CDN(rst_n), .Q(cnt_out[1]));
  DFF_RST cnt_out_reg_2_ ( .D(n32), .CP(clk), .CDN(rst_n), .Q(cnt_out[2]));
  DFF_RST cnt_out_reg_3_ ( .D(n31), .CP(clk), .CDN(rst_n), .Q(cnt_out[3]));
  DFF_RST cnt_out_reg_4_ ( .D(n30), .CP(clk), .CDN(rst_n), .Q(cnt_out[4]));
  DFF_RST cnt_out_reg_5_ ( .D(n29), .CP(clk), .CDN(rst_n), .Q(cnt_out[5]));
  DFF_RST cnt_out_reg_6_ ( .D(n28), .CP(clk), .CDN(rst_n), .Q(cnt_out[6]));
  OR4 U32 ( .A1(cnt_out[0]), .A2(cnt_out[1]), .A3(cnt_out[2]), .A4(cnt_out[3]), .Z(n24) );
  OR4 U33 ( .A1(cnt_out[4]), .A2(cnt_out[5]), .A3(cnt_out[6]), .A4(cnt_out[7]), .Z(n23) );
  count_WIDTH8_DW01_inc_0 add_24 (.A(cnt_out), .SUM({N18, N17, N16, N15, N14, N13, N12, N11}));
  INV U3 ( .I(ld_n), .ZN(n40) );
  NOR2 U4 ( .A1(n7), .A2(n40), .ZN(n22) );
  NOR2 U5 ( .A1(cen), .A2(n40), .ZN(n7) );
  NOR2 U6 ( .A1(n25), .A2(n26), .ZN(tc) );
  I_NOR2 U7 ( .A1(n22), .B1(up_dn), .ZN(n5) );
  AND2 U8 ( .A1(up_dn), .A2(n22), .Z(n6) );
  NAND2 U9 ( .A1(n10), .A2(n11), .ZN(n29) );
  AOI22 U10 ( .A1(N16), .A2(n6), .B1(cnt_out[5]), .B2(n7), .ZN(n10) );
  AOI22 U11 ( .A1(din[5]), .A2(n40), .B1(N24), .B2(n5), .ZN(n11) );
  NAND2 U12 ( .A1(n14), .A2(n15), .ZN(n31) );
  AOI22 U13 ( .A1(N14), .A2(n6), .B1(cnt_out[3]), .B2(n7), .ZN(n14) );
  AOI22 U14 ( .A1(din[3]), .A2(n40), .B1(N22), .B2(n5), .ZN(n15) );
  NAND2 U15 ( .A1(n16), .A2(n17), .ZN(n32) );
  AOI22 U16 ( .A1(N13), .A2(n6), .B1(cnt_out[2]), .B2(n7), .ZN(n16) );
  AOI22 U17 ( .A1(din[2]), .A2(n40), .B1(N21), .B2(n5), .ZN(n17) );
  NAND2 U18 ( .A1(n3), .A2(n4), .ZN(n27) );
  AOI22 U19 ( .A1(N18), .A2(n6), .B1(cnt_out[7]), .B2(n7), .ZN(n3) );
  AOI22 U20 ( .A1(din[7]), .A2(n40), .B1(N26), .B2(n5), .ZN(n4) );
  NOR2 U21 ( .A1(n23), .A2(n24), .ZN(zero) );
  NAND2 U22 ( .A1(n8), .A2(n9), .ZN(n28) );
  AOI22 U23 ( .A1(N17), .A2(n6), .B1(cnt_out[6]), .B2(n7), .ZN(n8) );
  AOI22 U24 ( .A1(din[6]), .A2(n40), .B1(N25), .B2(n5), .ZN(n9) );
  NAND2 U25 ( .A1(n12), .A2(n13), .ZN(n30) );
  AOI22 U26 ( .A1(N15), .A2(n6), .B1(cnt_out[4]), .B2(n7), .ZN(n12) );
  AOI22 U27 ( .A1(din[4]), .A2(n40), .B1(N23), .B2(n5), .ZN(n13) );
  NAND2 U28 ( .A1(n18), .A2(n19), .ZN(n33) );
  AOI22 U29 ( .A1(N12), .A2(n6), .B1(cnt_out[1]), .B2(n7), .ZN(n18) );
  AOI22 U30 ( .A1(din[1]), .A2(n40), .B1(N20), .B2(n5), .ZN(n19) );
  NAND2 U31 ( .A1(n20), .A2(n21), .ZN(n34) );
  AOI22 U34 ( .A1(din[0]), .A2(n40), .B1(N19), .B2(n5), .ZN(n21) );
  AOI22 U35 ( .A1(N11), .A2(n6), .B1(cnt_out[0]), .B2(n7), .ZN(n20) );
  NAND4 U36 ( .A1(cnt_out[0]), .A2(cnt_out[1]), .A3(cnt_out[2]), .A4(cnt_out[3]), .ZN(n26) );
  NAND4 U37 ( .A1(cnt_out[4]), .A2(cnt_out[5]), .A3(cnt_out[6]), .A4(cnt_out[7]), .ZN(n25) );
  I_NAND2 U38 ( .A1(cnt_out[1]), .B1(N19), .ZN(n1) );
  IOA21 U39 ( .A1(cnt_out[0]), .A2(cnt_out[1]), .B(n1), .ZN(N20) );
  OR2 U40 ( .A1(n1), .A2(cnt_out[2]), .Z(n2) );
  IOA21 U41 ( .A1(n1), .A2(cnt_out[2]), .B(n2), .ZN(N21) );
  OR2 U42 ( .A1(n2), .A2(cnt_out[3]), .Z(n35) );
  IOA21 U43 ( .A1(n2), .A2(cnt_out[3]), .B(n35), .ZN(N22) );
  NOR2 U44 ( .A1(n35), .A2(cnt_out[4]), .ZN(n36) );
  AO21 U45 ( .A1(n35), .A2(cnt_out[4]), .B(n36), .Z(N23) );
  NAND2 U46 ( .A1(n36), .A2(n39), .ZN(n37) );
  OAI21 U47 ( .A1(n36), .A2(n39), .B(n37), .ZN(N24) );
  XNOR2 U48 ( .A1(n37), .A2(cnt_out[6]), .ZN(N25) );
  NOR2 U49 ( .A1(cnt_out[6]), .A2(n37), .ZN(n38) );
  XOR2 U50 ( .A1(cnt_out[7]), .A2(n38), .Z(N26) );
  INV U51 ( .I(cnt_out[5]), .ZN(n39) );
  INV U52 ( .I(cnt_out[0]), .ZN(N19) );
endmodule


module rdyacpt_WIDTH8_0 ( clk, reset_n, upstream_rdy, downstream_acpt, 
        upstream_data, downstream_rdy, upstream_acpt, downstream_data );
  input [7:0] upstream_data;
  output [7:0] downstream_data;
  input clk, reset_n, upstream_rdy, downstream_acpt;
  output downstream_rdy, upstream_acpt;
  wire   v1, ready_reg, N3, N29, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n1;
  wire   [7:0] d1;

  DFF_RST v0_reg ( .D(n16), .CP(clk), .CDN(reset_n), .Q(downstream_rdy) );
  DFF_EN d1_reg_7_ ( .D(upstream_data[7]), .E(N29), .CP(clk), .Q(d1[7]) );
  DFF_EN d1_reg_5_ ( .D(upstream_data[5]), .E(N29), .CP(clk), .Q(d1[5]) );
  DFF_EN d1_reg_3_ ( .D(upstream_data[3]), .E(N29), .CP(clk), .Q(d1[3]) );
  DFF_EN d1_reg_1_ ( .D(upstream_data[1]), .E(N29), .CP(clk), .Q(d1[1]) );
  DFF_EN d1_reg_0_ ( .D(upstream_data[0]), .E(N29), .CP(clk), .Q(d1[0]) );
  DFF_EN d1_reg_2_ ( .D(upstream_data[2]), .E(N29), .CP(clk), .Q(d1[2]) );
  DFF_EN d1_reg_4_ ( .D(upstream_data[4]), .E(N29), .CP(clk), .Q(d1[4]) );
  DFF_EN d1_reg_6_ ( .D(upstream_data[6]), .E(N29), .CP(clk), .Q(d1[6]) );
  DFF d0_reg_7_ ( .D(n8), .CP(clk), .Q(downstream_data[7]) );
  DFF d0_reg_5_ ( .D(n10), .CP(clk), .Q(downstream_data[5]) );
  DFF d0_reg_3_ ( .D(n12), .CP(clk), .Q(downstream_data[3]) );
  DFF d0_reg_1_ ( .D(n14), .CP(clk), .Q(downstream_data[1]) );
  DFF d0_reg_0_ ( .D(n15), .CP(clk), .Q(downstream_data[0]) );
  DFF d0_reg_2_ ( .D(n13), .CP(clk), .Q(downstream_data[2]) );
  DFF d0_reg_4_ ( .D(n11), .CP(clk), .Q(downstream_data[4]) );
  DFF d0_reg_6_ ( .D(n9), .CP(clk), .Q(downstream_data[6]) );
  DFF_EN ready_reg_reg ( .D(N3), .E(reset_n), .CP(clk), .Q(ready_reg) );
  DFF_EN_RST v1_reg (.D(upstream_rdy), .E(upstream_acpt), .CP(clk), .CDN(reset_n), .Q(v1));
  INV U2 ( .I(reset_n), .ZN(n1) );
  NOR2 U3 ( .A1(n6), .A2(upstream_acpt), .ZN(n4) );
  I_NAND3 U4 ( .A1(upstream_rdy), .B1(upstream_acpt), .B2(N3), .ZN(n16) );
  INV U5 ( .I(n7), .ZN(upstream_acpt) );
  NOR2 U6 ( .A1(n6), .A2(n7), .ZN(n5) );
  NAND2 U7 ( .A1(N3), .A2(reset_n), .ZN(n6) );
  NOR2 U8 ( .A1(n7), .A2(n1), .ZN(N29) );
  AO222 U9 ( .A1(d1[6]), .A2(n4), .B1(upstream_data[6]), .B2(n5), .C1(downstream_data[6]), .C2(n6), .Z(n9) );
  AO222 U10 ( .A1(d1[4]), .A2(n4), .B1(upstream_data[4]), .B2(n5), .C1(downstream_data[4]), .C2(n6), .Z(n11) );
  AO222 U11 ( .A1(d1[2]), .A2(n4), .B1(upstream_data[2]), .B2(n5), .C1(downstream_data[2]), .C2(n6), .Z(n13) );
  AO222 U12 ( .A1(d1[0]), .A2(n4), .B1(upstream_data[0]), .B2(n5), .C1(downstream_data[0]), .C2(n6), .Z(n15) );
  AO222 U13 ( .A1(d1[1]), .A2(n4), .B1(upstream_data[1]), .B2(n5), .C1(downstream_data[1]), .C2(n6), .Z(n14) );
  AO222 U14 ( .A1(d1[3]), .A2(n4), .B1(upstream_data[3]), .B2(n5), .C1(downstream_data[3]), .C2(n6), .Z(n12) );
  AO222 U15 ( .A1(d1[5]), .A2(n4), .B1(upstream_data[5]), .B2(n5), .C1(downstream_data[5]), .C2(n6), .Z(n10) );
  AO222 U16 ( .A1(d1[7]), .A2(n4), .B1(upstream_data[7]), .B2(n5), .C1(downstream_data[7]), .C2(n6), .Z(n8) );
  I_NOR2 U17 ( .A1(v1), .B1(ready_reg), .ZN(n7) );
  I_NAND2 U18 ( .A1(downstream_acpt), .B1(downstream_rdy), .ZN(N3) );
endmodule


module mem_ctrl ( clk, rstn, do_rdy, mc_pwr, memsel, mc_save, mc_restore, 
        mc_pwr_ack, do_acpt, ceb, web, addr );
  input [1:0] memsel;
  output [3:0] ceb;
  output [3:0] web;
  output [7:0] addr;
  input clk, rstn, do_rdy, mc_pwr, mc_save, mc_restore;
  output mc_pwr_ack, do_acpt;
  wire   n66, n67, n68, N8, N9, N10, N11, N12, N13, N14, N15, n3, n9, n10, n11,
         n14, n28, n31, n34, n37, n40, n43, n46, n49, n6, n7, n8, n12, n13,
         n15, n16, n17, n18, n19, n52, n53, n54, n55, n56, n57, n58, n59, n60;
  wire   [69:70] n;
  wire   [3:0] next_state;
  wire   [3:0] present_state;

  DFF_RET present_state_reg_1_ ( .SAVE(mc_save), .NRESTORE(mc_restore), 
        .D(next_state[1]), .SI(1'b0), .SE(1'b0), .CP(n66), .CDN(n67), .SDN(
        1'b1), .Q(present_state[1]) ); //synopsys retention_upf mem_ctrl_ret+PD_mem_ctrl
  DFF_RET present_state_reg_2_ ( .SAVE(mc_save), .NRESTORE(mc_restore), 
        .D(next_state[2]), .SI(1'b0), .SE(1'b0), .CP(n66), .CDN(n67), .SDN(
        1'b1), .Q(present_state[2]) ); //synopsys retention_upf mem_ctrl_ret+PD_mem_ctrl
  mem_ctrl_DW01_inc_0 add_34 ( .A(addr), .SUM({N15, N14, N13, N12, N11, N10, 
        N9, N8}) );
  DFF_RET present_state_reg_0_ ( .SAVE(mc_save), .NRESTORE(mc_restore), 
        .D(next_state[0]), .SI(1'b0), .SE(1'b0), .CP(n66), .CDN(n67), .SDN(
        1'b1), .Q(present_state[0]) ); //synopsys retention_upf mem_ctrl_ret+PD_mem_ctrl
  DFF_RET addr_reg_7_ ( .SAVE(mc_save), .NRESTORE(mc_restore), .D(n49), 
        .SI(1'b0), .SE(1'b0), .CP(n66), .CDN(n67), .SDN(1'b1), .Q(addr[7]) ); //synopsys retention_upf mem_ctrl_ret+PD_mem_ctrl
  DFF_RET addr_reg_6_ ( .SAVE(mc_save), .NRESTORE(mc_restore), .D(n28), 
        .SI(1'b0), .SE(1'b0), .CP(n66), .CDN(n67), .SDN(1'b1), .Q(addr[6]) ); //synopsys retention_upf mem_ctrl_ret+PD_mem_ctrl
  DFF_RET addr_reg_4_ ( .SAVE(mc_save), .NRESTORE(mc_restore), .D(n34), 
        .SI(1'b0), .SE(1'b0), .CP(n66), .CDN(n67), .SDN(1'b1), .Q(addr[4]) ); //synopsys retention_upf mem_ctrl_ret+PD_mem_ctrl
  DFF_RET addr_reg_3_ ( .SAVE(mc_save), .NRESTORE(mc_restore), .D(n37), 
        .SI(1'b0), .SE(1'b0), .CP(n66), .CDN(n67), .SDN(1'b1), .Q(addr[3]) ); //synopsys retention_upf mem_ctrl_ret+PD_mem_ctrl
  DFF_RET addr_reg_5_ ( .SAVE(mc_save), .NRESTORE(mc_restore), .D(n31), 
        .SI(1'b0), .SE(1'b0), .CP(n66), .CDN(n67), .SDN(1'b1), .Q(addr[5]) ); //synopsys retention_upf mem_ctrl_ret+PD_mem_ctrl
  DFF_RET addr_reg_2_ ( .SAVE(mc_save), .NRESTORE(mc_restore), .D(n40), 
        .SI(1'b0), .SE(1'b0), .CP(n66), .CDN(n67), .SDN(1'b1), .Q(addr[2]) ); //synopsys retention_upf mem_ctrl_ret+PD_mem_ctrl
  DFF_RET addr_reg_1_ ( .SAVE(mc_save), .NRESTORE(mc_restore), .D(n43), 
        .SI(1'b0), .SE(1'b0), .CP(n66), .CDN(n67), .SDN(1'b1), .Q(addr[1]) ); //synopsys retention_upf mem_ctrl_ret+PD_mem_ctrl
  DFF_RET addr_reg_0_ ( .SAVE(mc_save), .NRESTORE(mc_restore), .D(n46), 
        .SI(1'b0), .SE(1'b0), .CP(n66), .CDN(n67), .SDN(1'b1), .Q(addr[0]) ); //synopsys retention_upf mem_ctrl_ret+PD_mem_ctrl
  DFF_RET present_state_reg_3_ ( .SAVE(mc_save), .NRESTORE(mc_restore), 
        .D(next_state[3]), .SI(1'b0), .SE(1'b0), .CP(n66), .CDN(n67), .SDN(
        1'b1), .Q(present_state[3]) ); //synopsys retention_upf mem_ctrl_ret+PD_mem_ctrl
  LS_HL LS_clk_UPF_LS ( .I(clk), .Z(n66) );
  OR2 U3 ( .A1(ceb[3]), .A2(present_state[2]), .Z(web[3]) );
  AO211 U9 ( .A1(n59), .A2(present_state[0]), .B(n57), .C(n56), .Z(
        next_state[1]) );
  AO211 U8 ( .A1(n56), .A2(present_state[2]), .B(n57), .C(do_acpt), .Z(
        next_state[2]) );
  LS_HL LS_do_rdy_UPF_LS ( .I(do_rdy), .Z(n68) );
  AOI22 U11 ( .A1(n68), .A2(n58), .B1(present_state[1]), .B2(n60), .ZN(n11) );
  AOI31 U10 ( .A1(n9), .A2(n10), .A3(n11), .B(present_state[0]), .ZN(
        next_state[0]) );
  NAND2 U21 ( .A1(n58), .A2(present_state[0]), .ZN(n14) );
  LS_HL LS_memsel_0__UPF_LS ( .I(memsel[0]), .Z(n[70]) );
  LS_HL LS_memsel_1__UPF_LS ( .I(memsel[1]), .Z(n[69]) );
  LS_HL LS_rstn_UPF_LS ( .I(rstn), .Z(n67) );
  I_NOR2 U7 ( .A1(n55), .B1(present_state[2]), .ZN(n3) );
  INV U4 ( .I(1'b1), .ZN(mc_pwr_ack) );
  I_NAND2 U6 ( .A1(n60), .B1(n59), .ZN(n10) );
  I_NAND3 U12 ( .A1(n9), .B1(present_state[0]), .B2(n7), .ZN(n52) );
  I_NAND3 U13 ( .A1(n[70]), .B1(n55), .B2(n54), .ZN(ceb[0]) );
  NOR2 U14 ( .A1(n9), .A2(present_state[1]), .ZN(n16) );
  NOR2 U15 ( .A1(n13), .A2(present_state[2]), .ZN(n15) );
  OAI21 U16 ( .A1(n17), .A2(n9), .B(n10), .ZN(next_state[3]) );
  I_NAND3 U17 ( .A1(n[69]), .B1(n53), .B2(n3), .ZN(web[0]) );
  I_NAND3 U18 ( .A1(n[70]), .B1(n[69]), .B2(n3), .ZN(web[2]) );
  I_NAND3 U19 ( .A1(n[69]), .B1(n[70]), .B2(n3), .ZN(web[1]) );
  I_NAND3 U20 ( .A1(n[70]), .B1(n55), .B2(n[69]), .ZN(ceb[2]) );
  I_NAND3 U22 ( .A1(n[69]), .B1(n55), .B2(n[70]), .ZN(ceb[1]) );
  NAND3 U23 ( .A1(n[70]), .A2(n[69]), .A3(n56), .ZN(ceb[3]) );
  I_NAND2 U24 ( .A1(next_state[3]), .B1(n18), .ZN(n19) );
  I_NAND2 U25 ( .A1(present_state[3]), .B1(present_state[2]), .ZN(n9) );
  NAND2 U26 ( .A1(present_state[0]), .A2(present_state[1]), .ZN(n17) );
  I_NAND2 U27 ( .A1(present_state[3]), .B1(present_state[1]), .ZN(n13) );
  OR2 U28 ( .A1(present_state[2]), .A2(present_state[1]), .Z(n18) );
  I_NAND2 U29 ( .A1(present_state[0]), .B1(n8), .ZN(n12) );
  I_NAND2 U30 ( .A1(present_state[3]), .B1(n59), .ZN(n6) );
  INV U31 ( .I(n18), .ZN(n59) );
  INV U32 ( .I(n6), .ZN(n58) );
  INV U33 ( .I(present_state[3]), .ZN(n60) );
  INV U34 ( .I(present_state[1]), .ZN(n7) );
  INV U35 ( .I(n52), .ZN(n57) );
  INV U36 ( .I(n13), .ZN(n8) );
  INV U37 ( .I(n12), .ZN(n56) );
  MUX21 U38 ( .I0(n16), .I1(n15), .S(present_state[0]), .Z(do_acpt) );
  I_NOR4 U39 ( .A1(n52), .B1(do_acpt), .B2(present_state[3]), .B3(n19), .ZN(n55) );
  INV U40 ( .I(n[70]), .ZN(n53) );
  INV U41 ( .I(n[69]), .ZN(n54) );
  MUX21 U66 ( .I0(N14), .I1(addr[6]), .S(n14), .Z(n28) );
  MUX21 U67 ( .I0(N13), .I1(addr[5]), .S(n14), .Z(n31) );
  MUX21 U68 ( .I0(N12), .I1(addr[4]), .S(n14), .Z(n34) );
  MUX21 U69 ( .I0(N11), .I1(addr[3]), .S(n14), .Z(n37) );
  MUX21 U70 ( .I0(N10), .I1(addr[2]), .S(n14), .Z(n40) );
  MUX21 U71 ( .I0(N9), .I1(addr[1]), .S(n14), .Z(n43) );
  MUX21 U72 ( .I0(N8), .I1(addr[0]), .S(n14), .Z(n46) );
  MUX21 U73 ( .I0(N15), .I1(addr[7]), .S(n14), .Z(n49) );
endmodule


module async_bridge ( clk1, clk2, rstn, do_rdy_in, do_acpt_in, do_acpt_out, 
        do_rdy_out );
  input clk1, clk2, rstn, do_rdy_in, do_acpt_in;
  output do_acpt_out, do_rdy_out;
  wire   do_rdy_in_d2, do_rdy_in_d1, do_rdy, N3, do_acpt, ready_tmp, acpt_tmp1,
         acpt_tmp3, acpt_tmp2, n2;

  DFF_RST do_rdy_in_d2_reg ( .D(do_rdy_in_d1), .CP(clk1), .CDN(rstn), .Q(
        do_rdy_in_d2) );
  DFF_RST do_rdy_out_reg ( .D(ready_tmp), .CP(clk2), .CDN(rstn), .Q(
        do_rdy_out) );
  DFF_RST do_rdy_in_d1_reg ( .D(do_rdy_in), .CP(clk1), .CDN(rstn), .Q(
        do_rdy_in_d1) );
  DFF_RST acpt_tmp2_reg ( .D(acpt_tmp1), .CP(clk1), .CDN(rstn), .Q(
        acpt_tmp2) );
  DFF_RST acpt_tmp3_reg ( .D(acpt_tmp2), .CP(clk1), .CDN(rstn), .Q(
        acpt_tmp3) );
  DFF_RST do_rdy_reg ( .D(N3), .CP(clk1), .CDN(rstn), .Q(do_rdy) );
  DFF_RST do_acpt_reg ( .D(do_acpt_in), .CP(clk2), .CDN(rstn), .Q(do_acpt)
         );
  DFF_RST ready_tmp_reg ( .D(do_rdy), .CP(clk2), .CDN(rstn), .Q(ready_tmp)
         );
  DFF_RST acpt_tmp1_reg ( .D(do_acpt), .CP(clk1), .CDN(rstn), .Q(acpt_tmp1)
         );
  I_NOR2 U3 ( .A1(acpt_tmp2), .B1(acpt_tmp3), .ZN(do_acpt_out) );
  MOAI22 U4 ( .A1(do_rdy_in_d2), .A2(n2), .B1(do_rdy_in), .B2(
        do_rdy_in_d1), .ZN(N3) );
  NOR2 U5 ( .A1(do_rdy_in), .A2(do_rdy_in_d1), .ZN(n2) );
endmodule


module interleaver ( clk, reset_n, di_rdy, do_acpt, enable, di_data, do_rdy, 
        di_acpt, do_data );
  input [7:0] di_data;
  output [7:0] do_data;
  input clk, reset_n, di_rdy, do_acpt, enable;
  output do_rdy, di_acpt;
  wire   n93, n94, n95, n96, n97, in_acpt, in_rdy, out_acpt, out_rdy, pkt_zero,
         pkt_cen, N56, N57, N58, N59, N60, N61, N62, N63, N531, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75,
         n76, n77, n78, n79, n1, n2, n16, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92;
  wire   [98:105] n;
  wire   [4:0] int_state;
  wire   [3:0] data_sel;
  wire   [10:0] push;
  wire   [7:0] do_reg;
  wire   [7:0] input_down_data;
  wire   [7:0] fifo_data;
  wire   [4:0] nxt_state;

  DFF_RST int_state_reg_0_ ( .D(nxt_state[0]), .CP(n93), .CDN(n1), .Q(int_state[0]) );
  DFF_RST int_state_reg_1_ ( .D(nxt_state[1]), .CP(n93), .CDN(n1), .Q(int_state[1]) );
  DFF_RST int_state_reg_4_ ( .D(nxt_state[4]), .CP(n93), .CDN(n1), .Q(int_state[4]) );
  DFF_RST int_state_reg_2_ ( .D(nxt_state[2]), .CP(n93), .CDN(n1), .Q(int_state[2]) );
  rdyacpt_WIDTH8_0 in2wire ( .clk(n93), .reset_n(n1), .upstream_rdy(n95), 
        .downstream_acpt(in_acpt), .upstream_data(n), .downstream_rdy(in_rdy), 
        .upstream_acpt(di_acpt), .downstream_data(input_down_data) );
  count_WIDTH8 pkt_counter ( .clk(n93), .rst_n(n1), .ld_n(N531), .up_dn(1'b0), 
        .cen(pkt_cen), .din({1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b0, 1'b1, 1'b1}), 
        .zero(pkt_zero) );
  fifo_shift_ram fifo ( .clk(n93), .reset_n(n1), .ram_re(n16), .push({
        push[10:1], n80}), .din(input_down_data), .sel(data_sel), .dout(
        fifo_data) );
  rdyacpt_WIDTH8_1 out2wire ( .clk(n93), .reset_n(n1), .upstream_rdy(out_rdy), 
        .downstream_acpt(n96), .upstream_data(do_reg), .downstream_rdy(do_rdy), 
        .upstream_acpt(out_acpt), .downstream_data(do_data) );
  LS_HL LS_clk_UPF_LS ( .I(clk), .Z(n93) );
  DFF do_reg_reg_0_ ( .D(N56), .CP(n93), .Q(do_reg[0]) );
  DFF do_reg_reg_7_ ( .D(N63), .CP(n93), .Q(do_reg[7]) );
  DFF do_reg_reg_6_ ( .D(N62), .CP(n93), .Q(do_reg[6]) );
  DFF do_reg_reg_5_ ( .D(N61), .CP(n93), .Q(do_reg[5]) );
  DFF do_reg_reg_4_ ( .D(N60), .CP(n93), .Q(do_reg[4]) );
  DFF do_reg_reg_3_ ( .D(N59), .CP(n93), .Q(do_reg[3]) );
  DFF do_reg_reg_2_ ( .D(N58), .CP(n93), .Q(do_reg[2]) );
  DFF do_reg_reg_1_ ( .D(N57), .CP(n93), .Q(do_reg[1]) );
  DFF_RST int_state_reg_3_ ( .D(nxt_state[3]), .CP(n93), .CDN(n1), .Q(int_state[3]) );
  LS_HL LS_do_acpt_UPF_LS ( .I(do_acpt), .Z(n96) );
  LS_HL LS_enable_UPF_LS ( .I(enable), .Z(n97) );
  LS_HL LS_reset_n_UPF_LS ( .I(reset_n), .Z(n94) );
  LS_HL LS_di_rdy_UPF_LS ( .I(di_rdy), .Z(n95) );
  LS_HL LS_di_data_7__UPF_LS ( .I(di_data[7]), .Z(n[98]) );
  LS_HL LS_di_data_5__UPF_LS ( .I(di_data[5]), .Z(n[100]) );
  LS_HL LS_di_data_3__UPF_LS ( .I(di_data[3]), .Z(n[102]) );
  LS_HL LS_di_data_1__UPF_LS ( .I(di_data[1]), .Z(n[104]) );
  LS_HL LS_di_data_0__UPF_LS ( .I(di_data[0]), .Z(n[105]) );
  LS_HL LS_di_data_2__UPF_LS ( .I(di_data[2]), .Z(n[103]) );
  LS_HL LS_di_data_4__UPF_LS ( .I(di_data[4]), .Z(n[101]) );
  LS_HL LS_di_data_6__UPF_LS ( .I(di_data[6]), .Z(n[99]) );
  I_NAND4 U3 ( .A1(n52), .B1(n53), .B2(n50), .B3(n54), .ZN(data_sel[3]) );
  NAND4 U4 ( .A1(n84), .A2(n43), .A3(n57), .A4(n85), .ZN(data_sel[2]) );
  INV U5 ( .I(n2), .ZN(n1) );
  NAND2 U6 ( .A1(in_rdy), .A2(in_acpt), .ZN(n18) );
  I_NOR2 U7 ( .A1(n35), .B1(n82), .ZN(n57) );
  I_NAND4 U8 ( .A1(n41), .B1(n87), .B2(n43), .B3(n85), .ZN(data_sel[1]) );
  NAND2 U9 ( .A1(n28), .A2(n60), .ZN(n20) );
  NAND2 U10 ( .A1(n20), .A2(n69), .ZN(n24) );
  AND2 U11 ( .A1(n48), .A2(n59), .Z(n43) );
  NAND2 U12 ( .A1(n40), .A2(n70), .ZN(n32) );
  NAND2 U13 ( .A1(n39), .A2(n66), .ZN(n52) );
  AND2 U14 ( .A1(n47), .A2(n62), .Z(n53) );
  NOR2 U15 ( .A1(n71), .A2(n72), .ZN(n51) );
  I_NAND4 U16 ( .A1(push[10]), .B1(n17), .B2(n73), .B3(n74), .ZN(n71) );
  NOR3 U17 ( .A1(push[1]), .A2(push[3]), .A3(push[2]), .ZN(n73) );
  NOR4 U18 ( .A1(n75), .A2(push[4]), .A3(push[6]), .A4(push[5]), .ZN(n74));
  OR3 U19 ( .A1(push[8]), .A2(push[9]), .A3(push[7]), .Z(n75) );
  NAND2 U20 ( .A1(out_acpt), .A2(out_rdy), .ZN(n21) );
  AND2 U21 ( .A1(n28), .A2(n29), .Z(n25) );
  NAND4 U22 ( .A1(n84), .A2(n85), .A3(n87), .A4(n64), .ZN(data_sel[0]) );
  I_NOR3 U23 ( .A1(n38), .B1(n52), .B2(n65), .ZN(n64) );
  NOR2 U24 ( .A1(n88), .A2(n86), .ZN(n28) );
  I_NOR2 U25 ( .A1(n78), .B1(n92), .ZN(n60) );
  I_NOR2 U26 ( .A1(n79), .B1(n92), .ZN(n29) );
  NAND3 U27 ( .A1(n46), .A2(n61), .A3(n53), .ZN(n41) );
  NAND2 U28 ( .A1(n29), .A2(n76), .ZN(n66) );
  NAND2 U29 ( .A1(n60), .A2(n76), .ZN(n70) );
  NAND2 U30 ( .A1(n55), .A2(n58), .ZN(n34) );
  NAND2 U31 ( .A1(n77), .A2(n29), .ZN(n62) );
  NAND2 U32 ( .A1(n55), .A2(n60), .ZN(n48) );
  NAND2 U33 ( .A1(n55), .A2(n29), .ZN(n47) );
  NAND2 U34 ( .A1(n60), .A2(n77), .ZN(n59) );
  NAND2 U35 ( .A1(n28), .A2(n56), .ZN(n39) );
  AND2 U36 ( .A1(n63), .A2(n76), .Z(n65) );
  NAND2 U37 ( .A1(n55), .A2(n63), .ZN(n46) );
  NAND2 U38 ( .A1(n58), .A2(n77), .ZN(n35) );
  NAND2 U39 ( .A1(n27), .A2(n68), .ZN(n33) );
  NAND2 U40 ( .A1(n77), .A2(n56), .ZN(n54) );
  NAND2 U41 ( .A1(n56), .A2(n76), .ZN(n69) );
  NAND2 U42 ( .A1(n58), .A2(n76), .ZN(n68) );
  NAND2 U43 ( .A1(n55), .A2(n56), .ZN(n50) );
  NAND2 U44 ( .A1(n28), .A2(n58), .ZN(n40) );
  NAND3 U45 ( .A1(n81), .A2(n92), .A3(n67), .ZN(n17) );
  NOR2 U46 ( .A1(n61), .A2(n18), .ZN(push[2]) );
  NOR2 U47 ( .A1(n70), .A2(n18), .ZN(push[5]) );
  NOR2 U48 ( .A1(n18), .A2(n66), .ZN(push[9]) );
  NOR2 U49 ( .A1(n59), .A2(n18), .ZN(push[6]) );
  NOR2 U50 ( .A1(n35), .A2(n18), .ZN(push[4]) );
  NOR2 U51 ( .A1(n68), .A2(n18), .ZN(push[3]) );
  I_NOR2 U52 ( .A1(n65), .B1(n18), .ZN(push[1]) );
  NOR2 U53 ( .A1(n54), .A2(n18), .ZN(push[8]) );
  NOR2 U54 ( .A1(n69), .A2(n18), .ZN(push[7]) );
  OAI21 U55 ( .A1(n16), .A2(n86), .B(n51), .ZN(nxt_state[0]) );
  NOR2 U56 ( .A1(n62), .A2(n18), .ZN(push[10]) );
  AOI21 U57 ( .A1(n42), .A2(N531), .B(n18), .ZN(n72) );
  NAND2 U58 ( .A1(n49), .A2(n86), .ZN(N531) );
  OAI221 U59 ( .A1(n16), .A2(n20), .B1(n81), .B2(n42), .C(n43), .ZN(n30));
  I_NAND3 U60 ( .A1(pkt_zero), .B1(n25), .B2(n16), .ZN(n22) );
  NOR3 U61 ( .A1(n18), .A2(pkt_zero), .A3(n2), .ZN(pkt_cen) );
  NOR2 U62 ( .A1(n86), .A2(n90), .ZN(out_rdy) );
  OAI221 U63 ( .A1(n26), .A2(n89), .B1(n27), .B2(n21), .C(n22), .ZN(nxt_state[3]) );
  NOR4 U64 ( .A1(n30), .A2(n31), .A3(n32), .A4(n33), .ZN(n26) );
  NAND2 U65 ( .A1(n34), .A2(n35), .ZN(n31) );
  OAI221 U66 ( .A1(n19), .A2(n91), .B1(n20), .B2(n21), .C(n22), .ZN(nxt_state[4]) );
  AOI211 U67 ( .A1(n90), .A2(n18), .B(n23), .C(n24), .ZN(n19) );
  AO21 U68 ( .A1(n21), .A2(n25), .B(data_sel[3]), .Z(n23) );
  INV U69 ( .I(n94), .ZN(n2) );
  NOR2 U70 ( .A1(n86), .A2(int_state[1]), .ZN(n55) );
  NOR3 U71 ( .A1(int_state[3]), .A2(int_state[4]), .A3(n88), .ZN(n67) );
  NAND3 U72 ( .A1(int_state[2]), .A2(n86), .A3(n67), .ZN(n61) );
  NAND3 U73 ( .A1(int_state[2]), .A2(int_state[0]), .A3(n67), .ZN(n27) );
  NAND3 U74 ( .A1(int_state[0]), .A2(n92), .A3(n67), .ZN(n38) );
  NOR2 U75 ( .A1(int_state[1]), .A2(int_state[0]), .ZN(n76) );
  I_NOR2 U76 ( .A1(n79), .B1(int_state[2]), .ZN(n56) );
  I_NOR2 U77 ( .A1(n78), .B1(int_state[2]), .ZN(n58) );
  NOR2 U78 ( .A1(n88), .A2(int_state[0]), .ZN(n77) );
  NOR2 U79 ( .A1(n91), .A2(int_state[3]), .ZN(n79) );
  INV U80 ( .I(int_state[3]), .ZN(n89) );
  NOR2 U81 ( .A1(n89), .A2(int_state[4]), .ZN(n78) );
  MOAI22 U82 ( .A1(int_state[0]), .A2(n90), .B1(n92), .B2(n76), .ZN(in_acpt) );
  AO222 U83 ( .A1(fifo_data[1]), .A2(n71), .B1(do_reg[1]), .B2(n51), .C1(input_down_data[1]), .C2(n72), .Z(N57) );
  AO222 U84 ( .A1(fifo_data[2]), .A2(n71), .B1(do_reg[2]), .B2(n51), .C1(input_down_data[2]), .C2(n72), .Z(N58) );
  AO222 U85 ( .A1(fifo_data[3]), .A2(n71), .B1(do_reg[3]), .B2(n51), .C1(input_down_data[3]), .C2(n72), .Z(N59) );
  AO222 U86 ( .A1(fifo_data[4]), .A2(n71), .B1(do_reg[4]), .B2(n51), .C1(input_down_data[4]), .C2(n72), .Z(N60) );
  AO222 U87 ( .A1(fifo_data[5]), .A2(n71), .B1(do_reg[5]), .B2(n51), .C1(input_down_data[5]), .C2(n72), .Z(N61) );
  AO222 U88 ( .A1(fifo_data[6]), .A2(n71), .B1(do_reg[6]), .B2(n51), .C1(input_down_data[6]), .C2(n72), .Z(N62) );
  AO222 U89 ( .A1(fifo_data[7]), .A2(n71), .B1(do_reg[7]), .B2(n51), .C1(input_down_data[7]), .C2(n72), .Z(N63) );
  AO222 U90 ( .A1(fifo_data[0]), .A2(n71), .B1(do_reg[0]), .B2(n51), .C1(input_down_data[0]), .C2(n72), .Z(N56) );
  NAND2 U91 ( .A1(n36), .A2(n37), .ZN(nxt_state[2]) );
  AO31 U92 ( .A1(n38), .A2(n39), .A3(n40), .B(n21), .Z(n37) );
  OAI31 U93 ( .A1(n41), .A2(n21), .A3(n30), .B(int_state[2]), .ZN(n36) );
  OAI221 U94 ( .A1(n16), .A2(n88), .B1(n21), .B2(n44), .C(n45), .ZN(nxt_state[1]) );
  AOI211 U95 ( .A1(n97), .A2(n49), .B(n83), .C(n82), .ZN(n44) );
  AO31 U96 ( .A1(n46), .A2(n47), .A3(n48), .B(n21), .Z(n45) );
  NOR4 U97 ( .A1(int_state[1]), .A2(int_state[2]), .A3(int_state[3]), .A4(int_state[4]), .ZN(n49) );
  NAND2 U98 ( .A1(int_state[4]), .A2(int_state[3]), .ZN(n42) );
  NOR3 U99 ( .A1(int_state[3]), .A2(int_state[4]), .A3(n92), .ZN(n63) );
  INV U100 ( .I(n21), .ZN(n16) );
  INV U101 ( .I(n17), .ZN(n80) );
  INV U102 ( .I(n18), .ZN(n81) );
  INV U103 ( .I(n34), .ZN(n82) );
  INV U104 ( .I(n50), .ZN(n83) );
  INV U105 ( .I(n32), .ZN(n84) );
  INV U106 ( .I(n24), .ZN(n85) );
  INV U107 ( .I(int_state[0]), .ZN(n86) );
  INV U108 ( .I(n33), .ZN(n87) );
  INV U109 ( .I(int_state[1]), .ZN(n88) );
  INV U110 ( .I(n42), .ZN(n90) );
  INV U111 ( .I(int_state[4]), .ZN(n91) );
  INV U112 ( .I(int_state[2]), .ZN(n92) );
endmodule


module design_top ( clk1, clk2, reset_n, di_rdy, mc_pwr, mc_save, mc_restore, 
        mc_iso, mc_clk_gate, sram_pwr, memsel, di_data, di_acpt, mc_pwr_ack, 
        q1, q2, q3, q4 );
  input [1:0] memsel;
  input [7:0] di_data;
  output [15:0] q1;
  output [15:0] q2;
  output [15:0] q3;
  output [15:0] q4;
  input clk1, clk2, reset_n, di_rdy, mc_pwr, mc_save, mc_restore, mc_iso,
         mc_clk_gate, sram_pwr;
  output di_acpt, mc_pwr_ack;
  wire   clk1_c, clk2_c, reset_n_c, di_rdy_c, mc_pwr_c, mc_save_c,
         mc_restore_c, mc_clk_gate_c, sram_pwr_c, di_acpt_i, do_acpt_out,
         do_rdy, do_acpt, do_rdy_out, clk2_gate, n2, n3, n4, n5, n6, n7, n8,
         n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22,
         n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36,
         n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50,
         n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175;
  wire   [1:0] memsel_c;
  wire   [7:0] di_data_c;
  wire   [15:0] q1_i;
  wire   [15:0] q2_i;
  wire   [15:0] q3_i;
  wire   [15:0] q4_i;
  wire   [7:0] do_data;
  wire   [3:0] ceb;
  wire   [3:0] web;
  wire   [7:0] address;

  PAD_IN pi0 ( .PAD(clk1), .C(clk1_c) );
  PAD_IN pi1 ( .PAD(clk2), .C(clk2_c) );
  PAD_IN pi2 ( .PAD(reset_n), .C(reset_n_c) );
  PAD_IN pi3 ( .PAD(di_rdy), .C(di_rdy_c) );
  PAD_IN pi4 ( .PAD(mc_pwr), .C(mc_pwr_c) );
  PAD_IN pi5 ( .PAD(mc_save), .C(mc_save_c) );
  PAD_IN pi6 ( .PAD(mc_restore), .C(mc_restore_c) );
  PAD_IN pi7 ( .PAD(mc_iso), .C(n174) );
  PAD_IN pi8 ( .PAD(mc_clk_gate), .C(mc_clk_gate_c) );
  PAD_IN pi9 ( .PAD(sram_pwr), .C(sram_pwr_c) );
  PAD_IN pi_10 ( .PAD(memsel[0]), .C(memsel_c[0]) );
  PAD_IN pi_11 ( .PAD(memsel[1]), .C(memsel_c[1]) );
  PAD_IN di_data_slice_0__pi_12 ( .PAD(di_data[0]), .C(di_data_c[0]) );
  PAD_IN di_data_slice_1__pi_12 ( .PAD(di_data[1]), .C(di_data_c[1]) );
  PAD_IN di_data_slice_2__pi_12 ( .PAD(di_data[2]), .C(di_data_c[2]) );
  PAD_IN di_data_slice_3__pi_12 ( .PAD(di_data[3]), .C(di_data_c[3]) );
  PAD_IN di_data_slice_4__pi_12 ( .PAD(di_data[4]), .C(di_data_c[4]) );
  PAD_IN di_data_slice_5__pi_12 ( .PAD(di_data[5]), .C(di_data_c[5]) );
  PAD_IN di_data_slice_6__pi_12 ( .PAD(di_data[6]), .C(di_data_c[6]) );
  PAD_IN di_data_slice_7__pi_12 ( .PAD(di_data[7]), .C(di_data_c[7]) );
  PAD_OUT po0 ( .I(di_acpt_i), .PAD(di_acpt) );
  PAD_OUT po1 ( .I(1'b0), .PAD(mc_pwr_ack) );
  PAD_OUT q1_slice_0__po2 ( .I(n99), .PAD(q1[0]) );
  PAD_OUT q1_slice_1__po2 ( .I(n101), .PAD(q1[1]) );
  PAD_OUT q1_slice_2__po2 ( .I(n103), .PAD(q1[2]) );
  PAD_OUT q1_slice_3__po2 ( .I(n105), .PAD(q1[3]) );
  PAD_OUT q1_slice_4__po2 ( .I(n107), .PAD(q1[4]) );
  PAD_OUT q1_slice_5__po2 ( .I(n109), .PAD(q1[5]) );
  PAD_OUT q1_slice_6__po2 ( .I(n111), .PAD(q1[6]) );
  PAD_OUT q1_slice_7__po2 ( .I(n113), .PAD(q1[7]) );
  PAD_OUT q1_slice_8__po2 ( .I(n115), .PAD(q1[8]) );
  PAD_OUT q1_slice_9__po2 ( .I(n117), .PAD(q1[9]) );
  PAD_OUT q1_slice_10__po2 ( .I(n119), .PAD(q1[10]) );
  PAD_OUT q1_slice_11__po2 ( .I(n121), .PAD(q1[11]) );
  PAD_OUT q1_slice_12__po2 ( .I(n123), .PAD(q1[12]) );
  PAD_OUT q1_slice_13__po2 ( .I(n125), .PAD(q1[13]) );
  PAD_OUT q1_slice_14__po2 ( .I(n127), .PAD(q1[14]) );
  PAD_OUT q1_slice_15__po2 ( .I(n129), .PAD(q1[15]) );
  PAD_OUT q2_slice_0__po3 ( .I(n67), .PAD(q2[0]) );
  PAD_OUT q2_slice_1__po3 ( .I(n69), .PAD(q2[1]) );
  PAD_OUT q2_slice_2__po3 ( .I(n71), .PAD(q2[2]) );
  PAD_OUT q2_slice_3__po3 ( .I(n73), .PAD(q2[3]) );
  PAD_OUT q2_slice_4__po3 ( .I(n75), .PAD(q2[4]) );
  PAD_OUT q2_slice_5__po3 ( .I(n77), .PAD(q2[5]) );
  PAD_OUT q2_slice_6__po3 ( .I(n79), .PAD(q2[6]) );
  PAD_OUT q2_slice_7__po3 ( .I(n81), .PAD(q2[7]) );
  PAD_OUT q2_slice_8__po3 ( .I(n83), .PAD(q2[8]) );
  PAD_OUT q2_slice_9__po3 ( .I(n85), .PAD(q2[9]) );
  PAD_OUT q2_slice_10__po3 ( .I(n87), .PAD(q2[10]) );
  PAD_OUT q2_slice_11__po3 ( .I(n89), .PAD(q2[11]) );
  PAD_OUT q2_slice_12__po3 ( .I(n91), .PAD(q2[12]) );
  PAD_OUT q2_slice_13__po3 ( .I(n93), .PAD(q2[13]) );
  PAD_OUT q2_slice_14__po3 ( .I(n95), .PAD(q2[14]) );
  PAD_OUT q2_slice_15__po3 ( .I(n97), .PAD(q2[15]) );
  PAD_OUT q3_slice_0__po4 ( .I(n35), .PAD(q3[0]) );
  PAD_OUT q3_slice_1__po4 ( .I(n37), .PAD(q3[1]) );
  PAD_OUT q3_slice_2__po4 ( .I(n39), .PAD(q3[2]) );
  PAD_OUT q3_slice_3__po4 ( .I(n41), .PAD(q3[3]) );
  PAD_OUT q3_slice_4__po4 ( .I(n43), .PAD(q3[4]) );
  PAD_OUT q3_slice_5__po4 ( .I(n45), .PAD(q3[5]) );
  PAD_OUT q3_slice_6__po4 ( .I(n47), .PAD(q3[6]) );
  PAD_OUT q3_slice_7__po4 ( .I(n49), .PAD(q3[7]) );
  PAD_OUT q3_slice_8__po4 ( .I(n51), .PAD(q3[8]) );
  PAD_OUT q3_slice_9__po4 ( .I(n53), .PAD(q3[9]) );
  PAD_OUT q3_slice_10__po4 ( .I(n55), .PAD(q3[10]) );
  PAD_OUT q3_slice_11__po4 ( .I(n57), .PAD(q3[11]) );
  PAD_OUT q3_slice_12__po4 ( .I(n59), .PAD(q3[12]) );
  PAD_OUT q3_slice_13__po4 ( .I(n61), .PAD(q3[13]) );
  PAD_OUT q3_slice_14__po4 ( .I(n63), .PAD(q3[14]) );
  PAD_OUT q3_slice_15__po4 ( .I(n65), .PAD(q3[15]) );
  PAD_OUT q4_slice_0__po5 ( .I(n3), .PAD(q4[0]) );
  PAD_OUT q4_slice_1__po5 ( .I(n5), .PAD(q4[1]) );
  PAD_OUT q4_slice_2__po5 ( .I(n7), .PAD(q4[2]) );
  PAD_OUT q4_slice_3__po5 ( .I(n9), .PAD(q4[3]) );
  PAD_OUT q4_slice_4__po5 ( .I(n11), .PAD(q4[4]) );
  PAD_OUT q4_slice_5__po5 ( .I(n13), .PAD(q4[5]) );
  PAD_OUT q4_slice_6__po5 ( .I(n15), .PAD(q4[6]) );
  PAD_OUT q4_slice_7__po5 ( .I(n17), .PAD(q4[7]) );
  PAD_OUT q4_slice_8__po5 ( .I(n19), .PAD(q4[8]) );
  PAD_OUT q4_slice_9__po5 ( .I(n21), .PAD(q4[9]) );
  PAD_OUT q4_slice_10__po5 ( .I(n23), .PAD(q4[10]) );
  PAD_OUT q4_slice_11__po5 ( .I(n25), .PAD(q4[11]) );
  PAD_OUT q4_slice_12__po5 ( .I(n27), .PAD(q4[12]) );
  PAD_OUT q4_slice_13__po5 ( .I(n29), .PAD(q4[13]) );
  PAD_OUT q4_slice_14__po5 ( .I(n31), .PAD(q4[14]) );
  PAD_OUT q4_slice_15__po5 ( .I(n33), .PAD(q4[15]) );
  interleaver i0 ( .clk(clk1_c), .reset_n(reset_n_c), .di_rdy(di_rdy_c), 
        .do_acpt(do_acpt_out), .enable(1'b1), .di_data(di_data_c), .do_rdy(
        n132), .di_acpt(n131), .do_data({n133, n134, n135, n136, n137, n138, 
        n139, n140}) );
  async_bridge i1 ( .clk1(clk1_c), .clk2(clk2_c), .rstn(reset_n_c), 
        .do_rdy_in(do_rdy), .do_acpt_in(do_acpt), .do_acpt_out(do_acpt_out), 
        .do_rdy_out(do_rdy_out) );
  mem_ctrl mc0 ( .clk(clk2_gate), .rstn(reset_n_c), .do_rdy(do_rdy_out), 
        .mc_pwr(mc_pwr_c), .memsel(memsel_c), .mc_save(mc_save_c), 
        .mc_restore(mc_restore_c), .do_acpt(n141), .ceb({n142, n143, n144, 
        n145}), .web({n146, n147, n148, n149}), .addr({n150, n151, n152, n153, 
        n154, n155, n156, n157}) );
  sram_256x16 m1 ( .Q(q1_i), .A(address), .RSTB(reset_n_c),
        .D({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, do_data}),
        .PD(sram_pwr_c), .CLK(clk2_c), .CEB(ceb[0]), .WEB(web[0]));
  sram_256x16 m2 ( .Q(q2_i), .A(address), .RSTB(reset_n_c),
        .D({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, do_data}),
        .PD(sram_pwr_c), .CLK(clk2_c), .CEB(ceb[1]), .WEB(web[1]));
  sram_256x16 m3 (  .Q(q3_i), .A(address),.RSTB(reset_n_c),
        .D({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, do_data}),
        .PD(sram_pwr_c), .CLK(clk2_c), .CEB(ceb[2]), .WEB(web[2]));
  sram_256x16 m4 ( .Q(q4_i), .A(address), .RSTB(reset_n_c),
        .D({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, do_data}),
        .PD(sram_pwr_c), .CLK(clk2_c), .CEB(ceb[3]), .WEB(web[3]));
  ISO_LO ISO_addr_0__UPF_ISO ( .I(n158), .ISO(n174), .Z(address[0]) ); //synopsys isolation_upf mem_ctrl_iso_0+PD_mem_ctrl
  ISO_LO ISO_addr_1__UPF_ISO ( .I(n159), .ISO(n174), .Z(address[1]) ); //synopsys isolation_upf mem_ctrl_iso_0+PD_mem_ctrl
  ISO_LO ISO_addr_2__UPF_ISO ( .I(n160), .ISO(n174), .Z(address[2]) ); //synopsys isolation_upf mem_ctrl_iso_0+PD_mem_ctrl
  ISO_LO ISO_addr_3__UPF_ISO ( .I(n161), .ISO(n174), .Z(address[3]) ); //synopsys isolation_upf mem_ctrl_iso_0+PD_mem_ctrl
  ISO_LO ISO_addr_4__UPF_ISO ( .I(n162), .ISO(n174), .Z(address[4]) ); //synopsys isolation_upf mem_ctrl_iso_0+PD_mem_ctrl
  ISO_LO ISO_addr_5__UPF_ISO ( .I(n163), .ISO(n174), .Z(address[5]) ); //synopsys isolation_upf mem_ctrl_iso_0+PD_mem_ctrl
  ISO_LO ISO_addr_6__UPF_ISO ( .I(n164), .ISO(n174), .Z(address[6]) ); //synopsys isolation_upf mem_ctrl_iso_0+PD_mem_ctrl
  ISO_LO ISO_addr_7__UPF_ISO ( .I(n165), .ISO(n174), .Z(address[7]) ); //synopsys isolation_upf mem_ctrl_iso_0+PD_mem_ctrl
  ISO_HI ISO_web_0__UPF_ISO ( .I(n166), .ISO(n174), .Z(web[0]) ); //synopsys isolation_upf mem_ctrl_iso_1+PD_mem_ctrl
  ISO_HI ISO_web_1__UPF_ISO ( .I(n167), .ISO(n174), .Z(web[1]) ); //synopsys isolation_upf mem_ctrl_iso_1+PD_mem_ctrl
  ISO_HI ISO_web_2__UPF_ISO ( .I(n168), .ISO(n174), .Z(web[2]) ); //synopsys isolation_upf mem_ctrl_iso_1+PD_mem_ctrl
  ISO_HI ISO_web_3__UPF_ISO ( .I(n169), .ISO(n174), .Z(web[3]) ); //synopsys isolation_upf mem_ctrl_iso_1+PD_mem_ctrl
  ISO_HI ISO_ceb_0__UPF_ISO ( .I(n170), .ISO(n174), .Z(ceb[0]) ); //synopsys isolation_upf mem_ctrl_iso_1+PD_mem_ctrl
  ISO_HI ISO_ceb_1__UPF_ISO ( .I(n171), .ISO(n174), .Z(ceb[1]) ); //synopsys isolation_upf mem_ctrl_iso_1+PD_mem_ctrl
  ISO_HI ISO_ceb_2__UPF_ISO ( .I(n172), .ISO(n174), .Z(ceb[2]) ); //synopsys isolation_upf mem_ctrl_iso_1+PD_mem_ctrl
  ISO_HI ISO_ceb_3__UPF_ISO ( .I(n173), .ISO(n174), .Z(ceb[3]) ); //synopsys isolation_upf mem_ctrl_iso_1+PD_mem_ctrl
  ISO_LO ISO_do_acpt_UPF_ISO ( .I(n175), .ISO(n174), .Z(do_acpt) ); //synopsys isolation_upf mem_ctrl_iso_0+PD_mem_ctrl
  LS_LH LS_web_3__UPF_LS ( .I(n146), .Z(n169) );
  LS_LH LS_do_acpt_UPF_LS ( .I(n141), .Z(n175) );
  LS_LH LS_ceb_3__UPF_LS ( .I(n142), .Z(n173) );
  LS_LH LS_ceb_1__UPF_LS ( .I(n144), .Z(n171) );
  LS_LH LS_ceb_2__UPF_LS ( .I(n143), .Z(n172) );
  LS_LH LS_ceb_0__UPF_LS ( .I(n145), .Z(n170) );
  LS_LH LS_web_1__UPF_LS ( .I(n148), .Z(n167) );
  LS_LH LS_web_2__UPF_LS ( .I(n147), .Z(n168) );
  LS_LH LS_web_0__UPF_LS ( .I(n149), .Z(n166) );
  LS_LH LS_addr_4__UPF_LS ( .I(n153), .Z(n162) );
  LS_LH LS_addr_3__UPF_LS ( .I(n154), .Z(n161) );
  LS_LH LS_addr_2__UPF_LS ( .I(n155), .Z(n160) );
  LS_LH LS_addr_1__UPF_LS ( .I(n156), .Z(n159) );
  LS_LH LS_addr_0__UPF_LS ( .I(n157), .Z(n158) );
  LS_LH LS_do_data_7__UPF_LS ( .I(n133), .Z(do_data[7]) );
  LS_LH LS_do_data_6__UPF_LS ( .I(n134), .Z(do_data[6]) );
  LS_LH LS_do_data_5__UPF_LS ( .I(n135), .Z(do_data[5]) );
  LS_LH LS_do_data_4__UPF_LS ( .I(n136), .Z(do_data[4]) );
  LS_LH LS_do_data_3__UPF_LS ( .I(n137), .Z(do_data[3]) );
  LS_LH LS_do_data_2__UPF_LS ( .I(n138), .Z(do_data[2]) );
  LS_LH LS_do_data_1__UPF_LS ( .I(n139), .Z(do_data[1]) );
  LS_LH LS_do_data_0__UPF_LS ( .I(n140), .Z(do_data[0]) );
  LS_LH LS_do_rdy_UPF_LS ( .I(n132), .Z(do_rdy) );
  LS_LH LS_addr_5__UPF_LS ( .I(n152), .Z(n163) );
  LS_LH LS_addr_7__UPF_LS ( .I(n150), .Z(n165) );
  LS_LH LS_addr_6__UPF_LS ( .I(n151), .Z(n164) );
  LS_LH LS_di_acpt_UPF_LS ( .I(n131), .Z(di_acpt_i) );
  INV U5 ( .I(n2), .ZN(n3) );
  INV U6 ( .I(q4_i[0]), .ZN(n2) );
  INV U7 ( .I(n4), .ZN(n5) );
  INV U8 ( .I(q4_i[1]), .ZN(n4) );
  INV U9 ( .I(n6), .ZN(n7) );
  INV U10 ( .I(q4_i[2]), .ZN(n6) );
  INV U11 ( .I(n8), .ZN(n9) );
  INV U12 ( .I(q4_i[3]), .ZN(n8) );
  INV U13 ( .I(n10), .ZN(n11) );
  INV U14 ( .I(q4_i[4]), .ZN(n10) );
  INV U15 ( .I(n12), .ZN(n13) );
  INV U16 ( .I(q4_i[5]), .ZN(n12) );
  INV U17 ( .I(n14), .ZN(n15) );
  INV U18 ( .I(q4_i[6]), .ZN(n14) );
  INV U19 ( .I(n16), .ZN(n17) );
  INV U20 ( .I(q4_i[7]), .ZN(n16) );
  INV U21 ( .I(n18), .ZN(n19) );
  INV U22 ( .I(q4_i[8]), .ZN(n18) );
  INV U23 ( .I(n20), .ZN(n21) );
  INV U24 ( .I(q4_i[9]), .ZN(n20) );
  INV U25 ( .I(n22), .ZN(n23) );
  INV U26 ( .I(q4_i[10]), .ZN(n22) );
  INV U27 ( .I(n24), .ZN(n25) );
  INV U28 ( .I(q4_i[11]), .ZN(n24) );
  INV U29 ( .I(n26), .ZN(n27) );
  INV U30 ( .I(q4_i[12]), .ZN(n26) );
  INV U31 ( .I(n28), .ZN(n29) );
  INV U32 ( .I(q4_i[13]), .ZN(n28) );
  INV U33 ( .I(n30), .ZN(n31) );
  INV U34 ( .I(q4_i[14]), .ZN(n30) );
  INV U35 ( .I(n32), .ZN(n33) );
  INV U36 ( .I(q4_i[15]), .ZN(n32) );
  INV U37 ( .I(n34), .ZN(n35) );
  INV U38 ( .I(q3_i[0]), .ZN(n34) );
  INV U39 ( .I(n36), .ZN(n37) );
  INV U40 ( .I(q3_i[1]), .ZN(n36) );
  INV U41 ( .I(n38), .ZN(n39) );
  INV U42 ( .I(q3_i[2]), .ZN(n38) );
  INV U43 ( .I(n40), .ZN(n41) );
  INV U44 ( .I(q3_i[3]), .ZN(n40) );
  INV U45 ( .I(n42), .ZN(n43) );
  INV U46 ( .I(q3_i[4]), .ZN(n42) );
  INV U47 ( .I(n44), .ZN(n45) );
  INV U48 ( .I(q3_i[5]), .ZN(n44) );
  INV U49 ( .I(n46), .ZN(n47) );
  INV U50 ( .I(q3_i[6]), .ZN(n46) );
  INV U51 ( .I(n48), .ZN(n49) );
  INV U52 ( .I(q3_i[7]), .ZN(n48) );
  INV U53 ( .I(n50), .ZN(n51) );
  INV U54 ( .I(q3_i[8]), .ZN(n50) );
  INV U55 ( .I(n52), .ZN(n53) );
  INV U56 ( .I(q3_i[9]), .ZN(n52) );
  INV U57 ( .I(n54), .ZN(n55) );
  INV U58 ( .I(q3_i[10]), .ZN(n54) );
  INV U59 ( .I(n56), .ZN(n57) );
  INV U60 ( .I(q3_i[11]), .ZN(n56) );
  INV U61 ( .I(n58), .ZN(n59) );
  INV U62 ( .I(q3_i[12]), .ZN(n58) );
  INV U63 ( .I(n60), .ZN(n61) );
  INV U64 ( .I(q3_i[13]), .ZN(n60) );
  INV U65 ( .I(n62), .ZN(n63) );
  INV U66 ( .I(q3_i[14]), .ZN(n62) );
  INV U67 ( .I(n64), .ZN(n65) );
  INV U68 ( .I(q3_i[15]), .ZN(n64) );
  INV U69 ( .I(n66), .ZN(n67) );
  INV U70 ( .I(q2_i[0]), .ZN(n66) );
  INV U71 ( .I(n68), .ZN(n69) );
  INV U72 ( .I(q2_i[1]), .ZN(n68) );
  INV U73 ( .I(n70), .ZN(n71) );
  INV U74 ( .I(q2_i[2]), .ZN(n70) );
  INV U75 ( .I(n72), .ZN(n73) );
  INV U76 ( .I(q2_i[3]), .ZN(n72) );
  INV U77 ( .I(n74), .ZN(n75) );
  INV U78 ( .I(q2_i[4]), .ZN(n74) );
  INV U79 ( .I(n76), .ZN(n77) );
  INV U80 ( .I(q2_i[5]), .ZN(n76) );
  INV U81 ( .I(n78), .ZN(n79) );
  INV U82 ( .I(q2_i[6]), .ZN(n78) );
  INV U83 ( .I(n80), .ZN(n81) );
  INV U84 ( .I(q2_i[7]), .ZN(n80) );
  INV U85 ( .I(n82), .ZN(n83) );
  INV U86 ( .I(q2_i[8]), .ZN(n82) );
  INV U87 ( .I(n84), .ZN(n85) );
  INV U88 ( .I(q2_i[9]), .ZN(n84) );
  INV U89 ( .I(n86), .ZN(n87) );
  INV U90 ( .I(q2_i[10]), .ZN(n86) );
  INV U91 ( .I(n88), .ZN(n89) );
  INV U92 ( .I(q2_i[11]), .ZN(n88) );
  INV U93 ( .I(n90), .ZN(n91) );
  INV U94 ( .I(q2_i[12]), .ZN(n90) );
  INV U95 ( .I(n92), .ZN(n93) );
  INV U96 ( .I(q2_i[13]), .ZN(n92) );
  INV U97 ( .I(n94), .ZN(n95) );
  INV U98 ( .I(q2_i[14]), .ZN(n94) );
  INV U99 ( .I(n96), .ZN(n97) );
  INV U100 ( .I(q2_i[15]), .ZN(n96) );
  INV U101 ( .I(n98), .ZN(n99) );
  INV U102 ( .I(q1_i[0]), .ZN(n98) );
  INV U103 ( .I(n100), .ZN(n101) );
  INV U104 ( .I(q1_i[1]), .ZN(n100) );
  INV U105 ( .I(n102), .ZN(n103) );
  INV U106 ( .I(q1_i[2]), .ZN(n102) );
  INV U107 ( .I(n104), .ZN(n105) );
  INV U108 ( .I(q1_i[3]), .ZN(n104) );
  INV U109 ( .I(n106), .ZN(n107) );
  INV U110 ( .I(q1_i[4]), .ZN(n106) );
  INV U111 ( .I(q1_i[5]), .ZN(n108) );
  INV U112 ( .I(q1_i[6]), .ZN(n110) );
  INV U113 ( .I(q1_i[7]), .ZN(n112) );
  INV U114 ( .I(q1_i[8]), .ZN(n114) );
  INV U115 ( .I(q1_i[9]), .ZN(n116) );
  INV U116 ( .I(q1_i[10]), .ZN(n118) );
  INV U117 ( .I(q1_i[11]), .ZN(n120) );
  INV U118 ( .I(q1_i[12]), .ZN(n122) );
  INV U119 ( .I(q1_i[13]), .ZN(n124) );
  INV U120 ( .I(q1_i[14]), .ZN(n126) );
  INV U121 ( .I(q1_i[15]), .ZN(n128) );
  I_NOR2 U122 ( .A1(mc_clk_gate_c), .B1(n130), .ZN(clk2_gate) );
  INV U123 ( .I(n108), .ZN(n109) );
  INV U124 ( .I(n110), .ZN(n111) );
  INV U125 ( .I(n112), .ZN(n113) );
  INV U126 ( .I(n114), .ZN(n115) );
  INV U127 ( .I(n116), .ZN(n117) );
  INV U128 ( .I(n118), .ZN(n119) );
  INV U129 ( .I(n120), .ZN(n121) );
  INV U130 ( .I(n122), .ZN(n123) );
  INV U131 ( .I(n124), .ZN(n125) );
  INV U132 ( .I(n126), .ZN(n127) );
  INV U133 ( .I(n128), .ZN(n129) );
  INV U134 ( .I(clk2_c), .ZN(n130) );
endmodule

