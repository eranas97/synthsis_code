package interleaver_tr_pkg;

    import avm_pkg::*;
    `include "interleaver_transaction.svh"

endpackage // interleaver_tr_pkg
