module ripplecarryadder4(input [0:3]a,b,input cin,output cout);
wire [0:2]c;
