module testforsr;