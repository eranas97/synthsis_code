module bind_wrapper;
	bind send_receive receive_send inst_receive_send (.data_received(data_sent));
endmodule
