package fpu_agent_pkg;

import ovm_pkg::*;
`include "ovm_macros.svh";

`include "fpu_sv_utils.svh";
`include "fpu_tr.svh";

`include "fpu_sequencer.svh";
`include "fpu_sequence_driver.svh";
`include "fpu_monitor.svh";
`include "fpu_coverage.svh";

`include "fpu_agent.svh";


`include "fpu_sequence_library.svh";

endpackage // fpu_agent_pkg

