module 4_1mux(I0,I1,I2,I3,Y);
input I0,I1,I2,I3;
output Y;