module multiclock();
reg clk, clk1, clk2, clk3;
reg b0, b1, b2, b3, b4;

initial clk = 0; always #50 clk = ~clk;
initial clk1 = 0; always #51 clk1 = ~clk1;

assert property (@(posedge clk) b0 ##1 (1 ##1 (@(posedge clk1) b1) and (@(posedge clk) b2)) |=> b3);

initial
begin
    #100     b0 = 1;   b1 = 0;   b2 = 0;    b3 = 0; //100
    #100     b0 = 0;   b1 = 1;   b2 = 1;    b3 = 0; //200
    #100     b0 = 0;   b1 = 0;   b2 = 0;    b3 = 1; //300
    #100     b0 = 0;   b1 = 0;   b2 = 0;    b3 = 0; //400
    #100     b0 = 0;   b1 = 0;   b2 = 0;    b3 = 0; //500
    #100     b0 = 1;   b1 = 0;   b2 = 0;    b3 = 0; //600
    #100     b0 = 0;   b1 = 1;   b2 = 0;    b3 = 0; //700
    #100     b0 = 0;   b1 = 0;   b2 = 0;    b3 = 0; //800
    #100     b0 = 1;   b1 = 0;   b2 = 0;    b3 = 0; //900
    #100     b0 = 0;   b1 = 1;   b2 = 1;    b3 = 0; //1000
    #100     b0 = 1;   b1 = 0;   b2 = 0;    b3 = 0; //1100
    #100     b0 = 0;   b1 = 1;   b2 = 1;    b3 = 0; //1200
    #100     b0 = 0;   b1 = 0;   b2 = 0;    b3 = 1; //1300
    #100     b0 = 0;   b1 = 0;   b2 = 0;    b3 = 0; //1400
    #100     b0 = 0;   b1 = 0;   b2 = 0;    b3 = 0; //1500
    #100     b0 = 0;   b1 = 0;   b2 = 0;    b3 = 0; //1600
    #100     b0 = 0;   b1 = 0;   b2 = 0;    b3 = 0; //1700
    #100     b0 = 0;   b1 = 0;   b2 = 0;    b3 = 0; //1800
    #100     b0 = 0;   b1 = 0;   b2 = 0;    b3 = 0; //1900
    #100     b0 = 0;   b1 = 0;   b2 = 0;    b3 = 0; //2000
    #100     b0 = 0;   b1 = 0;   b2 = 0;    b3 = 0; //2100
    #100     b0 = 0;   b1 = 0;   b2 = 0;    b3 = 0; //2200
    #100     b0 = 0;   b1 = 0;   b2 = 0;    b3 = 0; //2300
    #100     b0 = 0;   b1 = 0;   b2 = 0;    b3 = 0; //2400
    #100     b0 = 0;   b1 = 0;   b2 = 0;    b3 = 0; //2500
    #100     b0 = 0;   b1 = 0;   b2 = 0;    b3 = 0; //2600
	#500 $finish;
end
endmodule




